

module bsg_link_iddr_phy_width_p9
(
  clk_i,
  data_i,
  data_r_o,
  rst
);

  input [8:0] data_i;
  output [17:0] data_r_o;
  input clk_i;
  input rst;
  wire [17:0] data_r_o;
  wire N0;
  wire [8:0] data_p_r,data_n_r;
  reg data_p_r_8_sv2v_reg,data_p_r_7_sv2v_reg,data_p_r_6_sv2v_reg,data_p_r_5_sv2v_reg,
  data_p_r_4_sv2v_reg,data_p_r_3_sv2v_reg,data_p_r_2_sv2v_reg,data_p_r_1_sv2v_reg,
  data_p_r_0_sv2v_reg,data_n_r_8_sv2v_reg,data_n_r_7_sv2v_reg,data_n_r_6_sv2v_reg,
  data_n_r_5_sv2v_reg,data_n_r_4_sv2v_reg,data_n_r_3_sv2v_reg,data_n_r_2_sv2v_reg,
  data_n_r_1_sv2v_reg,data_n_r_0_sv2v_reg,data_r_o_17_sv2v_reg,
  data_r_o_16_sv2v_reg,data_r_o_15_sv2v_reg,data_r_o_14_sv2v_reg,data_r_o_13_sv2v_reg,
  data_r_o_12_sv2v_reg,data_r_o_11_sv2v_reg,data_r_o_10_sv2v_reg,data_r_o_9_sv2v_reg,
  data_r_o_8_sv2v_reg,data_r_o_7_sv2v_reg,data_r_o_6_sv2v_reg,data_r_o_5_sv2v_reg,
  data_r_o_4_sv2v_reg,data_r_o_3_sv2v_reg,data_r_o_2_sv2v_reg,data_r_o_1_sv2v_reg,
  data_r_o_0_sv2v_reg;
  assign data_p_r[8] = data_p_r_8_sv2v_reg;
  assign data_p_r[7] = data_p_r_7_sv2v_reg;
  assign data_p_r[6] = data_p_r_6_sv2v_reg;
  assign data_p_r[5] = data_p_r_5_sv2v_reg;
  assign data_p_r[4] = data_p_r_4_sv2v_reg;
  assign data_p_r[3] = data_p_r_3_sv2v_reg;
  assign data_p_r[2] = data_p_r_2_sv2v_reg;
  assign data_p_r[1] = data_p_r_1_sv2v_reg;
  assign data_p_r[0] = data_p_r_0_sv2v_reg;
  assign data_n_r[8] = data_n_r_8_sv2v_reg;
  assign data_n_r[7] = data_n_r_7_sv2v_reg;
  assign data_n_r[6] = data_n_r_6_sv2v_reg;
  assign data_n_r[5] = data_n_r_5_sv2v_reg;
  assign data_n_r[4] = data_n_r_4_sv2v_reg;
  assign data_n_r[3] = data_n_r_3_sv2v_reg;
  assign data_n_r[2] = data_n_r_2_sv2v_reg;
  assign data_n_r[1] = data_n_r_1_sv2v_reg;
  assign data_n_r[0] = data_n_r_0_sv2v_reg;
  assign data_r_o[17] = data_r_o_17_sv2v_reg;
  assign data_r_o[16] = data_r_o_16_sv2v_reg;
  assign data_r_o[15] = data_r_o_15_sv2v_reg;
  assign data_r_o[14] = data_r_o_14_sv2v_reg;
  assign data_r_o[13] = data_r_o_13_sv2v_reg;
  assign data_r_o[12] = data_r_o_12_sv2v_reg;
  assign data_r_o[11] = data_r_o_11_sv2v_reg;
  assign data_r_o[10] = data_r_o_10_sv2v_reg;
  assign data_r_o[9] = data_r_o_9_sv2v_reg;
  assign data_r_o[8] = data_r_o_8_sv2v_reg;
  assign data_r_o[7] = data_r_o_7_sv2v_reg;
  assign data_r_o[6] = data_r_o_6_sv2v_reg;
  assign data_r_o[5] = data_r_o_5_sv2v_reg;
  assign data_r_o[4] = data_r_o_4_sv2v_reg;
  assign data_r_o[3] = data_r_o_3_sv2v_reg;
  assign data_r_o[2] = data_r_o_2_sv2v_reg;
  assign data_r_o[1] = data_r_o_1_sv2v_reg;
  assign data_r_o[0] = data_r_o_0_sv2v_reg;
  assign N0 = ~clk_i;

  always @(posedge clk_i) begin
  if (rst) begin
    data_p_r_8_sv2v_reg <= 1'b0;
    data_r_o_8_sv2v_reg <= 1'b0;
    
  end
  else begin
      data_p_r_8_sv2v_reg <= data_i[8];
      data_p_r_7_sv2v_reg <= data_i[7];
      data_p_r_6_sv2v_reg <= data_i[6];
      data_p_r_5_sv2v_reg <= data_i[5];
      data_p_r_4_sv2v_reg <= data_i[4];
      data_p_r_3_sv2v_reg <= data_i[3];
      data_p_r_2_sv2v_reg <= data_i[2];
      data_p_r_1_sv2v_reg <= data_i[1];
      data_p_r_0_sv2v_reg <= data_i[0];
      data_r_o_17_sv2v_reg <= data_n_r[8];
      data_r_o_16_sv2v_reg <= data_n_r[7];
      data_r_o_15_sv2v_reg <= data_n_r[6];
      data_r_o_14_sv2v_reg <= data_n_r[5];
      data_r_o_13_sv2v_reg <= data_n_r[4];
      data_r_o_12_sv2v_reg <= data_n_r[3];
      data_r_o_11_sv2v_reg <= data_n_r[2];
      data_r_o_10_sv2v_reg <= data_n_r[1];
      data_r_o_9_sv2v_reg <= data_n_r[0];
      data_r_o_8_sv2v_reg <= data_p_r[8];
      data_r_o_7_sv2v_reg <= data_p_r[7];
      data_r_o_6_sv2v_reg <= data_p_r[6];
      data_r_o_5_sv2v_reg <= data_p_r[5];
      data_r_o_4_sv2v_reg <= data_p_r[4];
      data_r_o_3_sv2v_reg <= data_p_r[3];
      data_r_o_2_sv2v_reg <= data_p_r[2];
      data_r_o_1_sv2v_reg <= data_p_r[1];
      data_r_o_0_sv2v_reg <= data_p_r[0];
    end 
  end


  always @(posedge N0) begin
    if(1'b1) begin
      data_n_r_8_sv2v_reg <= data_i[8];
      data_n_r_7_sv2v_reg <= data_i[7];
      data_n_r_6_sv2v_reg <= data_i[6];
      data_n_r_5_sv2v_reg <= data_i[5];
      data_n_r_4_sv2v_reg <= data_i[4];
      data_n_r_3_sv2v_reg <= data_i[3];
      data_n_r_2_sv2v_reg <= data_i[2];
      data_n_r_1_sv2v_reg <= data_i[1];
      data_n_r_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_synth_width_p16_els_p64_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [5:0] w_addr_i;
  input [15:0] w_data_i;
  input [5:0] r_addr_i;
  output [15:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [15:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294;
  wire [1023:0] mem;
  reg mem_1023_sv2v_reg,mem_1022_sv2v_reg,mem_1021_sv2v_reg,mem_1020_sv2v_reg,
  mem_1019_sv2v_reg,mem_1018_sv2v_reg,mem_1017_sv2v_reg,mem_1016_sv2v_reg,
  mem_1015_sv2v_reg,mem_1014_sv2v_reg,mem_1013_sv2v_reg,mem_1012_sv2v_reg,mem_1011_sv2v_reg,
  mem_1010_sv2v_reg,mem_1009_sv2v_reg,mem_1008_sv2v_reg,mem_1007_sv2v_reg,
  mem_1006_sv2v_reg,mem_1005_sv2v_reg,mem_1004_sv2v_reg,mem_1003_sv2v_reg,mem_1002_sv2v_reg,
  mem_1001_sv2v_reg,mem_1000_sv2v_reg,mem_999_sv2v_reg,mem_998_sv2v_reg,
  mem_997_sv2v_reg,mem_996_sv2v_reg,mem_995_sv2v_reg,mem_994_sv2v_reg,mem_993_sv2v_reg,
  mem_992_sv2v_reg,mem_991_sv2v_reg,mem_990_sv2v_reg,mem_989_sv2v_reg,mem_988_sv2v_reg,
  mem_987_sv2v_reg,mem_986_sv2v_reg,mem_985_sv2v_reg,mem_984_sv2v_reg,
  mem_983_sv2v_reg,mem_982_sv2v_reg,mem_981_sv2v_reg,mem_980_sv2v_reg,mem_979_sv2v_reg,
  mem_978_sv2v_reg,mem_977_sv2v_reg,mem_976_sv2v_reg,mem_975_sv2v_reg,mem_974_sv2v_reg,
  mem_973_sv2v_reg,mem_972_sv2v_reg,mem_971_sv2v_reg,mem_970_sv2v_reg,mem_969_sv2v_reg,
  mem_968_sv2v_reg,mem_967_sv2v_reg,mem_966_sv2v_reg,mem_965_sv2v_reg,
  mem_964_sv2v_reg,mem_963_sv2v_reg,mem_962_sv2v_reg,mem_961_sv2v_reg,mem_960_sv2v_reg,
  mem_959_sv2v_reg,mem_958_sv2v_reg,mem_957_sv2v_reg,mem_956_sv2v_reg,mem_955_sv2v_reg,
  mem_954_sv2v_reg,mem_953_sv2v_reg,mem_952_sv2v_reg,mem_951_sv2v_reg,
  mem_950_sv2v_reg,mem_949_sv2v_reg,mem_948_sv2v_reg,mem_947_sv2v_reg,mem_946_sv2v_reg,
  mem_945_sv2v_reg,mem_944_sv2v_reg,mem_943_sv2v_reg,mem_942_sv2v_reg,mem_941_sv2v_reg,
  mem_940_sv2v_reg,mem_939_sv2v_reg,mem_938_sv2v_reg,mem_937_sv2v_reg,mem_936_sv2v_reg,
  mem_935_sv2v_reg,mem_934_sv2v_reg,mem_933_sv2v_reg,mem_932_sv2v_reg,
  mem_931_sv2v_reg,mem_930_sv2v_reg,mem_929_sv2v_reg,mem_928_sv2v_reg,mem_927_sv2v_reg,
  mem_926_sv2v_reg,mem_925_sv2v_reg,mem_924_sv2v_reg,mem_923_sv2v_reg,mem_922_sv2v_reg,
  mem_921_sv2v_reg,mem_920_sv2v_reg,mem_919_sv2v_reg,mem_918_sv2v_reg,
  mem_917_sv2v_reg,mem_916_sv2v_reg,mem_915_sv2v_reg,mem_914_sv2v_reg,mem_913_sv2v_reg,
  mem_912_sv2v_reg,mem_911_sv2v_reg,mem_910_sv2v_reg,mem_909_sv2v_reg,mem_908_sv2v_reg,
  mem_907_sv2v_reg,mem_906_sv2v_reg,mem_905_sv2v_reg,mem_904_sv2v_reg,
  mem_903_sv2v_reg,mem_902_sv2v_reg,mem_901_sv2v_reg,mem_900_sv2v_reg,mem_899_sv2v_reg,
  mem_898_sv2v_reg,mem_897_sv2v_reg,mem_896_sv2v_reg,mem_895_sv2v_reg,mem_894_sv2v_reg,
  mem_893_sv2v_reg,mem_892_sv2v_reg,mem_891_sv2v_reg,mem_890_sv2v_reg,mem_889_sv2v_reg,
  mem_888_sv2v_reg,mem_887_sv2v_reg,mem_886_sv2v_reg,mem_885_sv2v_reg,
  mem_884_sv2v_reg,mem_883_sv2v_reg,mem_882_sv2v_reg,mem_881_sv2v_reg,mem_880_sv2v_reg,
  mem_879_sv2v_reg,mem_878_sv2v_reg,mem_877_sv2v_reg,mem_876_sv2v_reg,mem_875_sv2v_reg,
  mem_874_sv2v_reg,mem_873_sv2v_reg,mem_872_sv2v_reg,mem_871_sv2v_reg,
  mem_870_sv2v_reg,mem_869_sv2v_reg,mem_868_sv2v_reg,mem_867_sv2v_reg,mem_866_sv2v_reg,
  mem_865_sv2v_reg,mem_864_sv2v_reg,mem_863_sv2v_reg,mem_862_sv2v_reg,mem_861_sv2v_reg,
  mem_860_sv2v_reg,mem_859_sv2v_reg,mem_858_sv2v_reg,mem_857_sv2v_reg,mem_856_sv2v_reg,
  mem_855_sv2v_reg,mem_854_sv2v_reg,mem_853_sv2v_reg,mem_852_sv2v_reg,
  mem_851_sv2v_reg,mem_850_sv2v_reg,mem_849_sv2v_reg,mem_848_sv2v_reg,mem_847_sv2v_reg,
  mem_846_sv2v_reg,mem_845_sv2v_reg,mem_844_sv2v_reg,mem_843_sv2v_reg,mem_842_sv2v_reg,
  mem_841_sv2v_reg,mem_840_sv2v_reg,mem_839_sv2v_reg,mem_838_sv2v_reg,
  mem_837_sv2v_reg,mem_836_sv2v_reg,mem_835_sv2v_reg,mem_834_sv2v_reg,mem_833_sv2v_reg,
  mem_832_sv2v_reg,mem_831_sv2v_reg,mem_830_sv2v_reg,mem_829_sv2v_reg,mem_828_sv2v_reg,
  mem_827_sv2v_reg,mem_826_sv2v_reg,mem_825_sv2v_reg,mem_824_sv2v_reg,
  mem_823_sv2v_reg,mem_822_sv2v_reg,mem_821_sv2v_reg,mem_820_sv2v_reg,mem_819_sv2v_reg,
  mem_818_sv2v_reg,mem_817_sv2v_reg,mem_816_sv2v_reg,mem_815_sv2v_reg,mem_814_sv2v_reg,
  mem_813_sv2v_reg,mem_812_sv2v_reg,mem_811_sv2v_reg,mem_810_sv2v_reg,mem_809_sv2v_reg,
  mem_808_sv2v_reg,mem_807_sv2v_reg,mem_806_sv2v_reg,mem_805_sv2v_reg,
  mem_804_sv2v_reg,mem_803_sv2v_reg,mem_802_sv2v_reg,mem_801_sv2v_reg,mem_800_sv2v_reg,
  mem_799_sv2v_reg,mem_798_sv2v_reg,mem_797_sv2v_reg,mem_796_sv2v_reg,mem_795_sv2v_reg,
  mem_794_sv2v_reg,mem_793_sv2v_reg,mem_792_sv2v_reg,mem_791_sv2v_reg,
  mem_790_sv2v_reg,mem_789_sv2v_reg,mem_788_sv2v_reg,mem_787_sv2v_reg,mem_786_sv2v_reg,
  mem_785_sv2v_reg,mem_784_sv2v_reg,mem_783_sv2v_reg,mem_782_sv2v_reg,mem_781_sv2v_reg,
  mem_780_sv2v_reg,mem_779_sv2v_reg,mem_778_sv2v_reg,mem_777_sv2v_reg,mem_776_sv2v_reg,
  mem_775_sv2v_reg,mem_774_sv2v_reg,mem_773_sv2v_reg,mem_772_sv2v_reg,
  mem_771_sv2v_reg,mem_770_sv2v_reg,mem_769_sv2v_reg,mem_768_sv2v_reg,mem_767_sv2v_reg,
  mem_766_sv2v_reg,mem_765_sv2v_reg,mem_764_sv2v_reg,mem_763_sv2v_reg,mem_762_sv2v_reg,
  mem_761_sv2v_reg,mem_760_sv2v_reg,mem_759_sv2v_reg,mem_758_sv2v_reg,
  mem_757_sv2v_reg,mem_756_sv2v_reg,mem_755_sv2v_reg,mem_754_sv2v_reg,mem_753_sv2v_reg,
  mem_752_sv2v_reg,mem_751_sv2v_reg,mem_750_sv2v_reg,mem_749_sv2v_reg,mem_748_sv2v_reg,
  mem_747_sv2v_reg,mem_746_sv2v_reg,mem_745_sv2v_reg,mem_744_sv2v_reg,
  mem_743_sv2v_reg,mem_742_sv2v_reg,mem_741_sv2v_reg,mem_740_sv2v_reg,mem_739_sv2v_reg,
  mem_738_sv2v_reg,mem_737_sv2v_reg,mem_736_sv2v_reg,mem_735_sv2v_reg,mem_734_sv2v_reg,
  mem_733_sv2v_reg,mem_732_sv2v_reg,mem_731_sv2v_reg,mem_730_sv2v_reg,mem_729_sv2v_reg,
  mem_728_sv2v_reg,mem_727_sv2v_reg,mem_726_sv2v_reg,mem_725_sv2v_reg,
  mem_724_sv2v_reg,mem_723_sv2v_reg,mem_722_sv2v_reg,mem_721_sv2v_reg,mem_720_sv2v_reg,
  mem_719_sv2v_reg,mem_718_sv2v_reg,mem_717_sv2v_reg,mem_716_sv2v_reg,mem_715_sv2v_reg,
  mem_714_sv2v_reg,mem_713_sv2v_reg,mem_712_sv2v_reg,mem_711_sv2v_reg,
  mem_710_sv2v_reg,mem_709_sv2v_reg,mem_708_sv2v_reg,mem_707_sv2v_reg,mem_706_sv2v_reg,
  mem_705_sv2v_reg,mem_704_sv2v_reg,mem_703_sv2v_reg,mem_702_sv2v_reg,mem_701_sv2v_reg,
  mem_700_sv2v_reg,mem_699_sv2v_reg,mem_698_sv2v_reg,mem_697_sv2v_reg,mem_696_sv2v_reg,
  mem_695_sv2v_reg,mem_694_sv2v_reg,mem_693_sv2v_reg,mem_692_sv2v_reg,
  mem_691_sv2v_reg,mem_690_sv2v_reg,mem_689_sv2v_reg,mem_688_sv2v_reg,mem_687_sv2v_reg,
  mem_686_sv2v_reg,mem_685_sv2v_reg,mem_684_sv2v_reg,mem_683_sv2v_reg,mem_682_sv2v_reg,
  mem_681_sv2v_reg,mem_680_sv2v_reg,mem_679_sv2v_reg,mem_678_sv2v_reg,
  mem_677_sv2v_reg,mem_676_sv2v_reg,mem_675_sv2v_reg,mem_674_sv2v_reg,mem_673_sv2v_reg,
  mem_672_sv2v_reg,mem_671_sv2v_reg,mem_670_sv2v_reg,mem_669_sv2v_reg,mem_668_sv2v_reg,
  mem_667_sv2v_reg,mem_666_sv2v_reg,mem_665_sv2v_reg,mem_664_sv2v_reg,
  mem_663_sv2v_reg,mem_662_sv2v_reg,mem_661_sv2v_reg,mem_660_sv2v_reg,mem_659_sv2v_reg,
  mem_658_sv2v_reg,mem_657_sv2v_reg,mem_656_sv2v_reg,mem_655_sv2v_reg,mem_654_sv2v_reg,
  mem_653_sv2v_reg,mem_652_sv2v_reg,mem_651_sv2v_reg,mem_650_sv2v_reg,mem_649_sv2v_reg,
  mem_648_sv2v_reg,mem_647_sv2v_reg,mem_646_sv2v_reg,mem_645_sv2v_reg,
  mem_644_sv2v_reg,mem_643_sv2v_reg,mem_642_sv2v_reg,mem_641_sv2v_reg,mem_640_sv2v_reg,
  mem_639_sv2v_reg,mem_638_sv2v_reg,mem_637_sv2v_reg,mem_636_sv2v_reg,mem_635_sv2v_reg,
  mem_634_sv2v_reg,mem_633_sv2v_reg,mem_632_sv2v_reg,mem_631_sv2v_reg,
  mem_630_sv2v_reg,mem_629_sv2v_reg,mem_628_sv2v_reg,mem_627_sv2v_reg,mem_626_sv2v_reg,
  mem_625_sv2v_reg,mem_624_sv2v_reg,mem_623_sv2v_reg,mem_622_sv2v_reg,mem_621_sv2v_reg,
  mem_620_sv2v_reg,mem_619_sv2v_reg,mem_618_sv2v_reg,mem_617_sv2v_reg,mem_616_sv2v_reg,
  mem_615_sv2v_reg,mem_614_sv2v_reg,mem_613_sv2v_reg,mem_612_sv2v_reg,
  mem_611_sv2v_reg,mem_610_sv2v_reg,mem_609_sv2v_reg,mem_608_sv2v_reg,mem_607_sv2v_reg,
  mem_606_sv2v_reg,mem_605_sv2v_reg,mem_604_sv2v_reg,mem_603_sv2v_reg,mem_602_sv2v_reg,
  mem_601_sv2v_reg,mem_600_sv2v_reg,mem_599_sv2v_reg,mem_598_sv2v_reg,
  mem_597_sv2v_reg,mem_596_sv2v_reg,mem_595_sv2v_reg,mem_594_sv2v_reg,mem_593_sv2v_reg,
  mem_592_sv2v_reg,mem_591_sv2v_reg,mem_590_sv2v_reg,mem_589_sv2v_reg,mem_588_sv2v_reg,
  mem_587_sv2v_reg,mem_586_sv2v_reg,mem_585_sv2v_reg,mem_584_sv2v_reg,
  mem_583_sv2v_reg,mem_582_sv2v_reg,mem_581_sv2v_reg,mem_580_sv2v_reg,mem_579_sv2v_reg,
  mem_578_sv2v_reg,mem_577_sv2v_reg,mem_576_sv2v_reg,mem_575_sv2v_reg,mem_574_sv2v_reg,
  mem_573_sv2v_reg,mem_572_sv2v_reg,mem_571_sv2v_reg,mem_570_sv2v_reg,mem_569_sv2v_reg,
  mem_568_sv2v_reg,mem_567_sv2v_reg,mem_566_sv2v_reg,mem_565_sv2v_reg,
  mem_564_sv2v_reg,mem_563_sv2v_reg,mem_562_sv2v_reg,mem_561_sv2v_reg,mem_560_sv2v_reg,
  mem_559_sv2v_reg,mem_558_sv2v_reg,mem_557_sv2v_reg,mem_556_sv2v_reg,mem_555_sv2v_reg,
  mem_554_sv2v_reg,mem_553_sv2v_reg,mem_552_sv2v_reg,mem_551_sv2v_reg,
  mem_550_sv2v_reg,mem_549_sv2v_reg,mem_548_sv2v_reg,mem_547_sv2v_reg,mem_546_sv2v_reg,
  mem_545_sv2v_reg,mem_544_sv2v_reg,mem_543_sv2v_reg,mem_542_sv2v_reg,mem_541_sv2v_reg,
  mem_540_sv2v_reg,mem_539_sv2v_reg,mem_538_sv2v_reg,mem_537_sv2v_reg,mem_536_sv2v_reg,
  mem_535_sv2v_reg,mem_534_sv2v_reg,mem_533_sv2v_reg,mem_532_sv2v_reg,
  mem_531_sv2v_reg,mem_530_sv2v_reg,mem_529_sv2v_reg,mem_528_sv2v_reg,mem_527_sv2v_reg,
  mem_526_sv2v_reg,mem_525_sv2v_reg,mem_524_sv2v_reg,mem_523_sv2v_reg,mem_522_sv2v_reg,
  mem_521_sv2v_reg,mem_520_sv2v_reg,mem_519_sv2v_reg,mem_518_sv2v_reg,
  mem_517_sv2v_reg,mem_516_sv2v_reg,mem_515_sv2v_reg,mem_514_sv2v_reg,mem_513_sv2v_reg,
  mem_512_sv2v_reg,mem_511_sv2v_reg,mem_510_sv2v_reg,mem_509_sv2v_reg,mem_508_sv2v_reg,
  mem_507_sv2v_reg,mem_506_sv2v_reg,mem_505_sv2v_reg,mem_504_sv2v_reg,
  mem_503_sv2v_reg,mem_502_sv2v_reg,mem_501_sv2v_reg,mem_500_sv2v_reg,mem_499_sv2v_reg,
  mem_498_sv2v_reg,mem_497_sv2v_reg,mem_496_sv2v_reg,mem_495_sv2v_reg,mem_494_sv2v_reg,
  mem_493_sv2v_reg,mem_492_sv2v_reg,mem_491_sv2v_reg,mem_490_sv2v_reg,mem_489_sv2v_reg,
  mem_488_sv2v_reg,mem_487_sv2v_reg,mem_486_sv2v_reg,mem_485_sv2v_reg,
  mem_484_sv2v_reg,mem_483_sv2v_reg,mem_482_sv2v_reg,mem_481_sv2v_reg,mem_480_sv2v_reg,
  mem_479_sv2v_reg,mem_478_sv2v_reg,mem_477_sv2v_reg,mem_476_sv2v_reg,mem_475_sv2v_reg,
  mem_474_sv2v_reg,mem_473_sv2v_reg,mem_472_sv2v_reg,mem_471_sv2v_reg,
  mem_470_sv2v_reg,mem_469_sv2v_reg,mem_468_sv2v_reg,mem_467_sv2v_reg,mem_466_sv2v_reg,
  mem_465_sv2v_reg,mem_464_sv2v_reg,mem_463_sv2v_reg,mem_462_sv2v_reg,mem_461_sv2v_reg,
  mem_460_sv2v_reg,mem_459_sv2v_reg,mem_458_sv2v_reg,mem_457_sv2v_reg,mem_456_sv2v_reg,
  mem_455_sv2v_reg,mem_454_sv2v_reg,mem_453_sv2v_reg,mem_452_sv2v_reg,
  mem_451_sv2v_reg,mem_450_sv2v_reg,mem_449_sv2v_reg,mem_448_sv2v_reg,mem_447_sv2v_reg,
  mem_446_sv2v_reg,mem_445_sv2v_reg,mem_444_sv2v_reg,mem_443_sv2v_reg,mem_442_sv2v_reg,
  mem_441_sv2v_reg,mem_440_sv2v_reg,mem_439_sv2v_reg,mem_438_sv2v_reg,
  mem_437_sv2v_reg,mem_436_sv2v_reg,mem_435_sv2v_reg,mem_434_sv2v_reg,mem_433_sv2v_reg,
  mem_432_sv2v_reg,mem_431_sv2v_reg,mem_430_sv2v_reg,mem_429_sv2v_reg,mem_428_sv2v_reg,
  mem_427_sv2v_reg,mem_426_sv2v_reg,mem_425_sv2v_reg,mem_424_sv2v_reg,
  mem_423_sv2v_reg,mem_422_sv2v_reg,mem_421_sv2v_reg,mem_420_sv2v_reg,mem_419_sv2v_reg,
  mem_418_sv2v_reg,mem_417_sv2v_reg,mem_416_sv2v_reg,mem_415_sv2v_reg,mem_414_sv2v_reg,
  mem_413_sv2v_reg,mem_412_sv2v_reg,mem_411_sv2v_reg,mem_410_sv2v_reg,mem_409_sv2v_reg,
  mem_408_sv2v_reg,mem_407_sv2v_reg,mem_406_sv2v_reg,mem_405_sv2v_reg,
  mem_404_sv2v_reg,mem_403_sv2v_reg,mem_402_sv2v_reg,mem_401_sv2v_reg,mem_400_sv2v_reg,
  mem_399_sv2v_reg,mem_398_sv2v_reg,mem_397_sv2v_reg,mem_396_sv2v_reg,mem_395_sv2v_reg,
  mem_394_sv2v_reg,mem_393_sv2v_reg,mem_392_sv2v_reg,mem_391_sv2v_reg,
  mem_390_sv2v_reg,mem_389_sv2v_reg,mem_388_sv2v_reg,mem_387_sv2v_reg,mem_386_sv2v_reg,
  mem_385_sv2v_reg,mem_384_sv2v_reg,mem_383_sv2v_reg,mem_382_sv2v_reg,mem_381_sv2v_reg,
  mem_380_sv2v_reg,mem_379_sv2v_reg,mem_378_sv2v_reg,mem_377_sv2v_reg,mem_376_sv2v_reg,
  mem_375_sv2v_reg,mem_374_sv2v_reg,mem_373_sv2v_reg,mem_372_sv2v_reg,
  mem_371_sv2v_reg,mem_370_sv2v_reg,mem_369_sv2v_reg,mem_368_sv2v_reg,mem_367_sv2v_reg,
  mem_366_sv2v_reg,mem_365_sv2v_reg,mem_364_sv2v_reg,mem_363_sv2v_reg,mem_362_sv2v_reg,
  mem_361_sv2v_reg,mem_360_sv2v_reg,mem_359_sv2v_reg,mem_358_sv2v_reg,
  mem_357_sv2v_reg,mem_356_sv2v_reg,mem_355_sv2v_reg,mem_354_sv2v_reg,mem_353_sv2v_reg,
  mem_352_sv2v_reg,mem_351_sv2v_reg,mem_350_sv2v_reg,mem_349_sv2v_reg,mem_348_sv2v_reg,
  mem_347_sv2v_reg,mem_346_sv2v_reg,mem_345_sv2v_reg,mem_344_sv2v_reg,
  mem_343_sv2v_reg,mem_342_sv2v_reg,mem_341_sv2v_reg,mem_340_sv2v_reg,mem_339_sv2v_reg,
  mem_338_sv2v_reg,mem_337_sv2v_reg,mem_336_sv2v_reg,mem_335_sv2v_reg,mem_334_sv2v_reg,
  mem_333_sv2v_reg,mem_332_sv2v_reg,mem_331_sv2v_reg,mem_330_sv2v_reg,mem_329_sv2v_reg,
  mem_328_sv2v_reg,mem_327_sv2v_reg,mem_326_sv2v_reg,mem_325_sv2v_reg,
  mem_324_sv2v_reg,mem_323_sv2v_reg,mem_322_sv2v_reg,mem_321_sv2v_reg,mem_320_sv2v_reg,
  mem_319_sv2v_reg,mem_318_sv2v_reg,mem_317_sv2v_reg,mem_316_sv2v_reg,mem_315_sv2v_reg,
  mem_314_sv2v_reg,mem_313_sv2v_reg,mem_312_sv2v_reg,mem_311_sv2v_reg,
  mem_310_sv2v_reg,mem_309_sv2v_reg,mem_308_sv2v_reg,mem_307_sv2v_reg,mem_306_sv2v_reg,
  mem_305_sv2v_reg,mem_304_sv2v_reg,mem_303_sv2v_reg,mem_302_sv2v_reg,mem_301_sv2v_reg,
  mem_300_sv2v_reg,mem_299_sv2v_reg,mem_298_sv2v_reg,mem_297_sv2v_reg,mem_296_sv2v_reg,
  mem_295_sv2v_reg,mem_294_sv2v_reg,mem_293_sv2v_reg,mem_292_sv2v_reg,
  mem_291_sv2v_reg,mem_290_sv2v_reg,mem_289_sv2v_reg,mem_288_sv2v_reg,mem_287_sv2v_reg,
  mem_286_sv2v_reg,mem_285_sv2v_reg,mem_284_sv2v_reg,mem_283_sv2v_reg,mem_282_sv2v_reg,
  mem_281_sv2v_reg,mem_280_sv2v_reg,mem_279_sv2v_reg,mem_278_sv2v_reg,
  mem_277_sv2v_reg,mem_276_sv2v_reg,mem_275_sv2v_reg,mem_274_sv2v_reg,mem_273_sv2v_reg,
  mem_272_sv2v_reg,mem_271_sv2v_reg,mem_270_sv2v_reg,mem_269_sv2v_reg,mem_268_sv2v_reg,
  mem_267_sv2v_reg,mem_266_sv2v_reg,mem_265_sv2v_reg,mem_264_sv2v_reg,
  mem_263_sv2v_reg,mem_262_sv2v_reg,mem_261_sv2v_reg,mem_260_sv2v_reg,mem_259_sv2v_reg,
  mem_258_sv2v_reg,mem_257_sv2v_reg,mem_256_sv2v_reg,mem_255_sv2v_reg,mem_254_sv2v_reg,
  mem_253_sv2v_reg,mem_252_sv2v_reg,mem_251_sv2v_reg,mem_250_sv2v_reg,mem_249_sv2v_reg,
  mem_248_sv2v_reg,mem_247_sv2v_reg,mem_246_sv2v_reg,mem_245_sv2v_reg,
  mem_244_sv2v_reg,mem_243_sv2v_reg,mem_242_sv2v_reg,mem_241_sv2v_reg,mem_240_sv2v_reg,
  mem_239_sv2v_reg,mem_238_sv2v_reg,mem_237_sv2v_reg,mem_236_sv2v_reg,mem_235_sv2v_reg,
  mem_234_sv2v_reg,mem_233_sv2v_reg,mem_232_sv2v_reg,mem_231_sv2v_reg,
  mem_230_sv2v_reg,mem_229_sv2v_reg,mem_228_sv2v_reg,mem_227_sv2v_reg,mem_226_sv2v_reg,
  mem_225_sv2v_reg,mem_224_sv2v_reg,mem_223_sv2v_reg,mem_222_sv2v_reg,mem_221_sv2v_reg,
  mem_220_sv2v_reg,mem_219_sv2v_reg,mem_218_sv2v_reg,mem_217_sv2v_reg,mem_216_sv2v_reg,
  mem_215_sv2v_reg,mem_214_sv2v_reg,mem_213_sv2v_reg,mem_212_sv2v_reg,
  mem_211_sv2v_reg,mem_210_sv2v_reg,mem_209_sv2v_reg,mem_208_sv2v_reg,mem_207_sv2v_reg,
  mem_206_sv2v_reg,mem_205_sv2v_reg,mem_204_sv2v_reg,mem_203_sv2v_reg,mem_202_sv2v_reg,
  mem_201_sv2v_reg,mem_200_sv2v_reg,mem_199_sv2v_reg,mem_198_sv2v_reg,
  mem_197_sv2v_reg,mem_196_sv2v_reg,mem_195_sv2v_reg,mem_194_sv2v_reg,mem_193_sv2v_reg,
  mem_192_sv2v_reg,mem_191_sv2v_reg,mem_190_sv2v_reg,mem_189_sv2v_reg,mem_188_sv2v_reg,
  mem_187_sv2v_reg,mem_186_sv2v_reg,mem_185_sv2v_reg,mem_184_sv2v_reg,
  mem_183_sv2v_reg,mem_182_sv2v_reg,mem_181_sv2v_reg,mem_180_sv2v_reg,mem_179_sv2v_reg,
  mem_178_sv2v_reg,mem_177_sv2v_reg,mem_176_sv2v_reg,mem_175_sv2v_reg,mem_174_sv2v_reg,
  mem_173_sv2v_reg,mem_172_sv2v_reg,mem_171_sv2v_reg,mem_170_sv2v_reg,mem_169_sv2v_reg,
  mem_168_sv2v_reg,mem_167_sv2v_reg,mem_166_sv2v_reg,mem_165_sv2v_reg,
  mem_164_sv2v_reg,mem_163_sv2v_reg,mem_162_sv2v_reg,mem_161_sv2v_reg,mem_160_sv2v_reg,
  mem_159_sv2v_reg,mem_158_sv2v_reg,mem_157_sv2v_reg,mem_156_sv2v_reg,mem_155_sv2v_reg,
  mem_154_sv2v_reg,mem_153_sv2v_reg,mem_152_sv2v_reg,mem_151_sv2v_reg,
  mem_150_sv2v_reg,mem_149_sv2v_reg,mem_148_sv2v_reg,mem_147_sv2v_reg,mem_146_sv2v_reg,
  mem_145_sv2v_reg,mem_144_sv2v_reg,mem_143_sv2v_reg,mem_142_sv2v_reg,mem_141_sv2v_reg,
  mem_140_sv2v_reg,mem_139_sv2v_reg,mem_138_sv2v_reg,mem_137_sv2v_reg,mem_136_sv2v_reg,
  mem_135_sv2v_reg,mem_134_sv2v_reg,mem_133_sv2v_reg,mem_132_sv2v_reg,
  mem_131_sv2v_reg,mem_130_sv2v_reg,mem_129_sv2v_reg,mem_128_sv2v_reg,mem_127_sv2v_reg,
  mem_126_sv2v_reg,mem_125_sv2v_reg,mem_124_sv2v_reg,mem_123_sv2v_reg,mem_122_sv2v_reg,
  mem_121_sv2v_reg,mem_120_sv2v_reg,mem_119_sv2v_reg,mem_118_sv2v_reg,
  mem_117_sv2v_reg,mem_116_sv2v_reg,mem_115_sv2v_reg,mem_114_sv2v_reg,mem_113_sv2v_reg,
  mem_112_sv2v_reg,mem_111_sv2v_reg,mem_110_sv2v_reg,mem_109_sv2v_reg,mem_108_sv2v_reg,
  mem_107_sv2v_reg,mem_106_sv2v_reg,mem_105_sv2v_reg,mem_104_sv2v_reg,
  mem_103_sv2v_reg,mem_102_sv2v_reg,mem_101_sv2v_reg,mem_100_sv2v_reg,mem_99_sv2v_reg,
  mem_98_sv2v_reg,mem_97_sv2v_reg,mem_96_sv2v_reg,mem_95_sv2v_reg,mem_94_sv2v_reg,
  mem_93_sv2v_reg,mem_92_sv2v_reg,mem_91_sv2v_reg,mem_90_sv2v_reg,mem_89_sv2v_reg,
  mem_88_sv2v_reg,mem_87_sv2v_reg,mem_86_sv2v_reg,mem_85_sv2v_reg,mem_84_sv2v_reg,
  mem_83_sv2v_reg,mem_82_sv2v_reg,mem_81_sv2v_reg,mem_80_sv2v_reg,mem_79_sv2v_reg,
  mem_78_sv2v_reg,mem_77_sv2v_reg,mem_76_sv2v_reg,mem_75_sv2v_reg,mem_74_sv2v_reg,
  mem_73_sv2v_reg,mem_72_sv2v_reg,mem_71_sv2v_reg,mem_70_sv2v_reg,mem_69_sv2v_reg,
  mem_68_sv2v_reg,mem_67_sv2v_reg,mem_66_sv2v_reg,mem_65_sv2v_reg,mem_64_sv2v_reg,
  mem_63_sv2v_reg,mem_62_sv2v_reg,mem_61_sv2v_reg,mem_60_sv2v_reg,mem_59_sv2v_reg,
  mem_58_sv2v_reg,mem_57_sv2v_reg,mem_56_sv2v_reg,mem_55_sv2v_reg,mem_54_sv2v_reg,
  mem_53_sv2v_reg,mem_52_sv2v_reg,mem_51_sv2v_reg,mem_50_sv2v_reg,mem_49_sv2v_reg,
  mem_48_sv2v_reg,mem_47_sv2v_reg,mem_46_sv2v_reg,mem_45_sv2v_reg,mem_44_sv2v_reg,
  mem_43_sv2v_reg,mem_42_sv2v_reg,mem_41_sv2v_reg,mem_40_sv2v_reg,mem_39_sv2v_reg,
  mem_38_sv2v_reg,mem_37_sv2v_reg,mem_36_sv2v_reg,mem_35_sv2v_reg,mem_34_sv2v_reg,
  mem_33_sv2v_reg,mem_32_sv2v_reg,mem_31_sv2v_reg,mem_30_sv2v_reg,mem_29_sv2v_reg,
  mem_28_sv2v_reg,mem_27_sv2v_reg,mem_26_sv2v_reg,mem_25_sv2v_reg,mem_24_sv2v_reg,
  mem_23_sv2v_reg,mem_22_sv2v_reg,mem_21_sv2v_reg,mem_20_sv2v_reg,mem_19_sv2v_reg,
  mem_18_sv2v_reg,mem_17_sv2v_reg,mem_16_sv2v_reg,mem_15_sv2v_reg,mem_14_sv2v_reg,
  mem_13_sv2v_reg,mem_12_sv2v_reg,mem_11_sv2v_reg,mem_10_sv2v_reg,mem_9_sv2v_reg,
  mem_8_sv2v_reg,mem_7_sv2v_reg,mem_6_sv2v_reg,mem_5_sv2v_reg,mem_4_sv2v_reg,mem_3_sv2v_reg,
  mem_2_sv2v_reg,mem_1_sv2v_reg,mem_0_sv2v_reg;
  assign mem[1023] = mem_1023_sv2v_reg;
  assign mem[1022] = mem_1022_sv2v_reg;
  assign mem[1021] = mem_1021_sv2v_reg;
  assign mem[1020] = mem_1020_sv2v_reg;
  assign mem[1019] = mem_1019_sv2v_reg;
  assign mem[1018] = mem_1018_sv2v_reg;
  assign mem[1017] = mem_1017_sv2v_reg;
  assign mem[1016] = mem_1016_sv2v_reg;
  assign mem[1015] = mem_1015_sv2v_reg;
  assign mem[1014] = mem_1014_sv2v_reg;
  assign mem[1013] = mem_1013_sv2v_reg;
  assign mem[1012] = mem_1012_sv2v_reg;
  assign mem[1011] = mem_1011_sv2v_reg;
  assign mem[1010] = mem_1010_sv2v_reg;
  assign mem[1009] = mem_1009_sv2v_reg;
  assign mem[1008] = mem_1008_sv2v_reg;
  assign mem[1007] = mem_1007_sv2v_reg;
  assign mem[1006] = mem_1006_sv2v_reg;
  assign mem[1005] = mem_1005_sv2v_reg;
  assign mem[1004] = mem_1004_sv2v_reg;
  assign mem[1003] = mem_1003_sv2v_reg;
  assign mem[1002] = mem_1002_sv2v_reg;
  assign mem[1001] = mem_1001_sv2v_reg;
  assign mem[1000] = mem_1000_sv2v_reg;
  assign mem[999] = mem_999_sv2v_reg;
  assign mem[998] = mem_998_sv2v_reg;
  assign mem[997] = mem_997_sv2v_reg;
  assign mem[996] = mem_996_sv2v_reg;
  assign mem[995] = mem_995_sv2v_reg;
  assign mem[994] = mem_994_sv2v_reg;
  assign mem[993] = mem_993_sv2v_reg;
  assign mem[992] = mem_992_sv2v_reg;
  assign mem[991] = mem_991_sv2v_reg;
  assign mem[990] = mem_990_sv2v_reg;
  assign mem[989] = mem_989_sv2v_reg;
  assign mem[988] = mem_988_sv2v_reg;
  assign mem[987] = mem_987_sv2v_reg;
  assign mem[986] = mem_986_sv2v_reg;
  assign mem[985] = mem_985_sv2v_reg;
  assign mem[984] = mem_984_sv2v_reg;
  assign mem[983] = mem_983_sv2v_reg;
  assign mem[982] = mem_982_sv2v_reg;
  assign mem[981] = mem_981_sv2v_reg;
  assign mem[980] = mem_980_sv2v_reg;
  assign mem[979] = mem_979_sv2v_reg;
  assign mem[978] = mem_978_sv2v_reg;
  assign mem[977] = mem_977_sv2v_reg;
  assign mem[976] = mem_976_sv2v_reg;
  assign mem[975] = mem_975_sv2v_reg;
  assign mem[974] = mem_974_sv2v_reg;
  assign mem[973] = mem_973_sv2v_reg;
  assign mem[972] = mem_972_sv2v_reg;
  assign mem[971] = mem_971_sv2v_reg;
  assign mem[970] = mem_970_sv2v_reg;
  assign mem[969] = mem_969_sv2v_reg;
  assign mem[968] = mem_968_sv2v_reg;
  assign mem[967] = mem_967_sv2v_reg;
  assign mem[966] = mem_966_sv2v_reg;
  assign mem[965] = mem_965_sv2v_reg;
  assign mem[964] = mem_964_sv2v_reg;
  assign mem[963] = mem_963_sv2v_reg;
  assign mem[962] = mem_962_sv2v_reg;
  assign mem[961] = mem_961_sv2v_reg;
  assign mem[960] = mem_960_sv2v_reg;
  assign mem[959] = mem_959_sv2v_reg;
  assign mem[958] = mem_958_sv2v_reg;
  assign mem[957] = mem_957_sv2v_reg;
  assign mem[956] = mem_956_sv2v_reg;
  assign mem[955] = mem_955_sv2v_reg;
  assign mem[954] = mem_954_sv2v_reg;
  assign mem[953] = mem_953_sv2v_reg;
  assign mem[952] = mem_952_sv2v_reg;
  assign mem[951] = mem_951_sv2v_reg;
  assign mem[950] = mem_950_sv2v_reg;
  assign mem[949] = mem_949_sv2v_reg;
  assign mem[948] = mem_948_sv2v_reg;
  assign mem[947] = mem_947_sv2v_reg;
  assign mem[946] = mem_946_sv2v_reg;
  assign mem[945] = mem_945_sv2v_reg;
  assign mem[944] = mem_944_sv2v_reg;
  assign mem[943] = mem_943_sv2v_reg;
  assign mem[942] = mem_942_sv2v_reg;
  assign mem[941] = mem_941_sv2v_reg;
  assign mem[940] = mem_940_sv2v_reg;
  assign mem[939] = mem_939_sv2v_reg;
  assign mem[938] = mem_938_sv2v_reg;
  assign mem[937] = mem_937_sv2v_reg;
  assign mem[936] = mem_936_sv2v_reg;
  assign mem[935] = mem_935_sv2v_reg;
  assign mem[934] = mem_934_sv2v_reg;
  assign mem[933] = mem_933_sv2v_reg;
  assign mem[932] = mem_932_sv2v_reg;
  assign mem[931] = mem_931_sv2v_reg;
  assign mem[930] = mem_930_sv2v_reg;
  assign mem[929] = mem_929_sv2v_reg;
  assign mem[928] = mem_928_sv2v_reg;
  assign mem[927] = mem_927_sv2v_reg;
  assign mem[926] = mem_926_sv2v_reg;
  assign mem[925] = mem_925_sv2v_reg;
  assign mem[924] = mem_924_sv2v_reg;
  assign mem[923] = mem_923_sv2v_reg;
  assign mem[922] = mem_922_sv2v_reg;
  assign mem[921] = mem_921_sv2v_reg;
  assign mem[920] = mem_920_sv2v_reg;
  assign mem[919] = mem_919_sv2v_reg;
  assign mem[918] = mem_918_sv2v_reg;
  assign mem[917] = mem_917_sv2v_reg;
  assign mem[916] = mem_916_sv2v_reg;
  assign mem[915] = mem_915_sv2v_reg;
  assign mem[914] = mem_914_sv2v_reg;
  assign mem[913] = mem_913_sv2v_reg;
  assign mem[912] = mem_912_sv2v_reg;
  assign mem[911] = mem_911_sv2v_reg;
  assign mem[910] = mem_910_sv2v_reg;
  assign mem[909] = mem_909_sv2v_reg;
  assign mem[908] = mem_908_sv2v_reg;
  assign mem[907] = mem_907_sv2v_reg;
  assign mem[906] = mem_906_sv2v_reg;
  assign mem[905] = mem_905_sv2v_reg;
  assign mem[904] = mem_904_sv2v_reg;
  assign mem[903] = mem_903_sv2v_reg;
  assign mem[902] = mem_902_sv2v_reg;
  assign mem[901] = mem_901_sv2v_reg;
  assign mem[900] = mem_900_sv2v_reg;
  assign mem[899] = mem_899_sv2v_reg;
  assign mem[898] = mem_898_sv2v_reg;
  assign mem[897] = mem_897_sv2v_reg;
  assign mem[896] = mem_896_sv2v_reg;
  assign mem[895] = mem_895_sv2v_reg;
  assign mem[894] = mem_894_sv2v_reg;
  assign mem[893] = mem_893_sv2v_reg;
  assign mem[892] = mem_892_sv2v_reg;
  assign mem[891] = mem_891_sv2v_reg;
  assign mem[890] = mem_890_sv2v_reg;
  assign mem[889] = mem_889_sv2v_reg;
  assign mem[888] = mem_888_sv2v_reg;
  assign mem[887] = mem_887_sv2v_reg;
  assign mem[886] = mem_886_sv2v_reg;
  assign mem[885] = mem_885_sv2v_reg;
  assign mem[884] = mem_884_sv2v_reg;
  assign mem[883] = mem_883_sv2v_reg;
  assign mem[882] = mem_882_sv2v_reg;
  assign mem[881] = mem_881_sv2v_reg;
  assign mem[880] = mem_880_sv2v_reg;
  assign mem[879] = mem_879_sv2v_reg;
  assign mem[878] = mem_878_sv2v_reg;
  assign mem[877] = mem_877_sv2v_reg;
  assign mem[876] = mem_876_sv2v_reg;
  assign mem[875] = mem_875_sv2v_reg;
  assign mem[874] = mem_874_sv2v_reg;
  assign mem[873] = mem_873_sv2v_reg;
  assign mem[872] = mem_872_sv2v_reg;
  assign mem[871] = mem_871_sv2v_reg;
  assign mem[870] = mem_870_sv2v_reg;
  assign mem[869] = mem_869_sv2v_reg;
  assign mem[868] = mem_868_sv2v_reg;
  assign mem[867] = mem_867_sv2v_reg;
  assign mem[866] = mem_866_sv2v_reg;
  assign mem[865] = mem_865_sv2v_reg;
  assign mem[864] = mem_864_sv2v_reg;
  assign mem[863] = mem_863_sv2v_reg;
  assign mem[862] = mem_862_sv2v_reg;
  assign mem[861] = mem_861_sv2v_reg;
  assign mem[860] = mem_860_sv2v_reg;
  assign mem[859] = mem_859_sv2v_reg;
  assign mem[858] = mem_858_sv2v_reg;
  assign mem[857] = mem_857_sv2v_reg;
  assign mem[856] = mem_856_sv2v_reg;
  assign mem[855] = mem_855_sv2v_reg;
  assign mem[854] = mem_854_sv2v_reg;
  assign mem[853] = mem_853_sv2v_reg;
  assign mem[852] = mem_852_sv2v_reg;
  assign mem[851] = mem_851_sv2v_reg;
  assign mem[850] = mem_850_sv2v_reg;
  assign mem[849] = mem_849_sv2v_reg;
  assign mem[848] = mem_848_sv2v_reg;
  assign mem[847] = mem_847_sv2v_reg;
  assign mem[846] = mem_846_sv2v_reg;
  assign mem[845] = mem_845_sv2v_reg;
  assign mem[844] = mem_844_sv2v_reg;
  assign mem[843] = mem_843_sv2v_reg;
  assign mem[842] = mem_842_sv2v_reg;
  assign mem[841] = mem_841_sv2v_reg;
  assign mem[840] = mem_840_sv2v_reg;
  assign mem[839] = mem_839_sv2v_reg;
  assign mem[838] = mem_838_sv2v_reg;
  assign mem[837] = mem_837_sv2v_reg;
  assign mem[836] = mem_836_sv2v_reg;
  assign mem[835] = mem_835_sv2v_reg;
  assign mem[834] = mem_834_sv2v_reg;
  assign mem[833] = mem_833_sv2v_reg;
  assign mem[832] = mem_832_sv2v_reg;
  assign mem[831] = mem_831_sv2v_reg;
  assign mem[830] = mem_830_sv2v_reg;
  assign mem[829] = mem_829_sv2v_reg;
  assign mem[828] = mem_828_sv2v_reg;
  assign mem[827] = mem_827_sv2v_reg;
  assign mem[826] = mem_826_sv2v_reg;
  assign mem[825] = mem_825_sv2v_reg;
  assign mem[824] = mem_824_sv2v_reg;
  assign mem[823] = mem_823_sv2v_reg;
  assign mem[822] = mem_822_sv2v_reg;
  assign mem[821] = mem_821_sv2v_reg;
  assign mem[820] = mem_820_sv2v_reg;
  assign mem[819] = mem_819_sv2v_reg;
  assign mem[818] = mem_818_sv2v_reg;
  assign mem[817] = mem_817_sv2v_reg;
  assign mem[816] = mem_816_sv2v_reg;
  assign mem[815] = mem_815_sv2v_reg;
  assign mem[814] = mem_814_sv2v_reg;
  assign mem[813] = mem_813_sv2v_reg;
  assign mem[812] = mem_812_sv2v_reg;
  assign mem[811] = mem_811_sv2v_reg;
  assign mem[810] = mem_810_sv2v_reg;
  assign mem[809] = mem_809_sv2v_reg;
  assign mem[808] = mem_808_sv2v_reg;
  assign mem[807] = mem_807_sv2v_reg;
  assign mem[806] = mem_806_sv2v_reg;
  assign mem[805] = mem_805_sv2v_reg;
  assign mem[804] = mem_804_sv2v_reg;
  assign mem[803] = mem_803_sv2v_reg;
  assign mem[802] = mem_802_sv2v_reg;
  assign mem[801] = mem_801_sv2v_reg;
  assign mem[800] = mem_800_sv2v_reg;
  assign mem[799] = mem_799_sv2v_reg;
  assign mem[798] = mem_798_sv2v_reg;
  assign mem[797] = mem_797_sv2v_reg;
  assign mem[796] = mem_796_sv2v_reg;
  assign mem[795] = mem_795_sv2v_reg;
  assign mem[794] = mem_794_sv2v_reg;
  assign mem[793] = mem_793_sv2v_reg;
  assign mem[792] = mem_792_sv2v_reg;
  assign mem[791] = mem_791_sv2v_reg;
  assign mem[790] = mem_790_sv2v_reg;
  assign mem[789] = mem_789_sv2v_reg;
  assign mem[788] = mem_788_sv2v_reg;
  assign mem[787] = mem_787_sv2v_reg;
  assign mem[786] = mem_786_sv2v_reg;
  assign mem[785] = mem_785_sv2v_reg;
  assign mem[784] = mem_784_sv2v_reg;
  assign mem[783] = mem_783_sv2v_reg;
  assign mem[782] = mem_782_sv2v_reg;
  assign mem[781] = mem_781_sv2v_reg;
  assign mem[780] = mem_780_sv2v_reg;
  assign mem[779] = mem_779_sv2v_reg;
  assign mem[778] = mem_778_sv2v_reg;
  assign mem[777] = mem_777_sv2v_reg;
  assign mem[776] = mem_776_sv2v_reg;
  assign mem[775] = mem_775_sv2v_reg;
  assign mem[774] = mem_774_sv2v_reg;
  assign mem[773] = mem_773_sv2v_reg;
  assign mem[772] = mem_772_sv2v_reg;
  assign mem[771] = mem_771_sv2v_reg;
  assign mem[770] = mem_770_sv2v_reg;
  assign mem[769] = mem_769_sv2v_reg;
  assign mem[768] = mem_768_sv2v_reg;
  assign mem[767] = mem_767_sv2v_reg;
  assign mem[766] = mem_766_sv2v_reg;
  assign mem[765] = mem_765_sv2v_reg;
  assign mem[764] = mem_764_sv2v_reg;
  assign mem[763] = mem_763_sv2v_reg;
  assign mem[762] = mem_762_sv2v_reg;
  assign mem[761] = mem_761_sv2v_reg;
  assign mem[760] = mem_760_sv2v_reg;
  assign mem[759] = mem_759_sv2v_reg;
  assign mem[758] = mem_758_sv2v_reg;
  assign mem[757] = mem_757_sv2v_reg;
  assign mem[756] = mem_756_sv2v_reg;
  assign mem[755] = mem_755_sv2v_reg;
  assign mem[754] = mem_754_sv2v_reg;
  assign mem[753] = mem_753_sv2v_reg;
  assign mem[752] = mem_752_sv2v_reg;
  assign mem[751] = mem_751_sv2v_reg;
  assign mem[750] = mem_750_sv2v_reg;
  assign mem[749] = mem_749_sv2v_reg;
  assign mem[748] = mem_748_sv2v_reg;
  assign mem[747] = mem_747_sv2v_reg;
  assign mem[746] = mem_746_sv2v_reg;
  assign mem[745] = mem_745_sv2v_reg;
  assign mem[744] = mem_744_sv2v_reg;
  assign mem[743] = mem_743_sv2v_reg;
  assign mem[742] = mem_742_sv2v_reg;
  assign mem[741] = mem_741_sv2v_reg;
  assign mem[740] = mem_740_sv2v_reg;
  assign mem[739] = mem_739_sv2v_reg;
  assign mem[738] = mem_738_sv2v_reg;
  assign mem[737] = mem_737_sv2v_reg;
  assign mem[736] = mem_736_sv2v_reg;
  assign mem[735] = mem_735_sv2v_reg;
  assign mem[734] = mem_734_sv2v_reg;
  assign mem[733] = mem_733_sv2v_reg;
  assign mem[732] = mem_732_sv2v_reg;
  assign mem[731] = mem_731_sv2v_reg;
  assign mem[730] = mem_730_sv2v_reg;
  assign mem[729] = mem_729_sv2v_reg;
  assign mem[728] = mem_728_sv2v_reg;
  assign mem[727] = mem_727_sv2v_reg;
  assign mem[726] = mem_726_sv2v_reg;
  assign mem[725] = mem_725_sv2v_reg;
  assign mem[724] = mem_724_sv2v_reg;
  assign mem[723] = mem_723_sv2v_reg;
  assign mem[722] = mem_722_sv2v_reg;
  assign mem[721] = mem_721_sv2v_reg;
  assign mem[720] = mem_720_sv2v_reg;
  assign mem[719] = mem_719_sv2v_reg;
  assign mem[718] = mem_718_sv2v_reg;
  assign mem[717] = mem_717_sv2v_reg;
  assign mem[716] = mem_716_sv2v_reg;
  assign mem[715] = mem_715_sv2v_reg;
  assign mem[714] = mem_714_sv2v_reg;
  assign mem[713] = mem_713_sv2v_reg;
  assign mem[712] = mem_712_sv2v_reg;
  assign mem[711] = mem_711_sv2v_reg;
  assign mem[710] = mem_710_sv2v_reg;
  assign mem[709] = mem_709_sv2v_reg;
  assign mem[708] = mem_708_sv2v_reg;
  assign mem[707] = mem_707_sv2v_reg;
  assign mem[706] = mem_706_sv2v_reg;
  assign mem[705] = mem_705_sv2v_reg;
  assign mem[704] = mem_704_sv2v_reg;
  assign mem[703] = mem_703_sv2v_reg;
  assign mem[702] = mem_702_sv2v_reg;
  assign mem[701] = mem_701_sv2v_reg;
  assign mem[700] = mem_700_sv2v_reg;
  assign mem[699] = mem_699_sv2v_reg;
  assign mem[698] = mem_698_sv2v_reg;
  assign mem[697] = mem_697_sv2v_reg;
  assign mem[696] = mem_696_sv2v_reg;
  assign mem[695] = mem_695_sv2v_reg;
  assign mem[694] = mem_694_sv2v_reg;
  assign mem[693] = mem_693_sv2v_reg;
  assign mem[692] = mem_692_sv2v_reg;
  assign mem[691] = mem_691_sv2v_reg;
  assign mem[690] = mem_690_sv2v_reg;
  assign mem[689] = mem_689_sv2v_reg;
  assign mem[688] = mem_688_sv2v_reg;
  assign mem[687] = mem_687_sv2v_reg;
  assign mem[686] = mem_686_sv2v_reg;
  assign mem[685] = mem_685_sv2v_reg;
  assign mem[684] = mem_684_sv2v_reg;
  assign mem[683] = mem_683_sv2v_reg;
  assign mem[682] = mem_682_sv2v_reg;
  assign mem[681] = mem_681_sv2v_reg;
  assign mem[680] = mem_680_sv2v_reg;
  assign mem[679] = mem_679_sv2v_reg;
  assign mem[678] = mem_678_sv2v_reg;
  assign mem[677] = mem_677_sv2v_reg;
  assign mem[676] = mem_676_sv2v_reg;
  assign mem[675] = mem_675_sv2v_reg;
  assign mem[674] = mem_674_sv2v_reg;
  assign mem[673] = mem_673_sv2v_reg;
  assign mem[672] = mem_672_sv2v_reg;
  assign mem[671] = mem_671_sv2v_reg;
  assign mem[670] = mem_670_sv2v_reg;
  assign mem[669] = mem_669_sv2v_reg;
  assign mem[668] = mem_668_sv2v_reg;
  assign mem[667] = mem_667_sv2v_reg;
  assign mem[666] = mem_666_sv2v_reg;
  assign mem[665] = mem_665_sv2v_reg;
  assign mem[664] = mem_664_sv2v_reg;
  assign mem[663] = mem_663_sv2v_reg;
  assign mem[662] = mem_662_sv2v_reg;
  assign mem[661] = mem_661_sv2v_reg;
  assign mem[660] = mem_660_sv2v_reg;
  assign mem[659] = mem_659_sv2v_reg;
  assign mem[658] = mem_658_sv2v_reg;
  assign mem[657] = mem_657_sv2v_reg;
  assign mem[656] = mem_656_sv2v_reg;
  assign mem[655] = mem_655_sv2v_reg;
  assign mem[654] = mem_654_sv2v_reg;
  assign mem[653] = mem_653_sv2v_reg;
  assign mem[652] = mem_652_sv2v_reg;
  assign mem[651] = mem_651_sv2v_reg;
  assign mem[650] = mem_650_sv2v_reg;
  assign mem[649] = mem_649_sv2v_reg;
  assign mem[648] = mem_648_sv2v_reg;
  assign mem[647] = mem_647_sv2v_reg;
  assign mem[646] = mem_646_sv2v_reg;
  assign mem[645] = mem_645_sv2v_reg;
  assign mem[644] = mem_644_sv2v_reg;
  assign mem[643] = mem_643_sv2v_reg;
  assign mem[642] = mem_642_sv2v_reg;
  assign mem[641] = mem_641_sv2v_reg;
  assign mem[640] = mem_640_sv2v_reg;
  assign mem[639] = mem_639_sv2v_reg;
  assign mem[638] = mem_638_sv2v_reg;
  assign mem[637] = mem_637_sv2v_reg;
  assign mem[636] = mem_636_sv2v_reg;
  assign mem[635] = mem_635_sv2v_reg;
  assign mem[634] = mem_634_sv2v_reg;
  assign mem[633] = mem_633_sv2v_reg;
  assign mem[632] = mem_632_sv2v_reg;
  assign mem[631] = mem_631_sv2v_reg;
  assign mem[630] = mem_630_sv2v_reg;
  assign mem[629] = mem_629_sv2v_reg;
  assign mem[628] = mem_628_sv2v_reg;
  assign mem[627] = mem_627_sv2v_reg;
  assign mem[626] = mem_626_sv2v_reg;
  assign mem[625] = mem_625_sv2v_reg;
  assign mem[624] = mem_624_sv2v_reg;
  assign mem[623] = mem_623_sv2v_reg;
  assign mem[622] = mem_622_sv2v_reg;
  assign mem[621] = mem_621_sv2v_reg;
  assign mem[620] = mem_620_sv2v_reg;
  assign mem[619] = mem_619_sv2v_reg;
  assign mem[618] = mem_618_sv2v_reg;
  assign mem[617] = mem_617_sv2v_reg;
  assign mem[616] = mem_616_sv2v_reg;
  assign mem[615] = mem_615_sv2v_reg;
  assign mem[614] = mem_614_sv2v_reg;
  assign mem[613] = mem_613_sv2v_reg;
  assign mem[612] = mem_612_sv2v_reg;
  assign mem[611] = mem_611_sv2v_reg;
  assign mem[610] = mem_610_sv2v_reg;
  assign mem[609] = mem_609_sv2v_reg;
  assign mem[608] = mem_608_sv2v_reg;
  assign mem[607] = mem_607_sv2v_reg;
  assign mem[606] = mem_606_sv2v_reg;
  assign mem[605] = mem_605_sv2v_reg;
  assign mem[604] = mem_604_sv2v_reg;
  assign mem[603] = mem_603_sv2v_reg;
  assign mem[602] = mem_602_sv2v_reg;
  assign mem[601] = mem_601_sv2v_reg;
  assign mem[600] = mem_600_sv2v_reg;
  assign mem[599] = mem_599_sv2v_reg;
  assign mem[598] = mem_598_sv2v_reg;
  assign mem[597] = mem_597_sv2v_reg;
  assign mem[596] = mem_596_sv2v_reg;
  assign mem[595] = mem_595_sv2v_reg;
  assign mem[594] = mem_594_sv2v_reg;
  assign mem[593] = mem_593_sv2v_reg;
  assign mem[592] = mem_592_sv2v_reg;
  assign mem[591] = mem_591_sv2v_reg;
  assign mem[590] = mem_590_sv2v_reg;
  assign mem[589] = mem_589_sv2v_reg;
  assign mem[588] = mem_588_sv2v_reg;
  assign mem[587] = mem_587_sv2v_reg;
  assign mem[586] = mem_586_sv2v_reg;
  assign mem[585] = mem_585_sv2v_reg;
  assign mem[584] = mem_584_sv2v_reg;
  assign mem[583] = mem_583_sv2v_reg;
  assign mem[582] = mem_582_sv2v_reg;
  assign mem[581] = mem_581_sv2v_reg;
  assign mem[580] = mem_580_sv2v_reg;
  assign mem[579] = mem_579_sv2v_reg;
  assign mem[578] = mem_578_sv2v_reg;
  assign mem[577] = mem_577_sv2v_reg;
  assign mem[576] = mem_576_sv2v_reg;
  assign mem[575] = mem_575_sv2v_reg;
  assign mem[574] = mem_574_sv2v_reg;
  assign mem[573] = mem_573_sv2v_reg;
  assign mem[572] = mem_572_sv2v_reg;
  assign mem[571] = mem_571_sv2v_reg;
  assign mem[570] = mem_570_sv2v_reg;
  assign mem[569] = mem_569_sv2v_reg;
  assign mem[568] = mem_568_sv2v_reg;
  assign mem[567] = mem_567_sv2v_reg;
  assign mem[566] = mem_566_sv2v_reg;
  assign mem[565] = mem_565_sv2v_reg;
  assign mem[564] = mem_564_sv2v_reg;
  assign mem[563] = mem_563_sv2v_reg;
  assign mem[562] = mem_562_sv2v_reg;
  assign mem[561] = mem_561_sv2v_reg;
  assign mem[560] = mem_560_sv2v_reg;
  assign mem[559] = mem_559_sv2v_reg;
  assign mem[558] = mem_558_sv2v_reg;
  assign mem[557] = mem_557_sv2v_reg;
  assign mem[556] = mem_556_sv2v_reg;
  assign mem[555] = mem_555_sv2v_reg;
  assign mem[554] = mem_554_sv2v_reg;
  assign mem[553] = mem_553_sv2v_reg;
  assign mem[552] = mem_552_sv2v_reg;
  assign mem[551] = mem_551_sv2v_reg;
  assign mem[550] = mem_550_sv2v_reg;
  assign mem[549] = mem_549_sv2v_reg;
  assign mem[548] = mem_548_sv2v_reg;
  assign mem[547] = mem_547_sv2v_reg;
  assign mem[546] = mem_546_sv2v_reg;
  assign mem[545] = mem_545_sv2v_reg;
  assign mem[544] = mem_544_sv2v_reg;
  assign mem[543] = mem_543_sv2v_reg;
  assign mem[542] = mem_542_sv2v_reg;
  assign mem[541] = mem_541_sv2v_reg;
  assign mem[540] = mem_540_sv2v_reg;
  assign mem[539] = mem_539_sv2v_reg;
  assign mem[538] = mem_538_sv2v_reg;
  assign mem[537] = mem_537_sv2v_reg;
  assign mem[536] = mem_536_sv2v_reg;
  assign mem[535] = mem_535_sv2v_reg;
  assign mem[534] = mem_534_sv2v_reg;
  assign mem[533] = mem_533_sv2v_reg;
  assign mem[532] = mem_532_sv2v_reg;
  assign mem[531] = mem_531_sv2v_reg;
  assign mem[530] = mem_530_sv2v_reg;
  assign mem[529] = mem_529_sv2v_reg;
  assign mem[528] = mem_528_sv2v_reg;
  assign mem[527] = mem_527_sv2v_reg;
  assign mem[526] = mem_526_sv2v_reg;
  assign mem[525] = mem_525_sv2v_reg;
  assign mem[524] = mem_524_sv2v_reg;
  assign mem[523] = mem_523_sv2v_reg;
  assign mem[522] = mem_522_sv2v_reg;
  assign mem[521] = mem_521_sv2v_reg;
  assign mem[520] = mem_520_sv2v_reg;
  assign mem[519] = mem_519_sv2v_reg;
  assign mem[518] = mem_518_sv2v_reg;
  assign mem[517] = mem_517_sv2v_reg;
  assign mem[516] = mem_516_sv2v_reg;
  assign mem[515] = mem_515_sv2v_reg;
  assign mem[514] = mem_514_sv2v_reg;
  assign mem[513] = mem_513_sv2v_reg;
  assign mem[512] = mem_512_sv2v_reg;
  assign mem[511] = mem_511_sv2v_reg;
  assign mem[510] = mem_510_sv2v_reg;
  assign mem[509] = mem_509_sv2v_reg;
  assign mem[508] = mem_508_sv2v_reg;
  assign mem[507] = mem_507_sv2v_reg;
  assign mem[506] = mem_506_sv2v_reg;
  assign mem[505] = mem_505_sv2v_reg;
  assign mem[504] = mem_504_sv2v_reg;
  assign mem[503] = mem_503_sv2v_reg;
  assign mem[502] = mem_502_sv2v_reg;
  assign mem[501] = mem_501_sv2v_reg;
  assign mem[500] = mem_500_sv2v_reg;
  assign mem[499] = mem_499_sv2v_reg;
  assign mem[498] = mem_498_sv2v_reg;
  assign mem[497] = mem_497_sv2v_reg;
  assign mem[496] = mem_496_sv2v_reg;
  assign mem[495] = mem_495_sv2v_reg;
  assign mem[494] = mem_494_sv2v_reg;
  assign mem[493] = mem_493_sv2v_reg;
  assign mem[492] = mem_492_sv2v_reg;
  assign mem[491] = mem_491_sv2v_reg;
  assign mem[490] = mem_490_sv2v_reg;
  assign mem[489] = mem_489_sv2v_reg;
  assign mem[488] = mem_488_sv2v_reg;
  assign mem[487] = mem_487_sv2v_reg;
  assign mem[486] = mem_486_sv2v_reg;
  assign mem[485] = mem_485_sv2v_reg;
  assign mem[484] = mem_484_sv2v_reg;
  assign mem[483] = mem_483_sv2v_reg;
  assign mem[482] = mem_482_sv2v_reg;
  assign mem[481] = mem_481_sv2v_reg;
  assign mem[480] = mem_480_sv2v_reg;
  assign mem[479] = mem_479_sv2v_reg;
  assign mem[478] = mem_478_sv2v_reg;
  assign mem[477] = mem_477_sv2v_reg;
  assign mem[476] = mem_476_sv2v_reg;
  assign mem[475] = mem_475_sv2v_reg;
  assign mem[474] = mem_474_sv2v_reg;
  assign mem[473] = mem_473_sv2v_reg;
  assign mem[472] = mem_472_sv2v_reg;
  assign mem[471] = mem_471_sv2v_reg;
  assign mem[470] = mem_470_sv2v_reg;
  assign mem[469] = mem_469_sv2v_reg;
  assign mem[468] = mem_468_sv2v_reg;
  assign mem[467] = mem_467_sv2v_reg;
  assign mem[466] = mem_466_sv2v_reg;
  assign mem[465] = mem_465_sv2v_reg;
  assign mem[464] = mem_464_sv2v_reg;
  assign mem[463] = mem_463_sv2v_reg;
  assign mem[462] = mem_462_sv2v_reg;
  assign mem[461] = mem_461_sv2v_reg;
  assign mem[460] = mem_460_sv2v_reg;
  assign mem[459] = mem_459_sv2v_reg;
  assign mem[458] = mem_458_sv2v_reg;
  assign mem[457] = mem_457_sv2v_reg;
  assign mem[456] = mem_456_sv2v_reg;
  assign mem[455] = mem_455_sv2v_reg;
  assign mem[454] = mem_454_sv2v_reg;
  assign mem[453] = mem_453_sv2v_reg;
  assign mem[452] = mem_452_sv2v_reg;
  assign mem[451] = mem_451_sv2v_reg;
  assign mem[450] = mem_450_sv2v_reg;
  assign mem[449] = mem_449_sv2v_reg;
  assign mem[448] = mem_448_sv2v_reg;
  assign mem[447] = mem_447_sv2v_reg;
  assign mem[446] = mem_446_sv2v_reg;
  assign mem[445] = mem_445_sv2v_reg;
  assign mem[444] = mem_444_sv2v_reg;
  assign mem[443] = mem_443_sv2v_reg;
  assign mem[442] = mem_442_sv2v_reg;
  assign mem[441] = mem_441_sv2v_reg;
  assign mem[440] = mem_440_sv2v_reg;
  assign mem[439] = mem_439_sv2v_reg;
  assign mem[438] = mem_438_sv2v_reg;
  assign mem[437] = mem_437_sv2v_reg;
  assign mem[436] = mem_436_sv2v_reg;
  assign mem[435] = mem_435_sv2v_reg;
  assign mem[434] = mem_434_sv2v_reg;
  assign mem[433] = mem_433_sv2v_reg;
  assign mem[432] = mem_432_sv2v_reg;
  assign mem[431] = mem_431_sv2v_reg;
  assign mem[430] = mem_430_sv2v_reg;
  assign mem[429] = mem_429_sv2v_reg;
  assign mem[428] = mem_428_sv2v_reg;
  assign mem[427] = mem_427_sv2v_reg;
  assign mem[426] = mem_426_sv2v_reg;
  assign mem[425] = mem_425_sv2v_reg;
  assign mem[424] = mem_424_sv2v_reg;
  assign mem[423] = mem_423_sv2v_reg;
  assign mem[422] = mem_422_sv2v_reg;
  assign mem[421] = mem_421_sv2v_reg;
  assign mem[420] = mem_420_sv2v_reg;
  assign mem[419] = mem_419_sv2v_reg;
  assign mem[418] = mem_418_sv2v_reg;
  assign mem[417] = mem_417_sv2v_reg;
  assign mem[416] = mem_416_sv2v_reg;
  assign mem[415] = mem_415_sv2v_reg;
  assign mem[414] = mem_414_sv2v_reg;
  assign mem[413] = mem_413_sv2v_reg;
  assign mem[412] = mem_412_sv2v_reg;
  assign mem[411] = mem_411_sv2v_reg;
  assign mem[410] = mem_410_sv2v_reg;
  assign mem[409] = mem_409_sv2v_reg;
  assign mem[408] = mem_408_sv2v_reg;
  assign mem[407] = mem_407_sv2v_reg;
  assign mem[406] = mem_406_sv2v_reg;
  assign mem[405] = mem_405_sv2v_reg;
  assign mem[404] = mem_404_sv2v_reg;
  assign mem[403] = mem_403_sv2v_reg;
  assign mem[402] = mem_402_sv2v_reg;
  assign mem[401] = mem_401_sv2v_reg;
  assign mem[400] = mem_400_sv2v_reg;
  assign mem[399] = mem_399_sv2v_reg;
  assign mem[398] = mem_398_sv2v_reg;
  assign mem[397] = mem_397_sv2v_reg;
  assign mem[396] = mem_396_sv2v_reg;
  assign mem[395] = mem_395_sv2v_reg;
  assign mem[394] = mem_394_sv2v_reg;
  assign mem[393] = mem_393_sv2v_reg;
  assign mem[392] = mem_392_sv2v_reg;
  assign mem[391] = mem_391_sv2v_reg;
  assign mem[390] = mem_390_sv2v_reg;
  assign mem[389] = mem_389_sv2v_reg;
  assign mem[388] = mem_388_sv2v_reg;
  assign mem[387] = mem_387_sv2v_reg;
  assign mem[386] = mem_386_sv2v_reg;
  assign mem[385] = mem_385_sv2v_reg;
  assign mem[384] = mem_384_sv2v_reg;
  assign mem[383] = mem_383_sv2v_reg;
  assign mem[382] = mem_382_sv2v_reg;
  assign mem[381] = mem_381_sv2v_reg;
  assign mem[380] = mem_380_sv2v_reg;
  assign mem[379] = mem_379_sv2v_reg;
  assign mem[378] = mem_378_sv2v_reg;
  assign mem[377] = mem_377_sv2v_reg;
  assign mem[376] = mem_376_sv2v_reg;
  assign mem[375] = mem_375_sv2v_reg;
  assign mem[374] = mem_374_sv2v_reg;
  assign mem[373] = mem_373_sv2v_reg;
  assign mem[372] = mem_372_sv2v_reg;
  assign mem[371] = mem_371_sv2v_reg;
  assign mem[370] = mem_370_sv2v_reg;
  assign mem[369] = mem_369_sv2v_reg;
  assign mem[368] = mem_368_sv2v_reg;
  assign mem[367] = mem_367_sv2v_reg;
  assign mem[366] = mem_366_sv2v_reg;
  assign mem[365] = mem_365_sv2v_reg;
  assign mem[364] = mem_364_sv2v_reg;
  assign mem[363] = mem_363_sv2v_reg;
  assign mem[362] = mem_362_sv2v_reg;
  assign mem[361] = mem_361_sv2v_reg;
  assign mem[360] = mem_360_sv2v_reg;
  assign mem[359] = mem_359_sv2v_reg;
  assign mem[358] = mem_358_sv2v_reg;
  assign mem[357] = mem_357_sv2v_reg;
  assign mem[356] = mem_356_sv2v_reg;
  assign mem[355] = mem_355_sv2v_reg;
  assign mem[354] = mem_354_sv2v_reg;
  assign mem[353] = mem_353_sv2v_reg;
  assign mem[352] = mem_352_sv2v_reg;
  assign mem[351] = mem_351_sv2v_reg;
  assign mem[350] = mem_350_sv2v_reg;
  assign mem[349] = mem_349_sv2v_reg;
  assign mem[348] = mem_348_sv2v_reg;
  assign mem[347] = mem_347_sv2v_reg;
  assign mem[346] = mem_346_sv2v_reg;
  assign mem[345] = mem_345_sv2v_reg;
  assign mem[344] = mem_344_sv2v_reg;
  assign mem[343] = mem_343_sv2v_reg;
  assign mem[342] = mem_342_sv2v_reg;
  assign mem[341] = mem_341_sv2v_reg;
  assign mem[340] = mem_340_sv2v_reg;
  assign mem[339] = mem_339_sv2v_reg;
  assign mem[338] = mem_338_sv2v_reg;
  assign mem[337] = mem_337_sv2v_reg;
  assign mem[336] = mem_336_sv2v_reg;
  assign mem[335] = mem_335_sv2v_reg;
  assign mem[334] = mem_334_sv2v_reg;
  assign mem[333] = mem_333_sv2v_reg;
  assign mem[332] = mem_332_sv2v_reg;
  assign mem[331] = mem_331_sv2v_reg;
  assign mem[330] = mem_330_sv2v_reg;
  assign mem[329] = mem_329_sv2v_reg;
  assign mem[328] = mem_328_sv2v_reg;
  assign mem[327] = mem_327_sv2v_reg;
  assign mem[326] = mem_326_sv2v_reg;
  assign mem[325] = mem_325_sv2v_reg;
  assign mem[324] = mem_324_sv2v_reg;
  assign mem[323] = mem_323_sv2v_reg;
  assign mem[322] = mem_322_sv2v_reg;
  assign mem[321] = mem_321_sv2v_reg;
  assign mem[320] = mem_320_sv2v_reg;
  assign mem[319] = mem_319_sv2v_reg;
  assign mem[318] = mem_318_sv2v_reg;
  assign mem[317] = mem_317_sv2v_reg;
  assign mem[316] = mem_316_sv2v_reg;
  assign mem[315] = mem_315_sv2v_reg;
  assign mem[314] = mem_314_sv2v_reg;
  assign mem[313] = mem_313_sv2v_reg;
  assign mem[312] = mem_312_sv2v_reg;
  assign mem[311] = mem_311_sv2v_reg;
  assign mem[310] = mem_310_sv2v_reg;
  assign mem[309] = mem_309_sv2v_reg;
  assign mem[308] = mem_308_sv2v_reg;
  assign mem[307] = mem_307_sv2v_reg;
  assign mem[306] = mem_306_sv2v_reg;
  assign mem[305] = mem_305_sv2v_reg;
  assign mem[304] = mem_304_sv2v_reg;
  assign mem[303] = mem_303_sv2v_reg;
  assign mem[302] = mem_302_sv2v_reg;
  assign mem[301] = mem_301_sv2v_reg;
  assign mem[300] = mem_300_sv2v_reg;
  assign mem[299] = mem_299_sv2v_reg;
  assign mem[298] = mem_298_sv2v_reg;
  assign mem[297] = mem_297_sv2v_reg;
  assign mem[296] = mem_296_sv2v_reg;
  assign mem[295] = mem_295_sv2v_reg;
  assign mem[294] = mem_294_sv2v_reg;
  assign mem[293] = mem_293_sv2v_reg;
  assign mem[292] = mem_292_sv2v_reg;
  assign mem[291] = mem_291_sv2v_reg;
  assign mem[290] = mem_290_sv2v_reg;
  assign mem[289] = mem_289_sv2v_reg;
  assign mem[288] = mem_288_sv2v_reg;
  assign mem[287] = mem_287_sv2v_reg;
  assign mem[286] = mem_286_sv2v_reg;
  assign mem[285] = mem_285_sv2v_reg;
  assign mem[284] = mem_284_sv2v_reg;
  assign mem[283] = mem_283_sv2v_reg;
  assign mem[282] = mem_282_sv2v_reg;
  assign mem[281] = mem_281_sv2v_reg;
  assign mem[280] = mem_280_sv2v_reg;
  assign mem[279] = mem_279_sv2v_reg;
  assign mem[278] = mem_278_sv2v_reg;
  assign mem[277] = mem_277_sv2v_reg;
  assign mem[276] = mem_276_sv2v_reg;
  assign mem[275] = mem_275_sv2v_reg;
  assign mem[274] = mem_274_sv2v_reg;
  assign mem[273] = mem_273_sv2v_reg;
  assign mem[272] = mem_272_sv2v_reg;
  assign mem[271] = mem_271_sv2v_reg;
  assign mem[270] = mem_270_sv2v_reg;
  assign mem[269] = mem_269_sv2v_reg;
  assign mem[268] = mem_268_sv2v_reg;
  assign mem[267] = mem_267_sv2v_reg;
  assign mem[266] = mem_266_sv2v_reg;
  assign mem[265] = mem_265_sv2v_reg;
  assign mem[264] = mem_264_sv2v_reg;
  assign mem[263] = mem_263_sv2v_reg;
  assign mem[262] = mem_262_sv2v_reg;
  assign mem[261] = mem_261_sv2v_reg;
  assign mem[260] = mem_260_sv2v_reg;
  assign mem[259] = mem_259_sv2v_reg;
  assign mem[258] = mem_258_sv2v_reg;
  assign mem[257] = mem_257_sv2v_reg;
  assign mem[256] = mem_256_sv2v_reg;
  assign mem[255] = mem_255_sv2v_reg;
  assign mem[254] = mem_254_sv2v_reg;
  assign mem[253] = mem_253_sv2v_reg;
  assign mem[252] = mem_252_sv2v_reg;
  assign mem[251] = mem_251_sv2v_reg;
  assign mem[250] = mem_250_sv2v_reg;
  assign mem[249] = mem_249_sv2v_reg;
  assign mem[248] = mem_248_sv2v_reg;
  assign mem[247] = mem_247_sv2v_reg;
  assign mem[246] = mem_246_sv2v_reg;
  assign mem[245] = mem_245_sv2v_reg;
  assign mem[244] = mem_244_sv2v_reg;
  assign mem[243] = mem_243_sv2v_reg;
  assign mem[242] = mem_242_sv2v_reg;
  assign mem[241] = mem_241_sv2v_reg;
  assign mem[240] = mem_240_sv2v_reg;
  assign mem[239] = mem_239_sv2v_reg;
  assign mem[238] = mem_238_sv2v_reg;
  assign mem[237] = mem_237_sv2v_reg;
  assign mem[236] = mem_236_sv2v_reg;
  assign mem[235] = mem_235_sv2v_reg;
  assign mem[234] = mem_234_sv2v_reg;
  assign mem[233] = mem_233_sv2v_reg;
  assign mem[232] = mem_232_sv2v_reg;
  assign mem[231] = mem_231_sv2v_reg;
  assign mem[230] = mem_230_sv2v_reg;
  assign mem[229] = mem_229_sv2v_reg;
  assign mem[228] = mem_228_sv2v_reg;
  assign mem[227] = mem_227_sv2v_reg;
  assign mem[226] = mem_226_sv2v_reg;
  assign mem[225] = mem_225_sv2v_reg;
  assign mem[224] = mem_224_sv2v_reg;
  assign mem[223] = mem_223_sv2v_reg;
  assign mem[222] = mem_222_sv2v_reg;
  assign mem[221] = mem_221_sv2v_reg;
  assign mem[220] = mem_220_sv2v_reg;
  assign mem[219] = mem_219_sv2v_reg;
  assign mem[218] = mem_218_sv2v_reg;
  assign mem[217] = mem_217_sv2v_reg;
  assign mem[216] = mem_216_sv2v_reg;
  assign mem[215] = mem_215_sv2v_reg;
  assign mem[214] = mem_214_sv2v_reg;
  assign mem[213] = mem_213_sv2v_reg;
  assign mem[212] = mem_212_sv2v_reg;
  assign mem[211] = mem_211_sv2v_reg;
  assign mem[210] = mem_210_sv2v_reg;
  assign mem[209] = mem_209_sv2v_reg;
  assign mem[208] = mem_208_sv2v_reg;
  assign mem[207] = mem_207_sv2v_reg;
  assign mem[206] = mem_206_sv2v_reg;
  assign mem[205] = mem_205_sv2v_reg;
  assign mem[204] = mem_204_sv2v_reg;
  assign mem[203] = mem_203_sv2v_reg;
  assign mem[202] = mem_202_sv2v_reg;
  assign mem[201] = mem_201_sv2v_reg;
  assign mem[200] = mem_200_sv2v_reg;
  assign mem[199] = mem_199_sv2v_reg;
  assign mem[198] = mem_198_sv2v_reg;
  assign mem[197] = mem_197_sv2v_reg;
  assign mem[196] = mem_196_sv2v_reg;
  assign mem[195] = mem_195_sv2v_reg;
  assign mem[194] = mem_194_sv2v_reg;
  assign mem[193] = mem_193_sv2v_reg;
  assign mem[192] = mem_192_sv2v_reg;
  assign mem[191] = mem_191_sv2v_reg;
  assign mem[190] = mem_190_sv2v_reg;
  assign mem[189] = mem_189_sv2v_reg;
  assign mem[188] = mem_188_sv2v_reg;
  assign mem[187] = mem_187_sv2v_reg;
  assign mem[186] = mem_186_sv2v_reg;
  assign mem[185] = mem_185_sv2v_reg;
  assign mem[184] = mem_184_sv2v_reg;
  assign mem[183] = mem_183_sv2v_reg;
  assign mem[182] = mem_182_sv2v_reg;
  assign mem[181] = mem_181_sv2v_reg;
  assign mem[180] = mem_180_sv2v_reg;
  assign mem[179] = mem_179_sv2v_reg;
  assign mem[178] = mem_178_sv2v_reg;
  assign mem[177] = mem_177_sv2v_reg;
  assign mem[176] = mem_176_sv2v_reg;
  assign mem[175] = mem_175_sv2v_reg;
  assign mem[174] = mem_174_sv2v_reg;
  assign mem[173] = mem_173_sv2v_reg;
  assign mem[172] = mem_172_sv2v_reg;
  assign mem[171] = mem_171_sv2v_reg;
  assign mem[170] = mem_170_sv2v_reg;
  assign mem[169] = mem_169_sv2v_reg;
  assign mem[168] = mem_168_sv2v_reg;
  assign mem[167] = mem_167_sv2v_reg;
  assign mem[166] = mem_166_sv2v_reg;
  assign mem[165] = mem_165_sv2v_reg;
  assign mem[164] = mem_164_sv2v_reg;
  assign mem[163] = mem_163_sv2v_reg;
  assign mem[162] = mem_162_sv2v_reg;
  assign mem[161] = mem_161_sv2v_reg;
  assign mem[160] = mem_160_sv2v_reg;
  assign mem[159] = mem_159_sv2v_reg;
  assign mem[158] = mem_158_sv2v_reg;
  assign mem[157] = mem_157_sv2v_reg;
  assign mem[156] = mem_156_sv2v_reg;
  assign mem[155] = mem_155_sv2v_reg;
  assign mem[154] = mem_154_sv2v_reg;
  assign mem[153] = mem_153_sv2v_reg;
  assign mem[152] = mem_152_sv2v_reg;
  assign mem[151] = mem_151_sv2v_reg;
  assign mem[150] = mem_150_sv2v_reg;
  assign mem[149] = mem_149_sv2v_reg;
  assign mem[148] = mem_148_sv2v_reg;
  assign mem[147] = mem_147_sv2v_reg;
  assign mem[146] = mem_146_sv2v_reg;
  assign mem[145] = mem_145_sv2v_reg;
  assign mem[144] = mem_144_sv2v_reg;
  assign mem[143] = mem_143_sv2v_reg;
  assign mem[142] = mem_142_sv2v_reg;
  assign mem[141] = mem_141_sv2v_reg;
  assign mem[140] = mem_140_sv2v_reg;
  assign mem[139] = mem_139_sv2v_reg;
  assign mem[138] = mem_138_sv2v_reg;
  assign mem[137] = mem_137_sv2v_reg;
  assign mem[136] = mem_136_sv2v_reg;
  assign mem[135] = mem_135_sv2v_reg;
  assign mem[134] = mem_134_sv2v_reg;
  assign mem[133] = mem_133_sv2v_reg;
  assign mem[132] = mem_132_sv2v_reg;
  assign mem[131] = mem_131_sv2v_reg;
  assign mem[130] = mem_130_sv2v_reg;
  assign mem[129] = mem_129_sv2v_reg;
  assign mem[128] = mem_128_sv2v_reg;
  assign mem[127] = mem_127_sv2v_reg;
  assign mem[126] = mem_126_sv2v_reg;
  assign mem[125] = mem_125_sv2v_reg;
  assign mem[124] = mem_124_sv2v_reg;
  assign mem[123] = mem_123_sv2v_reg;
  assign mem[122] = mem_122_sv2v_reg;
  assign mem[121] = mem_121_sv2v_reg;
  assign mem[120] = mem_120_sv2v_reg;
  assign mem[119] = mem_119_sv2v_reg;
  assign mem[118] = mem_118_sv2v_reg;
  assign mem[117] = mem_117_sv2v_reg;
  assign mem[116] = mem_116_sv2v_reg;
  assign mem[115] = mem_115_sv2v_reg;
  assign mem[114] = mem_114_sv2v_reg;
  assign mem[113] = mem_113_sv2v_reg;
  assign mem[112] = mem_112_sv2v_reg;
  assign mem[111] = mem_111_sv2v_reg;
  assign mem[110] = mem_110_sv2v_reg;
  assign mem[109] = mem_109_sv2v_reg;
  assign mem[108] = mem_108_sv2v_reg;
  assign mem[107] = mem_107_sv2v_reg;
  assign mem[106] = mem_106_sv2v_reg;
  assign mem[105] = mem_105_sv2v_reg;
  assign mem[104] = mem_104_sv2v_reg;
  assign mem[103] = mem_103_sv2v_reg;
  assign mem[102] = mem_102_sv2v_reg;
  assign mem[101] = mem_101_sv2v_reg;
  assign mem[100] = mem_100_sv2v_reg;
  assign mem[99] = mem_99_sv2v_reg;
  assign mem[98] = mem_98_sv2v_reg;
  assign mem[97] = mem_97_sv2v_reg;
  assign mem[96] = mem_96_sv2v_reg;
  assign mem[95] = mem_95_sv2v_reg;
  assign mem[94] = mem_94_sv2v_reg;
  assign mem[93] = mem_93_sv2v_reg;
  assign mem[92] = mem_92_sv2v_reg;
  assign mem[91] = mem_91_sv2v_reg;
  assign mem[90] = mem_90_sv2v_reg;
  assign mem[89] = mem_89_sv2v_reg;
  assign mem[88] = mem_88_sv2v_reg;
  assign mem[87] = mem_87_sv2v_reg;
  assign mem[86] = mem_86_sv2v_reg;
  assign mem[85] = mem_85_sv2v_reg;
  assign mem[84] = mem_84_sv2v_reg;
  assign mem[83] = mem_83_sv2v_reg;
  assign mem[82] = mem_82_sv2v_reg;
  assign mem[81] = mem_81_sv2v_reg;
  assign mem[80] = mem_80_sv2v_reg;
  assign mem[79] = mem_79_sv2v_reg;
  assign mem[78] = mem_78_sv2v_reg;
  assign mem[77] = mem_77_sv2v_reg;
  assign mem[76] = mem_76_sv2v_reg;
  assign mem[75] = mem_75_sv2v_reg;
  assign mem[74] = mem_74_sv2v_reg;
  assign mem[73] = mem_73_sv2v_reg;
  assign mem[72] = mem_72_sv2v_reg;
  assign mem[71] = mem_71_sv2v_reg;
  assign mem[70] = mem_70_sv2v_reg;
  assign mem[69] = mem_69_sv2v_reg;
  assign mem[68] = mem_68_sv2v_reg;
  assign mem[67] = mem_67_sv2v_reg;
  assign mem[66] = mem_66_sv2v_reg;
  assign mem[65] = mem_65_sv2v_reg;
  assign mem[64] = mem_64_sv2v_reg;
  assign mem[63] = mem_63_sv2v_reg;
  assign mem[62] = mem_62_sv2v_reg;
  assign mem[61] = mem_61_sv2v_reg;
  assign mem[60] = mem_60_sv2v_reg;
  assign mem[59] = mem_59_sv2v_reg;
  assign mem[58] = mem_58_sv2v_reg;
  assign mem[57] = mem_57_sv2v_reg;
  assign mem[56] = mem_56_sv2v_reg;
  assign mem[55] = mem_55_sv2v_reg;
  assign mem[54] = mem_54_sv2v_reg;
  assign mem[53] = mem_53_sv2v_reg;
  assign mem[52] = mem_52_sv2v_reg;
  assign mem[51] = mem_51_sv2v_reg;
  assign mem[50] = mem_50_sv2v_reg;
  assign mem[49] = mem_49_sv2v_reg;
  assign mem[48] = mem_48_sv2v_reg;
  assign mem[47] = mem_47_sv2v_reg;
  assign mem[46] = mem_46_sv2v_reg;
  assign mem[45] = mem_45_sv2v_reg;
  assign mem[44] = mem_44_sv2v_reg;
  assign mem[43] = mem_43_sv2v_reg;
  assign mem[42] = mem_42_sv2v_reg;
  assign mem[41] = mem_41_sv2v_reg;
  assign mem[40] = mem_40_sv2v_reg;
  assign mem[39] = mem_39_sv2v_reg;
  assign mem[38] = mem_38_sv2v_reg;
  assign mem[37] = mem_37_sv2v_reg;
  assign mem[36] = mem_36_sv2v_reg;
  assign mem[35] = mem_35_sv2v_reg;
  assign mem[34] = mem_34_sv2v_reg;
  assign mem[33] = mem_33_sv2v_reg;
  assign mem[32] = mem_32_sv2v_reg;
  assign mem[31] = mem_31_sv2v_reg;
  assign mem[30] = mem_30_sv2v_reg;
  assign mem[29] = mem_29_sv2v_reg;
  assign mem[28] = mem_28_sv2v_reg;
  assign mem[27] = mem_27_sv2v_reg;
  assign mem[26] = mem_26_sv2v_reg;
  assign mem[25] = mem_25_sv2v_reg;
  assign mem[24] = mem_24_sv2v_reg;
  assign mem[23] = mem_23_sv2v_reg;
  assign mem[22] = mem_22_sv2v_reg;
  assign mem[21] = mem_21_sv2v_reg;
  assign mem[20] = mem_20_sv2v_reg;
  assign mem[19] = mem_19_sv2v_reg;
  assign mem[18] = mem_18_sv2v_reg;
  assign mem[17] = mem_17_sv2v_reg;
  assign mem[16] = mem_16_sv2v_reg;
  assign mem[15] = mem_15_sv2v_reg;
  assign mem[14] = mem_14_sv2v_reg;
  assign mem[13] = mem_13_sv2v_reg;
  assign mem[12] = mem_12_sv2v_reg;
  assign mem[11] = mem_11_sv2v_reg;
  assign mem[10] = mem_10_sv2v_reg;
  assign mem[9] = mem_9_sv2v_reg;
  assign mem[8] = mem_8_sv2v_reg;
  assign mem[7] = mem_7_sv2v_reg;
  assign mem[6] = mem_6_sv2v_reg;
  assign mem[5] = mem_5_sv2v_reg;
  assign mem[4] = mem_4_sv2v_reg;
  assign mem[3] = mem_3_sv2v_reg;
  assign mem[2] = mem_2_sv2v_reg;
  assign mem[1] = mem_1_sv2v_reg;
  assign mem[0] = mem_0_sv2v_reg;
  assign r_data_o[15] = (N76)? mem[15] : 
                        (N78)? mem[31] : 
                        (N80)? mem[47] : 
                        (N82)? mem[63] : 
                        (N84)? mem[79] : 
                        (N86)? mem[95] : 
                        (N88)? mem[111] : 
                        (N90)? mem[127] : 
                        (N92)? mem[143] : 
                        (N94)? mem[159] : 
                        (N96)? mem[175] : 
                        (N98)? mem[191] : 
                        (N100)? mem[207] : 
                        (N102)? mem[223] : 
                        (N104)? mem[239] : 
                        (N106)? mem[255] : 
                        (N108)? mem[271] : 
                        (N110)? mem[287] : 
                        (N112)? mem[303] : 
                        (N114)? mem[319] : 
                        (N116)? mem[335] : 
                        (N118)? mem[351] : 
                        (N120)? mem[367] : 
                        (N122)? mem[383] : 
                        (N124)? mem[399] : 
                        (N126)? mem[415] : 
                        (N128)? mem[431] : 
                        (N130)? mem[447] : 
                        (N132)? mem[463] : 
                        (N134)? mem[479] : 
                        (N136)? mem[495] : 
                        (N138)? mem[511] : 
                        (N77)? mem[527] : 
                        (N79)? mem[543] : 
                        (N81)? mem[559] : 
                        (N83)? mem[575] : 
                        (N85)? mem[591] : 
                        (N87)? mem[607] : 
                        (N89)? mem[623] : 
                        (N91)? mem[639] : 
                        (N93)? mem[655] : 
                        (N95)? mem[671] : 
                        (N97)? mem[687] : 
                        (N99)? mem[703] : 
                        (N101)? mem[719] : 
                        (N103)? mem[735] : 
                        (N105)? mem[751] : 
                        (N107)? mem[767] : 
                        (N109)? mem[783] : 
                        (N111)? mem[799] : 
                        (N113)? mem[815] : 
                        (N115)? mem[831] : 
                        (N117)? mem[847] : 
                        (N119)? mem[863] : 
                        (N121)? mem[879] : 
                        (N123)? mem[895] : 
                        (N125)? mem[911] : 
                        (N127)? mem[927] : 
                        (N129)? mem[943] : 
                        (N131)? mem[959] : 
                        (N133)? mem[975] : 
                        (N135)? mem[991] : 
                        (N137)? mem[1007] : 
                        (N139)? mem[1023] : 1'b0;
  assign r_data_o[14] = (N76)? mem[14] : 
                        (N78)? mem[30] : 
                        (N80)? mem[46] : 
                        (N82)? mem[62] : 
                        (N84)? mem[78] : 
                        (N86)? mem[94] : 
                        (N88)? mem[110] : 
                        (N90)? mem[126] : 
                        (N92)? mem[142] : 
                        (N94)? mem[158] : 
                        (N96)? mem[174] : 
                        (N98)? mem[190] : 
                        (N100)? mem[206] : 
                        (N102)? mem[222] : 
                        (N104)? mem[238] : 
                        (N106)? mem[254] : 
                        (N108)? mem[270] : 
                        (N110)? mem[286] : 
                        (N112)? mem[302] : 
                        (N114)? mem[318] : 
                        (N116)? mem[334] : 
                        (N118)? mem[350] : 
                        (N120)? mem[366] : 
                        (N122)? mem[382] : 
                        (N124)? mem[398] : 
                        (N126)? mem[414] : 
                        (N128)? mem[430] : 
                        (N130)? mem[446] : 
                        (N132)? mem[462] : 
                        (N134)? mem[478] : 
                        (N136)? mem[494] : 
                        (N138)? mem[510] : 
                        (N77)? mem[526] : 
                        (N79)? mem[542] : 
                        (N81)? mem[558] : 
                        (N83)? mem[574] : 
                        (N85)? mem[590] : 
                        (N87)? mem[606] : 
                        (N89)? mem[622] : 
                        (N91)? mem[638] : 
                        (N93)? mem[654] : 
                        (N95)? mem[670] : 
                        (N97)? mem[686] : 
                        (N99)? mem[702] : 
                        (N101)? mem[718] : 
                        (N103)? mem[734] : 
                        (N105)? mem[750] : 
                        (N107)? mem[766] : 
                        (N109)? mem[782] : 
                        (N111)? mem[798] : 
                        (N113)? mem[814] : 
                        (N115)? mem[830] : 
                        (N117)? mem[846] : 
                        (N119)? mem[862] : 
                        (N121)? mem[878] : 
                        (N123)? mem[894] : 
                        (N125)? mem[910] : 
                        (N127)? mem[926] : 
                        (N129)? mem[942] : 
                        (N131)? mem[958] : 
                        (N133)? mem[974] : 
                        (N135)? mem[990] : 
                        (N137)? mem[1006] : 
                        (N139)? mem[1022] : 1'b0;
  assign r_data_o[13] = (N76)? mem[13] : 
                        (N78)? mem[29] : 
                        (N80)? mem[45] : 
                        (N82)? mem[61] : 
                        (N84)? mem[77] : 
                        (N86)? mem[93] : 
                        (N88)? mem[109] : 
                        (N90)? mem[125] : 
                        (N92)? mem[141] : 
                        (N94)? mem[157] : 
                        (N96)? mem[173] : 
                        (N98)? mem[189] : 
                        (N100)? mem[205] : 
                        (N102)? mem[221] : 
                        (N104)? mem[237] : 
                        (N106)? mem[253] : 
                        (N108)? mem[269] : 
                        (N110)? mem[285] : 
                        (N112)? mem[301] : 
                        (N114)? mem[317] : 
                        (N116)? mem[333] : 
                        (N118)? mem[349] : 
                        (N120)? mem[365] : 
                        (N122)? mem[381] : 
                        (N124)? mem[397] : 
                        (N126)? mem[413] : 
                        (N128)? mem[429] : 
                        (N130)? mem[445] : 
                        (N132)? mem[461] : 
                        (N134)? mem[477] : 
                        (N136)? mem[493] : 
                        (N138)? mem[509] : 
                        (N77)? mem[525] : 
                        (N79)? mem[541] : 
                        (N81)? mem[557] : 
                        (N83)? mem[573] : 
                        (N85)? mem[589] : 
                        (N87)? mem[605] : 
                        (N89)? mem[621] : 
                        (N91)? mem[637] : 
                        (N93)? mem[653] : 
                        (N95)? mem[669] : 
                        (N97)? mem[685] : 
                        (N99)? mem[701] : 
                        (N101)? mem[717] : 
                        (N103)? mem[733] : 
                        (N105)? mem[749] : 
                        (N107)? mem[765] : 
                        (N109)? mem[781] : 
                        (N111)? mem[797] : 
                        (N113)? mem[813] : 
                        (N115)? mem[829] : 
                        (N117)? mem[845] : 
                        (N119)? mem[861] : 
                        (N121)? mem[877] : 
                        (N123)? mem[893] : 
                        (N125)? mem[909] : 
                        (N127)? mem[925] : 
                        (N129)? mem[941] : 
                        (N131)? mem[957] : 
                        (N133)? mem[973] : 
                        (N135)? mem[989] : 
                        (N137)? mem[1005] : 
                        (N139)? mem[1021] : 1'b0;
  assign r_data_o[12] = (N76)? mem[12] : 
                        (N78)? mem[28] : 
                        (N80)? mem[44] : 
                        (N82)? mem[60] : 
                        (N84)? mem[76] : 
                        (N86)? mem[92] : 
                        (N88)? mem[108] : 
                        (N90)? mem[124] : 
                        (N92)? mem[140] : 
                        (N94)? mem[156] : 
                        (N96)? mem[172] : 
                        (N98)? mem[188] : 
                        (N100)? mem[204] : 
                        (N102)? mem[220] : 
                        (N104)? mem[236] : 
                        (N106)? mem[252] : 
                        (N108)? mem[268] : 
                        (N110)? mem[284] : 
                        (N112)? mem[300] : 
                        (N114)? mem[316] : 
                        (N116)? mem[332] : 
                        (N118)? mem[348] : 
                        (N120)? mem[364] : 
                        (N122)? mem[380] : 
                        (N124)? mem[396] : 
                        (N126)? mem[412] : 
                        (N128)? mem[428] : 
                        (N130)? mem[444] : 
                        (N132)? mem[460] : 
                        (N134)? mem[476] : 
                        (N136)? mem[492] : 
                        (N138)? mem[508] : 
                        (N77)? mem[524] : 
                        (N79)? mem[540] : 
                        (N81)? mem[556] : 
                        (N83)? mem[572] : 
                        (N85)? mem[588] : 
                        (N87)? mem[604] : 
                        (N89)? mem[620] : 
                        (N91)? mem[636] : 
                        (N93)? mem[652] : 
                        (N95)? mem[668] : 
                        (N97)? mem[684] : 
                        (N99)? mem[700] : 
                        (N101)? mem[716] : 
                        (N103)? mem[732] : 
                        (N105)? mem[748] : 
                        (N107)? mem[764] : 
                        (N109)? mem[780] : 
                        (N111)? mem[796] : 
                        (N113)? mem[812] : 
                        (N115)? mem[828] : 
                        (N117)? mem[844] : 
                        (N119)? mem[860] : 
                        (N121)? mem[876] : 
                        (N123)? mem[892] : 
                        (N125)? mem[908] : 
                        (N127)? mem[924] : 
                        (N129)? mem[940] : 
                        (N131)? mem[956] : 
                        (N133)? mem[972] : 
                        (N135)? mem[988] : 
                        (N137)? mem[1004] : 
                        (N139)? mem[1020] : 1'b0;
  assign r_data_o[11] = (N76)? mem[11] : 
                        (N78)? mem[27] : 
                        (N80)? mem[43] : 
                        (N82)? mem[59] : 
                        (N84)? mem[75] : 
                        (N86)? mem[91] : 
                        (N88)? mem[107] : 
                        (N90)? mem[123] : 
                        (N92)? mem[139] : 
                        (N94)? mem[155] : 
                        (N96)? mem[171] : 
                        (N98)? mem[187] : 
                        (N100)? mem[203] : 
                        (N102)? mem[219] : 
                        (N104)? mem[235] : 
                        (N106)? mem[251] : 
                        (N108)? mem[267] : 
                        (N110)? mem[283] : 
                        (N112)? mem[299] : 
                        (N114)? mem[315] : 
                        (N116)? mem[331] : 
                        (N118)? mem[347] : 
                        (N120)? mem[363] : 
                        (N122)? mem[379] : 
                        (N124)? mem[395] : 
                        (N126)? mem[411] : 
                        (N128)? mem[427] : 
                        (N130)? mem[443] : 
                        (N132)? mem[459] : 
                        (N134)? mem[475] : 
                        (N136)? mem[491] : 
                        (N138)? mem[507] : 
                        (N77)? mem[523] : 
                        (N79)? mem[539] : 
                        (N81)? mem[555] : 
                        (N83)? mem[571] : 
                        (N85)? mem[587] : 
                        (N87)? mem[603] : 
                        (N89)? mem[619] : 
                        (N91)? mem[635] : 
                        (N93)? mem[651] : 
                        (N95)? mem[667] : 
                        (N97)? mem[683] : 
                        (N99)? mem[699] : 
                        (N101)? mem[715] : 
                        (N103)? mem[731] : 
                        (N105)? mem[747] : 
                        (N107)? mem[763] : 
                        (N109)? mem[779] : 
                        (N111)? mem[795] : 
                        (N113)? mem[811] : 
                        (N115)? mem[827] : 
                        (N117)? mem[843] : 
                        (N119)? mem[859] : 
                        (N121)? mem[875] : 
                        (N123)? mem[891] : 
                        (N125)? mem[907] : 
                        (N127)? mem[923] : 
                        (N129)? mem[939] : 
                        (N131)? mem[955] : 
                        (N133)? mem[971] : 
                        (N135)? mem[987] : 
                        (N137)? mem[1003] : 
                        (N139)? mem[1019] : 1'b0;
  assign r_data_o[10] = (N76)? mem[10] : 
                        (N78)? mem[26] : 
                        (N80)? mem[42] : 
                        (N82)? mem[58] : 
                        (N84)? mem[74] : 
                        (N86)? mem[90] : 
                        (N88)? mem[106] : 
                        (N90)? mem[122] : 
                        (N92)? mem[138] : 
                        (N94)? mem[154] : 
                        (N96)? mem[170] : 
                        (N98)? mem[186] : 
                        (N100)? mem[202] : 
                        (N102)? mem[218] : 
                        (N104)? mem[234] : 
                        (N106)? mem[250] : 
                        (N108)? mem[266] : 
                        (N110)? mem[282] : 
                        (N112)? mem[298] : 
                        (N114)? mem[314] : 
                        (N116)? mem[330] : 
                        (N118)? mem[346] : 
                        (N120)? mem[362] : 
                        (N122)? mem[378] : 
                        (N124)? mem[394] : 
                        (N126)? mem[410] : 
                        (N128)? mem[426] : 
                        (N130)? mem[442] : 
                        (N132)? mem[458] : 
                        (N134)? mem[474] : 
                        (N136)? mem[490] : 
                        (N138)? mem[506] : 
                        (N77)? mem[522] : 
                        (N79)? mem[538] : 
                        (N81)? mem[554] : 
                        (N83)? mem[570] : 
                        (N85)? mem[586] : 
                        (N87)? mem[602] : 
                        (N89)? mem[618] : 
                        (N91)? mem[634] : 
                        (N93)? mem[650] : 
                        (N95)? mem[666] : 
                        (N97)? mem[682] : 
                        (N99)? mem[698] : 
                        (N101)? mem[714] : 
                        (N103)? mem[730] : 
                        (N105)? mem[746] : 
                        (N107)? mem[762] : 
                        (N109)? mem[778] : 
                        (N111)? mem[794] : 
                        (N113)? mem[810] : 
                        (N115)? mem[826] : 
                        (N117)? mem[842] : 
                        (N119)? mem[858] : 
                        (N121)? mem[874] : 
                        (N123)? mem[890] : 
                        (N125)? mem[906] : 
                        (N127)? mem[922] : 
                        (N129)? mem[938] : 
                        (N131)? mem[954] : 
                        (N133)? mem[970] : 
                        (N135)? mem[986] : 
                        (N137)? mem[1002] : 
                        (N139)? mem[1018] : 1'b0;
  assign r_data_o[9] = (N76)? mem[9] : 
                       (N78)? mem[25] : 
                       (N80)? mem[41] : 
                       (N82)? mem[57] : 
                       (N84)? mem[73] : 
                       (N86)? mem[89] : 
                       (N88)? mem[105] : 
                       (N90)? mem[121] : 
                       (N92)? mem[137] : 
                       (N94)? mem[153] : 
                       (N96)? mem[169] : 
                       (N98)? mem[185] : 
                       (N100)? mem[201] : 
                       (N102)? mem[217] : 
                       (N104)? mem[233] : 
                       (N106)? mem[249] : 
                       (N108)? mem[265] : 
                       (N110)? mem[281] : 
                       (N112)? mem[297] : 
                       (N114)? mem[313] : 
                       (N116)? mem[329] : 
                       (N118)? mem[345] : 
                       (N120)? mem[361] : 
                       (N122)? mem[377] : 
                       (N124)? mem[393] : 
                       (N126)? mem[409] : 
                       (N128)? mem[425] : 
                       (N130)? mem[441] : 
                       (N132)? mem[457] : 
                       (N134)? mem[473] : 
                       (N136)? mem[489] : 
                       (N138)? mem[505] : 
                       (N77)? mem[521] : 
                       (N79)? mem[537] : 
                       (N81)? mem[553] : 
                       (N83)? mem[569] : 
                       (N85)? mem[585] : 
                       (N87)? mem[601] : 
                       (N89)? mem[617] : 
                       (N91)? mem[633] : 
                       (N93)? mem[649] : 
                       (N95)? mem[665] : 
                       (N97)? mem[681] : 
                       (N99)? mem[697] : 
                       (N101)? mem[713] : 
                       (N103)? mem[729] : 
                       (N105)? mem[745] : 
                       (N107)? mem[761] : 
                       (N109)? mem[777] : 
                       (N111)? mem[793] : 
                       (N113)? mem[809] : 
                       (N115)? mem[825] : 
                       (N117)? mem[841] : 
                       (N119)? mem[857] : 
                       (N121)? mem[873] : 
                       (N123)? mem[889] : 
                       (N125)? mem[905] : 
                       (N127)? mem[921] : 
                       (N129)? mem[937] : 
                       (N131)? mem[953] : 
                       (N133)? mem[969] : 
                       (N135)? mem[985] : 
                       (N137)? mem[1001] : 
                       (N139)? mem[1017] : 1'b0;
  assign r_data_o[8] = (N76)? mem[8] : 
                       (N78)? mem[24] : 
                       (N80)? mem[40] : 
                       (N82)? mem[56] : 
                       (N84)? mem[72] : 
                       (N86)? mem[88] : 
                       (N88)? mem[104] : 
                       (N90)? mem[120] : 
                       (N92)? mem[136] : 
                       (N94)? mem[152] : 
                       (N96)? mem[168] : 
                       (N98)? mem[184] : 
                       (N100)? mem[200] : 
                       (N102)? mem[216] : 
                       (N104)? mem[232] : 
                       (N106)? mem[248] : 
                       (N108)? mem[264] : 
                       (N110)? mem[280] : 
                       (N112)? mem[296] : 
                       (N114)? mem[312] : 
                       (N116)? mem[328] : 
                       (N118)? mem[344] : 
                       (N120)? mem[360] : 
                       (N122)? mem[376] : 
                       (N124)? mem[392] : 
                       (N126)? mem[408] : 
                       (N128)? mem[424] : 
                       (N130)? mem[440] : 
                       (N132)? mem[456] : 
                       (N134)? mem[472] : 
                       (N136)? mem[488] : 
                       (N138)? mem[504] : 
                       (N77)? mem[520] : 
                       (N79)? mem[536] : 
                       (N81)? mem[552] : 
                       (N83)? mem[568] : 
                       (N85)? mem[584] : 
                       (N87)? mem[600] : 
                       (N89)? mem[616] : 
                       (N91)? mem[632] : 
                       (N93)? mem[648] : 
                       (N95)? mem[664] : 
                       (N97)? mem[680] : 
                       (N99)? mem[696] : 
                       (N101)? mem[712] : 
                       (N103)? mem[728] : 
                       (N105)? mem[744] : 
                       (N107)? mem[760] : 
                       (N109)? mem[776] : 
                       (N111)? mem[792] : 
                       (N113)? mem[808] : 
                       (N115)? mem[824] : 
                       (N117)? mem[840] : 
                       (N119)? mem[856] : 
                       (N121)? mem[872] : 
                       (N123)? mem[888] : 
                       (N125)? mem[904] : 
                       (N127)? mem[920] : 
                       (N129)? mem[936] : 
                       (N131)? mem[952] : 
                       (N133)? mem[968] : 
                       (N135)? mem[984] : 
                       (N137)? mem[1000] : 
                       (N139)? mem[1016] : 1'b0;
  assign r_data_o[7] = (N76)? mem[7] : 
                       (N78)? mem[23] : 
                       (N80)? mem[39] : 
                       (N82)? mem[55] : 
                       (N84)? mem[71] : 
                       (N86)? mem[87] : 
                       (N88)? mem[103] : 
                       (N90)? mem[119] : 
                       (N92)? mem[135] : 
                       (N94)? mem[151] : 
                       (N96)? mem[167] : 
                       (N98)? mem[183] : 
                       (N100)? mem[199] : 
                       (N102)? mem[215] : 
                       (N104)? mem[231] : 
                       (N106)? mem[247] : 
                       (N108)? mem[263] : 
                       (N110)? mem[279] : 
                       (N112)? mem[295] : 
                       (N114)? mem[311] : 
                       (N116)? mem[327] : 
                       (N118)? mem[343] : 
                       (N120)? mem[359] : 
                       (N122)? mem[375] : 
                       (N124)? mem[391] : 
                       (N126)? mem[407] : 
                       (N128)? mem[423] : 
                       (N130)? mem[439] : 
                       (N132)? mem[455] : 
                       (N134)? mem[471] : 
                       (N136)? mem[487] : 
                       (N138)? mem[503] : 
                       (N77)? mem[519] : 
                       (N79)? mem[535] : 
                       (N81)? mem[551] : 
                       (N83)? mem[567] : 
                       (N85)? mem[583] : 
                       (N87)? mem[599] : 
                       (N89)? mem[615] : 
                       (N91)? mem[631] : 
                       (N93)? mem[647] : 
                       (N95)? mem[663] : 
                       (N97)? mem[679] : 
                       (N99)? mem[695] : 
                       (N101)? mem[711] : 
                       (N103)? mem[727] : 
                       (N105)? mem[743] : 
                       (N107)? mem[759] : 
                       (N109)? mem[775] : 
                       (N111)? mem[791] : 
                       (N113)? mem[807] : 
                       (N115)? mem[823] : 
                       (N117)? mem[839] : 
                       (N119)? mem[855] : 
                       (N121)? mem[871] : 
                       (N123)? mem[887] : 
                       (N125)? mem[903] : 
                       (N127)? mem[919] : 
                       (N129)? mem[935] : 
                       (N131)? mem[951] : 
                       (N133)? mem[967] : 
                       (N135)? mem[983] : 
                       (N137)? mem[999] : 
                       (N139)? mem[1015] : 1'b0;
  assign r_data_o[6] = (N76)? mem[6] : 
                       (N78)? mem[22] : 
                       (N80)? mem[38] : 
                       (N82)? mem[54] : 
                       (N84)? mem[70] : 
                       (N86)? mem[86] : 
                       (N88)? mem[102] : 
                       (N90)? mem[118] : 
                       (N92)? mem[134] : 
                       (N94)? mem[150] : 
                       (N96)? mem[166] : 
                       (N98)? mem[182] : 
                       (N100)? mem[198] : 
                       (N102)? mem[214] : 
                       (N104)? mem[230] : 
                       (N106)? mem[246] : 
                       (N108)? mem[262] : 
                       (N110)? mem[278] : 
                       (N112)? mem[294] : 
                       (N114)? mem[310] : 
                       (N116)? mem[326] : 
                       (N118)? mem[342] : 
                       (N120)? mem[358] : 
                       (N122)? mem[374] : 
                       (N124)? mem[390] : 
                       (N126)? mem[406] : 
                       (N128)? mem[422] : 
                       (N130)? mem[438] : 
                       (N132)? mem[454] : 
                       (N134)? mem[470] : 
                       (N136)? mem[486] : 
                       (N138)? mem[502] : 
                       (N77)? mem[518] : 
                       (N79)? mem[534] : 
                       (N81)? mem[550] : 
                       (N83)? mem[566] : 
                       (N85)? mem[582] : 
                       (N87)? mem[598] : 
                       (N89)? mem[614] : 
                       (N91)? mem[630] : 
                       (N93)? mem[646] : 
                       (N95)? mem[662] : 
                       (N97)? mem[678] : 
                       (N99)? mem[694] : 
                       (N101)? mem[710] : 
                       (N103)? mem[726] : 
                       (N105)? mem[742] : 
                       (N107)? mem[758] : 
                       (N109)? mem[774] : 
                       (N111)? mem[790] : 
                       (N113)? mem[806] : 
                       (N115)? mem[822] : 
                       (N117)? mem[838] : 
                       (N119)? mem[854] : 
                       (N121)? mem[870] : 
                       (N123)? mem[886] : 
                       (N125)? mem[902] : 
                       (N127)? mem[918] : 
                       (N129)? mem[934] : 
                       (N131)? mem[950] : 
                       (N133)? mem[966] : 
                       (N135)? mem[982] : 
                       (N137)? mem[998] : 
                       (N139)? mem[1014] : 1'b0;
  assign r_data_o[5] = (N76)? mem[5] : 
                       (N78)? mem[21] : 
                       (N80)? mem[37] : 
                       (N82)? mem[53] : 
                       (N84)? mem[69] : 
                       (N86)? mem[85] : 
                       (N88)? mem[101] : 
                       (N90)? mem[117] : 
                       (N92)? mem[133] : 
                       (N94)? mem[149] : 
                       (N96)? mem[165] : 
                       (N98)? mem[181] : 
                       (N100)? mem[197] : 
                       (N102)? mem[213] : 
                       (N104)? mem[229] : 
                       (N106)? mem[245] : 
                       (N108)? mem[261] : 
                       (N110)? mem[277] : 
                       (N112)? mem[293] : 
                       (N114)? mem[309] : 
                       (N116)? mem[325] : 
                       (N118)? mem[341] : 
                       (N120)? mem[357] : 
                       (N122)? mem[373] : 
                       (N124)? mem[389] : 
                       (N126)? mem[405] : 
                       (N128)? mem[421] : 
                       (N130)? mem[437] : 
                       (N132)? mem[453] : 
                       (N134)? mem[469] : 
                       (N136)? mem[485] : 
                       (N138)? mem[501] : 
                       (N77)? mem[517] : 
                       (N79)? mem[533] : 
                       (N81)? mem[549] : 
                       (N83)? mem[565] : 
                       (N85)? mem[581] : 
                       (N87)? mem[597] : 
                       (N89)? mem[613] : 
                       (N91)? mem[629] : 
                       (N93)? mem[645] : 
                       (N95)? mem[661] : 
                       (N97)? mem[677] : 
                       (N99)? mem[693] : 
                       (N101)? mem[709] : 
                       (N103)? mem[725] : 
                       (N105)? mem[741] : 
                       (N107)? mem[757] : 
                       (N109)? mem[773] : 
                       (N111)? mem[789] : 
                       (N113)? mem[805] : 
                       (N115)? mem[821] : 
                       (N117)? mem[837] : 
                       (N119)? mem[853] : 
                       (N121)? mem[869] : 
                       (N123)? mem[885] : 
                       (N125)? mem[901] : 
                       (N127)? mem[917] : 
                       (N129)? mem[933] : 
                       (N131)? mem[949] : 
                       (N133)? mem[965] : 
                       (N135)? mem[981] : 
                       (N137)? mem[997] : 
                       (N139)? mem[1013] : 1'b0;
  assign r_data_o[4] = (N76)? mem[4] : 
                       (N78)? mem[20] : 
                       (N80)? mem[36] : 
                       (N82)? mem[52] : 
                       (N84)? mem[68] : 
                       (N86)? mem[84] : 
                       (N88)? mem[100] : 
                       (N90)? mem[116] : 
                       (N92)? mem[132] : 
                       (N94)? mem[148] : 
                       (N96)? mem[164] : 
                       (N98)? mem[180] : 
                       (N100)? mem[196] : 
                       (N102)? mem[212] : 
                       (N104)? mem[228] : 
                       (N106)? mem[244] : 
                       (N108)? mem[260] : 
                       (N110)? mem[276] : 
                       (N112)? mem[292] : 
                       (N114)? mem[308] : 
                       (N116)? mem[324] : 
                       (N118)? mem[340] : 
                       (N120)? mem[356] : 
                       (N122)? mem[372] : 
                       (N124)? mem[388] : 
                       (N126)? mem[404] : 
                       (N128)? mem[420] : 
                       (N130)? mem[436] : 
                       (N132)? mem[452] : 
                       (N134)? mem[468] : 
                       (N136)? mem[484] : 
                       (N138)? mem[500] : 
                       (N77)? mem[516] : 
                       (N79)? mem[532] : 
                       (N81)? mem[548] : 
                       (N83)? mem[564] : 
                       (N85)? mem[580] : 
                       (N87)? mem[596] : 
                       (N89)? mem[612] : 
                       (N91)? mem[628] : 
                       (N93)? mem[644] : 
                       (N95)? mem[660] : 
                       (N97)? mem[676] : 
                       (N99)? mem[692] : 
                       (N101)? mem[708] : 
                       (N103)? mem[724] : 
                       (N105)? mem[740] : 
                       (N107)? mem[756] : 
                       (N109)? mem[772] : 
                       (N111)? mem[788] : 
                       (N113)? mem[804] : 
                       (N115)? mem[820] : 
                       (N117)? mem[836] : 
                       (N119)? mem[852] : 
                       (N121)? mem[868] : 
                       (N123)? mem[884] : 
                       (N125)? mem[900] : 
                       (N127)? mem[916] : 
                       (N129)? mem[932] : 
                       (N131)? mem[948] : 
                       (N133)? mem[964] : 
                       (N135)? mem[980] : 
                       (N137)? mem[996] : 
                       (N139)? mem[1012] : 1'b0;
  assign r_data_o[3] = (N76)? mem[3] : 
                       (N78)? mem[19] : 
                       (N80)? mem[35] : 
                       (N82)? mem[51] : 
                       (N84)? mem[67] : 
                       (N86)? mem[83] : 
                       (N88)? mem[99] : 
                       (N90)? mem[115] : 
                       (N92)? mem[131] : 
                       (N94)? mem[147] : 
                       (N96)? mem[163] : 
                       (N98)? mem[179] : 
                       (N100)? mem[195] : 
                       (N102)? mem[211] : 
                       (N104)? mem[227] : 
                       (N106)? mem[243] : 
                       (N108)? mem[259] : 
                       (N110)? mem[275] : 
                       (N112)? mem[291] : 
                       (N114)? mem[307] : 
                       (N116)? mem[323] : 
                       (N118)? mem[339] : 
                       (N120)? mem[355] : 
                       (N122)? mem[371] : 
                       (N124)? mem[387] : 
                       (N126)? mem[403] : 
                       (N128)? mem[419] : 
                       (N130)? mem[435] : 
                       (N132)? mem[451] : 
                       (N134)? mem[467] : 
                       (N136)? mem[483] : 
                       (N138)? mem[499] : 
                       (N77)? mem[515] : 
                       (N79)? mem[531] : 
                       (N81)? mem[547] : 
                       (N83)? mem[563] : 
                       (N85)? mem[579] : 
                       (N87)? mem[595] : 
                       (N89)? mem[611] : 
                       (N91)? mem[627] : 
                       (N93)? mem[643] : 
                       (N95)? mem[659] : 
                       (N97)? mem[675] : 
                       (N99)? mem[691] : 
                       (N101)? mem[707] : 
                       (N103)? mem[723] : 
                       (N105)? mem[739] : 
                       (N107)? mem[755] : 
                       (N109)? mem[771] : 
                       (N111)? mem[787] : 
                       (N113)? mem[803] : 
                       (N115)? mem[819] : 
                       (N117)? mem[835] : 
                       (N119)? mem[851] : 
                       (N121)? mem[867] : 
                       (N123)? mem[883] : 
                       (N125)? mem[899] : 
                       (N127)? mem[915] : 
                       (N129)? mem[931] : 
                       (N131)? mem[947] : 
                       (N133)? mem[963] : 
                       (N135)? mem[979] : 
                       (N137)? mem[995] : 
                       (N139)? mem[1011] : 1'b0;
  assign r_data_o[2] = (N76)? mem[2] : 
                       (N78)? mem[18] : 
                       (N80)? mem[34] : 
                       (N82)? mem[50] : 
                       (N84)? mem[66] : 
                       (N86)? mem[82] : 
                       (N88)? mem[98] : 
                       (N90)? mem[114] : 
                       (N92)? mem[130] : 
                       (N94)? mem[146] : 
                       (N96)? mem[162] : 
                       (N98)? mem[178] : 
                       (N100)? mem[194] : 
                       (N102)? mem[210] : 
                       (N104)? mem[226] : 
                       (N106)? mem[242] : 
                       (N108)? mem[258] : 
                       (N110)? mem[274] : 
                       (N112)? mem[290] : 
                       (N114)? mem[306] : 
                       (N116)? mem[322] : 
                       (N118)? mem[338] : 
                       (N120)? mem[354] : 
                       (N122)? mem[370] : 
                       (N124)? mem[386] : 
                       (N126)? mem[402] : 
                       (N128)? mem[418] : 
                       (N130)? mem[434] : 
                       (N132)? mem[450] : 
                       (N134)? mem[466] : 
                       (N136)? mem[482] : 
                       (N138)? mem[498] : 
                       (N77)? mem[514] : 
                       (N79)? mem[530] : 
                       (N81)? mem[546] : 
                       (N83)? mem[562] : 
                       (N85)? mem[578] : 
                       (N87)? mem[594] : 
                       (N89)? mem[610] : 
                       (N91)? mem[626] : 
                       (N93)? mem[642] : 
                       (N95)? mem[658] : 
                       (N97)? mem[674] : 
                       (N99)? mem[690] : 
                       (N101)? mem[706] : 
                       (N103)? mem[722] : 
                       (N105)? mem[738] : 
                       (N107)? mem[754] : 
                       (N109)? mem[770] : 
                       (N111)? mem[786] : 
                       (N113)? mem[802] : 
                       (N115)? mem[818] : 
                       (N117)? mem[834] : 
                       (N119)? mem[850] : 
                       (N121)? mem[866] : 
                       (N123)? mem[882] : 
                       (N125)? mem[898] : 
                       (N127)? mem[914] : 
                       (N129)? mem[930] : 
                       (N131)? mem[946] : 
                       (N133)? mem[962] : 
                       (N135)? mem[978] : 
                       (N137)? mem[994] : 
                       (N139)? mem[1010] : 1'b0;
  assign r_data_o[1] = (N76)? mem[1] : 
                       (N78)? mem[17] : 
                       (N80)? mem[33] : 
                       (N82)? mem[49] : 
                       (N84)? mem[65] : 
                       (N86)? mem[81] : 
                       (N88)? mem[97] : 
                       (N90)? mem[113] : 
                       (N92)? mem[129] : 
                       (N94)? mem[145] : 
                       (N96)? mem[161] : 
                       (N98)? mem[177] : 
                       (N100)? mem[193] : 
                       (N102)? mem[209] : 
                       (N104)? mem[225] : 
                       (N106)? mem[241] : 
                       (N108)? mem[257] : 
                       (N110)? mem[273] : 
                       (N112)? mem[289] : 
                       (N114)? mem[305] : 
                       (N116)? mem[321] : 
                       (N118)? mem[337] : 
                       (N120)? mem[353] : 
                       (N122)? mem[369] : 
                       (N124)? mem[385] : 
                       (N126)? mem[401] : 
                       (N128)? mem[417] : 
                       (N130)? mem[433] : 
                       (N132)? mem[449] : 
                       (N134)? mem[465] : 
                       (N136)? mem[481] : 
                       (N138)? mem[497] : 
                       (N77)? mem[513] : 
                       (N79)? mem[529] : 
                       (N81)? mem[545] : 
                       (N83)? mem[561] : 
                       (N85)? mem[577] : 
                       (N87)? mem[593] : 
                       (N89)? mem[609] : 
                       (N91)? mem[625] : 
                       (N93)? mem[641] : 
                       (N95)? mem[657] : 
                       (N97)? mem[673] : 
                       (N99)? mem[689] : 
                       (N101)? mem[705] : 
                       (N103)? mem[721] : 
                       (N105)? mem[737] : 
                       (N107)? mem[753] : 
                       (N109)? mem[769] : 
                       (N111)? mem[785] : 
                       (N113)? mem[801] : 
                       (N115)? mem[817] : 
                       (N117)? mem[833] : 
                       (N119)? mem[849] : 
                       (N121)? mem[865] : 
                       (N123)? mem[881] : 
                       (N125)? mem[897] : 
                       (N127)? mem[913] : 
                       (N129)? mem[929] : 
                       (N131)? mem[945] : 
                       (N133)? mem[961] : 
                       (N135)? mem[977] : 
                       (N137)? mem[993] : 
                       (N139)? mem[1009] : 1'b0;
  assign r_data_o[0] = (N76)? mem[0] : 
                       (N78)? mem[16] : 
                       (N80)? mem[32] : 
                       (N82)? mem[48] : 
                       (N84)? mem[64] : 
                       (N86)? mem[80] : 
                       (N88)? mem[96] : 
                       (N90)? mem[112] : 
                       (N92)? mem[128] : 
                       (N94)? mem[144] : 
                       (N96)? mem[160] : 
                       (N98)? mem[176] : 
                       (N100)? mem[192] : 
                       (N102)? mem[208] : 
                       (N104)? mem[224] : 
                       (N106)? mem[240] : 
                       (N108)? mem[256] : 
                       (N110)? mem[272] : 
                       (N112)? mem[288] : 
                       (N114)? mem[304] : 
                       (N116)? mem[320] : 
                       (N118)? mem[336] : 
                       (N120)? mem[352] : 
                       (N122)? mem[368] : 
                       (N124)? mem[384] : 
                       (N126)? mem[400] : 
                       (N128)? mem[416] : 
                       (N130)? mem[432] : 
                       (N132)? mem[448] : 
                       (N134)? mem[464] : 
                       (N136)? mem[480] : 
                       (N138)? mem[496] : 
                       (N77)? mem[512] : 
                       (N79)? mem[528] : 
                       (N81)? mem[544] : 
                       (N83)? mem[560] : 
                       (N85)? mem[576] : 
                       (N87)? mem[592] : 
                       (N89)? mem[608] : 
                       (N91)? mem[624] : 
                       (N93)? mem[640] : 
                       (N95)? mem[656] : 
                       (N97)? mem[672] : 
                       (N99)? mem[688] : 
                       (N101)? mem[704] : 
                       (N103)? mem[720] : 
                       (N105)? mem[736] : 
                       (N107)? mem[752] : 
                       (N109)? mem[768] : 
                       (N111)? mem[784] : 
                       (N113)? mem[800] : 
                       (N115)? mem[816] : 
                       (N117)? mem[832] : 
                       (N119)? mem[848] : 
                       (N121)? mem[864] : 
                       (N123)? mem[880] : 
                       (N125)? mem[896] : 
                       (N127)? mem[912] : 
                       (N129)? mem[928] : 
                       (N131)? mem[944] : 
                       (N133)? mem[960] : 
                       (N135)? mem[976] : 
                       (N137)? mem[992] : 
                       (N139)? mem[1008] : 1'b0;
  assign N205 = ~w_addr_i[5];
  assign N206 = w_addr_i[3] & w_addr_i[4];
  assign N207 = N0 & w_addr_i[4];
  assign N0 = ~w_addr_i[3];
  assign N208 = w_addr_i[3] & N1;
  assign N1 = ~w_addr_i[4];
  assign N209 = N2 & N3;
  assign N2 = ~w_addr_i[3];
  assign N3 = ~w_addr_i[4];
  assign N210 = w_addr_i[5] & N206;
  assign N211 = w_addr_i[5] & N207;
  assign N212 = w_addr_i[5] & N208;
  assign N213 = w_addr_i[5] & N209;
  assign N214 = N205 & N206;
  assign N215 = N205 & N207;
  assign N216 = N205 & N208;
  assign N217 = N205 & N209;
  assign N218 = ~w_addr_i[2];
  assign N219 = w_addr_i[0] & w_addr_i[1];
  assign N220 = N4 & w_addr_i[1];
  assign N4 = ~w_addr_i[0];
  assign N221 = w_addr_i[0] & N5;
  assign N5 = ~w_addr_i[1];
  assign N222 = N6 & N7;
  assign N6 = ~w_addr_i[0];
  assign N7 = ~w_addr_i[1];
  assign N223 = w_addr_i[2] & N219;
  assign N224 = w_addr_i[2] & N220;
  assign N225 = w_addr_i[2] & N221;
  assign N226 = w_addr_i[2] & N222;
  assign N227 = N218 & N219;
  assign N228 = N218 & N220;
  assign N229 = N218 & N221;
  assign N230 = N218 & N222;
  assign N231 = N210 & N223;
  assign N232 = N210 & N224;
  assign N233 = N210 & N225;
  assign N234 = N210 & N226;
  assign N235 = N210 & N227;
  assign N236 = N210 & N228;
  assign N237 = N210 & N229;
  assign N238 = N210 & N230;
  assign N239 = N211 & N223;
  assign N240 = N211 & N224;
  assign N241 = N211 & N225;
  assign N242 = N211 & N226;
  assign N243 = N211 & N227;
  assign N244 = N211 & N228;
  assign N245 = N211 & N229;
  assign N246 = N211 & N230;
  assign N247 = N212 & N223;
  assign N248 = N212 & N224;
  assign N249 = N212 & N225;
  assign N250 = N212 & N226;
  assign N251 = N212 & N227;
  assign N252 = N212 & N228;
  assign N253 = N212 & N229;
  assign N254 = N212 & N230;
  assign N255 = N213 & N223;
  assign N256 = N213 & N224;
  assign N257 = N213 & N225;
  assign N258 = N213 & N226;
  assign N259 = N213 & N227;
  assign N260 = N213 & N228;
  assign N261 = N213 & N229;
  assign N262 = N213 & N230;
  assign N263 = N214 & N223;
  assign N264 = N214 & N224;
  assign N265 = N214 & N225;
  assign N266 = N214 & N226;
  assign N267 = N214 & N227;
  assign N268 = N214 & N228;
  assign N269 = N214 & N229;
  assign N270 = N214 & N230;
  assign N271 = N215 & N223;
  assign N272 = N215 & N224;
  assign N273 = N215 & N225;
  assign N274 = N215 & N226;
  assign N275 = N215 & N227;
  assign N276 = N215 & N228;
  assign N277 = N215 & N229;
  assign N278 = N215 & N230;
  assign N279 = N216 & N223;
  assign N280 = N216 & N224;
  assign N281 = N216 & N225;
  assign N282 = N216 & N226;
  assign N283 = N216 & N227;
  assign N284 = N216 & N228;
  assign N285 = N216 & N229;
  assign N286 = N216 & N230;
  assign N287 = N217 & N223;
  assign N288 = N217 & N224;
  assign N289 = N217 & N225;
  assign N290 = N217 & N226;
  assign N291 = N217 & N227;
  assign N292 = N217 & N228;
  assign N293 = N217 & N229;
  assign N294 = N217 & N230;
  assign { N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141 } = (N8)? { N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_v_i;
  assign N9 = N140;
  assign N10 = ~r_addr_i[0];
  assign N11 = ~r_addr_i[1];
  assign N12 = N10 & N11;
  assign N13 = N10 & r_addr_i[1];
  assign N14 = r_addr_i[0] & N11;
  assign N15 = r_addr_i[0] & r_addr_i[1];
  assign N16 = ~r_addr_i[2];
  assign N17 = N12 & N16;
  assign N18 = N12 & r_addr_i[2];
  assign N19 = N14 & N16;
  assign N20 = N14 & r_addr_i[2];
  assign N21 = N13 & N16;
  assign N22 = N13 & r_addr_i[2];
  assign N23 = N15 & N16;
  assign N24 = N15 & r_addr_i[2];
  assign N25 = ~r_addr_i[3];
  assign N26 = N17 & N25;
  assign N27 = N17 & r_addr_i[3];
  assign N28 = N19 & N25;
  assign N29 = N19 & r_addr_i[3];
  assign N30 = N21 & N25;
  assign N31 = N21 & r_addr_i[3];
  assign N32 = N23 & N25;
  assign N33 = N23 & r_addr_i[3];
  assign N34 = N18 & N25;
  assign N35 = N18 & r_addr_i[3];
  assign N36 = N20 & N25;
  assign N37 = N20 & r_addr_i[3];
  assign N38 = N22 & N25;
  assign N39 = N22 & r_addr_i[3];
  assign N40 = N24 & N25;
  assign N41 = N24 & r_addr_i[3];
  assign N42 = ~r_addr_i[4];
  assign N43 = N26 & N42;
  assign N44 = N26 & r_addr_i[4];
  assign N45 = N28 & N42;
  assign N46 = N28 & r_addr_i[4];
  assign N47 = N30 & N42;
  assign N48 = N30 & r_addr_i[4];
  assign N49 = N32 & N42;
  assign N50 = N32 & r_addr_i[4];
  assign N51 = N34 & N42;
  assign N52 = N34 & r_addr_i[4];
  assign N53 = N36 & N42;
  assign N54 = N36 & r_addr_i[4];
  assign N55 = N38 & N42;
  assign N56 = N38 & r_addr_i[4];
  assign N57 = N40 & N42;
  assign N58 = N40 & r_addr_i[4];
  assign N59 = N27 & N42;
  assign N60 = N27 & r_addr_i[4];
  assign N61 = N29 & N42;
  assign N62 = N29 & r_addr_i[4];
  assign N63 = N31 & N42;
  assign N64 = N31 & r_addr_i[4];
  assign N65 = N33 & N42;
  assign N66 = N33 & r_addr_i[4];
  assign N67 = N35 & N42;
  assign N68 = N35 & r_addr_i[4];
  assign N69 = N37 & N42;
  assign N70 = N37 & r_addr_i[4];
  assign N71 = N39 & N42;
  assign N72 = N39 & r_addr_i[4];
  assign N73 = N41 & N42;
  assign N74 = N41 & r_addr_i[4];
  assign N75 = ~r_addr_i[5];
  assign N76 = N43 & N75;
  assign N77 = N43 & r_addr_i[5];
  assign N78 = N45 & N75;
  assign N79 = N45 & r_addr_i[5];
  assign N80 = N47 & N75;
  assign N81 = N47 & r_addr_i[5];
  assign N82 = N49 & N75;
  assign N83 = N49 & r_addr_i[5];
  assign N84 = N51 & N75;
  assign N85 = N51 & r_addr_i[5];
  assign N86 = N53 & N75;
  assign N87 = N53 & r_addr_i[5];
  assign N88 = N55 & N75;
  assign N89 = N55 & r_addr_i[5];
  assign N90 = N57 & N75;
  assign N91 = N57 & r_addr_i[5];
  assign N92 = N59 & N75;
  assign N93 = N59 & r_addr_i[5];
  assign N94 = N61 & N75;
  assign N95 = N61 & r_addr_i[5];
  assign N96 = N63 & N75;
  assign N97 = N63 & r_addr_i[5];
  assign N98 = N65 & N75;
  assign N99 = N65 & r_addr_i[5];
  assign N100 = N67 & N75;
  assign N101 = N67 & r_addr_i[5];
  assign N102 = N69 & N75;
  assign N103 = N69 & r_addr_i[5];
  assign N104 = N71 & N75;
  assign N105 = N71 & r_addr_i[5];
  assign N106 = N73 & N75;
  assign N107 = N73 & r_addr_i[5];
  assign N108 = N44 & N75;
  assign N109 = N44 & r_addr_i[5];
  assign N110 = N46 & N75;
  assign N111 = N46 & r_addr_i[5];
  assign N112 = N48 & N75;
  assign N113 = N48 & r_addr_i[5];
  assign N114 = N50 & N75;
  assign N115 = N50 & r_addr_i[5];
  assign N116 = N52 & N75;
  assign N117 = N52 & r_addr_i[5];
  assign N118 = N54 & N75;
  assign N119 = N54 & r_addr_i[5];
  assign N120 = N56 & N75;
  assign N121 = N56 & r_addr_i[5];
  assign N122 = N58 & N75;
  assign N123 = N58 & r_addr_i[5];
  assign N124 = N60 & N75;
  assign N125 = N60 & r_addr_i[5];
  assign N126 = N62 & N75;
  assign N127 = N62 & r_addr_i[5];
  assign N128 = N64 & N75;
  assign N129 = N64 & r_addr_i[5];
  assign N130 = N66 & N75;
  assign N131 = N66 & r_addr_i[5];
  assign N132 = N68 & N75;
  assign N133 = N68 & r_addr_i[5];
  assign N134 = N70 & N75;
  assign N135 = N70 & r_addr_i[5];
  assign N136 = N72 & N75;
  assign N137 = N72 & r_addr_i[5];
  assign N138 = N74 & N75;
  assign N139 = N74 & r_addr_i[5];
  assign N140 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N204) begin
      mem_1023_sv2v_reg <= w_data_i[15];
      mem_1022_sv2v_reg <= w_data_i[14];
      mem_1021_sv2v_reg <= w_data_i[13];
      mem_1020_sv2v_reg <= w_data_i[12];
      mem_1019_sv2v_reg <= w_data_i[11];
      mem_1018_sv2v_reg <= w_data_i[10];
      mem_1017_sv2v_reg <= w_data_i[9];
      mem_1016_sv2v_reg <= w_data_i[8];
      mem_1015_sv2v_reg <= w_data_i[7];
      mem_1014_sv2v_reg <= w_data_i[6];
      mem_1013_sv2v_reg <= w_data_i[5];
      mem_1012_sv2v_reg <= w_data_i[4];
      mem_1011_sv2v_reg <= w_data_i[3];
      mem_1010_sv2v_reg <= w_data_i[2];
      mem_1009_sv2v_reg <= w_data_i[1];
      mem_1008_sv2v_reg <= w_data_i[0];
    end 
    if(N203) begin
      mem_1007_sv2v_reg <= w_data_i[15];
      mem_1006_sv2v_reg <= w_data_i[14];
      mem_1005_sv2v_reg <= w_data_i[13];
      mem_1004_sv2v_reg <= w_data_i[12];
      mem_1003_sv2v_reg <= w_data_i[11];
      mem_1002_sv2v_reg <= w_data_i[10];
      mem_1001_sv2v_reg <= w_data_i[9];
      mem_1000_sv2v_reg <= w_data_i[8];
      mem_999_sv2v_reg <= w_data_i[7];
      mem_998_sv2v_reg <= w_data_i[6];
      mem_997_sv2v_reg <= w_data_i[5];
      mem_996_sv2v_reg <= w_data_i[4];
      mem_995_sv2v_reg <= w_data_i[3];
      mem_994_sv2v_reg <= w_data_i[2];
      mem_993_sv2v_reg <= w_data_i[1];
      mem_992_sv2v_reg <= w_data_i[0];
    end 
    if(N202) begin
      mem_991_sv2v_reg <= w_data_i[15];
      mem_990_sv2v_reg <= w_data_i[14];
      mem_989_sv2v_reg <= w_data_i[13];
      mem_988_sv2v_reg <= w_data_i[12];
      mem_987_sv2v_reg <= w_data_i[11];
      mem_986_sv2v_reg <= w_data_i[10];
      mem_985_sv2v_reg <= w_data_i[9];
      mem_984_sv2v_reg <= w_data_i[8];
      mem_983_sv2v_reg <= w_data_i[7];
      mem_982_sv2v_reg <= w_data_i[6];
      mem_981_sv2v_reg <= w_data_i[5];
      mem_980_sv2v_reg <= w_data_i[4];
      mem_979_sv2v_reg <= w_data_i[3];
      mem_978_sv2v_reg <= w_data_i[2];
      mem_977_sv2v_reg <= w_data_i[1];
      mem_976_sv2v_reg <= w_data_i[0];
    end 
    if(N201) begin
      mem_975_sv2v_reg <= w_data_i[15];
      mem_974_sv2v_reg <= w_data_i[14];
      mem_973_sv2v_reg <= w_data_i[13];
      mem_972_sv2v_reg <= w_data_i[12];
      mem_971_sv2v_reg <= w_data_i[11];
      mem_970_sv2v_reg <= w_data_i[10];
      mem_969_sv2v_reg <= w_data_i[9];
      mem_968_sv2v_reg <= w_data_i[8];
      mem_967_sv2v_reg <= w_data_i[7];
      mem_966_sv2v_reg <= w_data_i[6];
      mem_965_sv2v_reg <= w_data_i[5];
      mem_964_sv2v_reg <= w_data_i[4];
      mem_963_sv2v_reg <= w_data_i[3];
      mem_962_sv2v_reg <= w_data_i[2];
      mem_961_sv2v_reg <= w_data_i[1];
      mem_960_sv2v_reg <= w_data_i[0];
    end 
    if(N200) begin
      mem_959_sv2v_reg <= w_data_i[15];
      mem_958_sv2v_reg <= w_data_i[14];
      mem_957_sv2v_reg <= w_data_i[13];
      mem_956_sv2v_reg <= w_data_i[12];
      mem_955_sv2v_reg <= w_data_i[11];
      mem_954_sv2v_reg <= w_data_i[10];
      mem_953_sv2v_reg <= w_data_i[9];
      mem_952_sv2v_reg <= w_data_i[8];
      mem_951_sv2v_reg <= w_data_i[7];
      mem_950_sv2v_reg <= w_data_i[6];
      mem_949_sv2v_reg <= w_data_i[5];
      mem_948_sv2v_reg <= w_data_i[4];
      mem_947_sv2v_reg <= w_data_i[3];
      mem_946_sv2v_reg <= w_data_i[2];
      mem_945_sv2v_reg <= w_data_i[1];
      mem_944_sv2v_reg <= w_data_i[0];
    end 
    if(N199) begin
      mem_943_sv2v_reg <= w_data_i[15];
      mem_942_sv2v_reg <= w_data_i[14];
      mem_941_sv2v_reg <= w_data_i[13];
      mem_940_sv2v_reg <= w_data_i[12];
      mem_939_sv2v_reg <= w_data_i[11];
      mem_938_sv2v_reg <= w_data_i[10];
      mem_937_sv2v_reg <= w_data_i[9];
      mem_936_sv2v_reg <= w_data_i[8];
      mem_935_sv2v_reg <= w_data_i[7];
      mem_934_sv2v_reg <= w_data_i[6];
      mem_933_sv2v_reg <= w_data_i[5];
      mem_932_sv2v_reg <= w_data_i[4];
      mem_931_sv2v_reg <= w_data_i[3];
      mem_930_sv2v_reg <= w_data_i[2];
      mem_929_sv2v_reg <= w_data_i[1];
      mem_928_sv2v_reg <= w_data_i[0];
    end 
    if(N198) begin
      mem_927_sv2v_reg <= w_data_i[15];
      mem_926_sv2v_reg <= w_data_i[14];
      mem_925_sv2v_reg <= w_data_i[13];
      mem_924_sv2v_reg <= w_data_i[12];
      mem_923_sv2v_reg <= w_data_i[11];
      mem_922_sv2v_reg <= w_data_i[10];
      mem_921_sv2v_reg <= w_data_i[9];
      mem_920_sv2v_reg <= w_data_i[8];
      mem_919_sv2v_reg <= w_data_i[7];
      mem_918_sv2v_reg <= w_data_i[6];
      mem_917_sv2v_reg <= w_data_i[5];
      mem_916_sv2v_reg <= w_data_i[4];
      mem_915_sv2v_reg <= w_data_i[3];
      mem_914_sv2v_reg <= w_data_i[2];
      mem_913_sv2v_reg <= w_data_i[1];
      mem_912_sv2v_reg <= w_data_i[0];
    end 
    if(N197) begin
      mem_911_sv2v_reg <= w_data_i[15];
      mem_910_sv2v_reg <= w_data_i[14];
      mem_909_sv2v_reg <= w_data_i[13];
      mem_908_sv2v_reg <= w_data_i[12];
      mem_907_sv2v_reg <= w_data_i[11];
      mem_906_sv2v_reg <= w_data_i[10];
      mem_905_sv2v_reg <= w_data_i[9];
      mem_904_sv2v_reg <= w_data_i[8];
      mem_903_sv2v_reg <= w_data_i[7];
      mem_902_sv2v_reg <= w_data_i[6];
      mem_901_sv2v_reg <= w_data_i[5];
      mem_900_sv2v_reg <= w_data_i[4];
      mem_899_sv2v_reg <= w_data_i[3];
      mem_898_sv2v_reg <= w_data_i[2];
      mem_897_sv2v_reg <= w_data_i[1];
      mem_896_sv2v_reg <= w_data_i[0];
    end 
    if(N196) begin
      mem_895_sv2v_reg <= w_data_i[15];
      mem_894_sv2v_reg <= w_data_i[14];
      mem_893_sv2v_reg <= w_data_i[13];
      mem_892_sv2v_reg <= w_data_i[12];
      mem_891_sv2v_reg <= w_data_i[11];
      mem_890_sv2v_reg <= w_data_i[10];
      mem_889_sv2v_reg <= w_data_i[9];
      mem_888_sv2v_reg <= w_data_i[8];
      mem_887_sv2v_reg <= w_data_i[7];
      mem_886_sv2v_reg <= w_data_i[6];
      mem_885_sv2v_reg <= w_data_i[5];
      mem_884_sv2v_reg <= w_data_i[4];
      mem_883_sv2v_reg <= w_data_i[3];
      mem_882_sv2v_reg <= w_data_i[2];
      mem_881_sv2v_reg <= w_data_i[1];
      mem_880_sv2v_reg <= w_data_i[0];
    end 
    if(N195) begin
      mem_879_sv2v_reg <= w_data_i[15];
      mem_878_sv2v_reg <= w_data_i[14];
      mem_877_sv2v_reg <= w_data_i[13];
      mem_876_sv2v_reg <= w_data_i[12];
      mem_875_sv2v_reg <= w_data_i[11];
      mem_874_sv2v_reg <= w_data_i[10];
      mem_873_sv2v_reg <= w_data_i[9];
      mem_872_sv2v_reg <= w_data_i[8];
      mem_871_sv2v_reg <= w_data_i[7];
      mem_870_sv2v_reg <= w_data_i[6];
      mem_869_sv2v_reg <= w_data_i[5];
      mem_868_sv2v_reg <= w_data_i[4];
      mem_867_sv2v_reg <= w_data_i[3];
      mem_866_sv2v_reg <= w_data_i[2];
      mem_865_sv2v_reg <= w_data_i[1];
      mem_864_sv2v_reg <= w_data_i[0];
    end 
    if(N194) begin
      mem_863_sv2v_reg <= w_data_i[15];
      mem_862_sv2v_reg <= w_data_i[14];
      mem_861_sv2v_reg <= w_data_i[13];
      mem_860_sv2v_reg <= w_data_i[12];
      mem_859_sv2v_reg <= w_data_i[11];
      mem_858_sv2v_reg <= w_data_i[10];
      mem_857_sv2v_reg <= w_data_i[9];
      mem_856_sv2v_reg <= w_data_i[8];
      mem_855_sv2v_reg <= w_data_i[7];
      mem_854_sv2v_reg <= w_data_i[6];
      mem_853_sv2v_reg <= w_data_i[5];
      mem_852_sv2v_reg <= w_data_i[4];
      mem_851_sv2v_reg <= w_data_i[3];
      mem_850_sv2v_reg <= w_data_i[2];
      mem_849_sv2v_reg <= w_data_i[1];
      mem_848_sv2v_reg <= w_data_i[0];
    end 
    if(N193) begin
      mem_847_sv2v_reg <= w_data_i[15];
      mem_846_sv2v_reg <= w_data_i[14];
      mem_845_sv2v_reg <= w_data_i[13];
      mem_844_sv2v_reg <= w_data_i[12];
      mem_843_sv2v_reg <= w_data_i[11];
      mem_842_sv2v_reg <= w_data_i[10];
      mem_841_sv2v_reg <= w_data_i[9];
      mem_840_sv2v_reg <= w_data_i[8];
      mem_839_sv2v_reg <= w_data_i[7];
      mem_838_sv2v_reg <= w_data_i[6];
      mem_837_sv2v_reg <= w_data_i[5];
      mem_836_sv2v_reg <= w_data_i[4];
      mem_835_sv2v_reg <= w_data_i[3];
      mem_834_sv2v_reg <= w_data_i[2];
      mem_833_sv2v_reg <= w_data_i[1];
      mem_832_sv2v_reg <= w_data_i[0];
    end 
    if(N192) begin
      mem_831_sv2v_reg <= w_data_i[15];
      mem_830_sv2v_reg <= w_data_i[14];
      mem_829_sv2v_reg <= w_data_i[13];
      mem_828_sv2v_reg <= w_data_i[12];
      mem_827_sv2v_reg <= w_data_i[11];
      mem_826_sv2v_reg <= w_data_i[10];
      mem_825_sv2v_reg <= w_data_i[9];
      mem_824_sv2v_reg <= w_data_i[8];
      mem_823_sv2v_reg <= w_data_i[7];
      mem_822_sv2v_reg <= w_data_i[6];
      mem_821_sv2v_reg <= w_data_i[5];
      mem_820_sv2v_reg <= w_data_i[4];
      mem_819_sv2v_reg <= w_data_i[3];
      mem_818_sv2v_reg <= w_data_i[2];
      mem_817_sv2v_reg <= w_data_i[1];
      mem_816_sv2v_reg <= w_data_i[0];
    end 
    if(N191) begin
      mem_815_sv2v_reg <= w_data_i[15];
      mem_814_sv2v_reg <= w_data_i[14];
      mem_813_sv2v_reg <= w_data_i[13];
      mem_812_sv2v_reg <= w_data_i[12];
      mem_811_sv2v_reg <= w_data_i[11];
      mem_810_sv2v_reg <= w_data_i[10];
      mem_809_sv2v_reg <= w_data_i[9];
      mem_808_sv2v_reg <= w_data_i[8];
      mem_807_sv2v_reg <= w_data_i[7];
      mem_806_sv2v_reg <= w_data_i[6];
      mem_805_sv2v_reg <= w_data_i[5];
      mem_804_sv2v_reg <= w_data_i[4];
      mem_803_sv2v_reg <= w_data_i[3];
      mem_802_sv2v_reg <= w_data_i[2];
      mem_801_sv2v_reg <= w_data_i[1];
      mem_800_sv2v_reg <= w_data_i[0];
    end 
    if(N190) begin
      mem_799_sv2v_reg <= w_data_i[15];
      mem_798_sv2v_reg <= w_data_i[14];
      mem_797_sv2v_reg <= w_data_i[13];
      mem_796_sv2v_reg <= w_data_i[12];
      mem_795_sv2v_reg <= w_data_i[11];
      mem_794_sv2v_reg <= w_data_i[10];
      mem_793_sv2v_reg <= w_data_i[9];
      mem_792_sv2v_reg <= w_data_i[8];
      mem_791_sv2v_reg <= w_data_i[7];
      mem_790_sv2v_reg <= w_data_i[6];
      mem_789_sv2v_reg <= w_data_i[5];
      mem_788_sv2v_reg <= w_data_i[4];
      mem_787_sv2v_reg <= w_data_i[3];
      mem_786_sv2v_reg <= w_data_i[2];
      mem_785_sv2v_reg <= w_data_i[1];
      mem_784_sv2v_reg <= w_data_i[0];
    end 
    if(N189) begin
      mem_783_sv2v_reg <= w_data_i[15];
      mem_782_sv2v_reg <= w_data_i[14];
      mem_781_sv2v_reg <= w_data_i[13];
      mem_780_sv2v_reg <= w_data_i[12];
      mem_779_sv2v_reg <= w_data_i[11];
      mem_778_sv2v_reg <= w_data_i[10];
      mem_777_sv2v_reg <= w_data_i[9];
      mem_776_sv2v_reg <= w_data_i[8];
      mem_775_sv2v_reg <= w_data_i[7];
      mem_774_sv2v_reg <= w_data_i[6];
      mem_773_sv2v_reg <= w_data_i[5];
      mem_772_sv2v_reg <= w_data_i[4];
      mem_771_sv2v_reg <= w_data_i[3];
      mem_770_sv2v_reg <= w_data_i[2];
      mem_769_sv2v_reg <= w_data_i[1];
      mem_768_sv2v_reg <= w_data_i[0];
    end 
    if(N188) begin
      mem_767_sv2v_reg <= w_data_i[15];
      mem_766_sv2v_reg <= w_data_i[14];
      mem_765_sv2v_reg <= w_data_i[13];
      mem_764_sv2v_reg <= w_data_i[12];
      mem_763_sv2v_reg <= w_data_i[11];
      mem_762_sv2v_reg <= w_data_i[10];
      mem_761_sv2v_reg <= w_data_i[9];
      mem_760_sv2v_reg <= w_data_i[8];
      mem_759_sv2v_reg <= w_data_i[7];
      mem_758_sv2v_reg <= w_data_i[6];
      mem_757_sv2v_reg <= w_data_i[5];
      mem_756_sv2v_reg <= w_data_i[4];
      mem_755_sv2v_reg <= w_data_i[3];
      mem_754_sv2v_reg <= w_data_i[2];
      mem_753_sv2v_reg <= w_data_i[1];
      mem_752_sv2v_reg <= w_data_i[0];
    end 
    if(N187) begin
      mem_751_sv2v_reg <= w_data_i[15];
      mem_750_sv2v_reg <= w_data_i[14];
      mem_749_sv2v_reg <= w_data_i[13];
      mem_748_sv2v_reg <= w_data_i[12];
      mem_747_sv2v_reg <= w_data_i[11];
      mem_746_sv2v_reg <= w_data_i[10];
      mem_745_sv2v_reg <= w_data_i[9];
      mem_744_sv2v_reg <= w_data_i[8];
      mem_743_sv2v_reg <= w_data_i[7];
      mem_742_sv2v_reg <= w_data_i[6];
      mem_741_sv2v_reg <= w_data_i[5];
      mem_740_sv2v_reg <= w_data_i[4];
      mem_739_sv2v_reg <= w_data_i[3];
      mem_738_sv2v_reg <= w_data_i[2];
      mem_737_sv2v_reg <= w_data_i[1];
      mem_736_sv2v_reg <= w_data_i[0];
    end 
    if(N186) begin
      mem_735_sv2v_reg <= w_data_i[15];
      mem_734_sv2v_reg <= w_data_i[14];
      mem_733_sv2v_reg <= w_data_i[13];
      mem_732_sv2v_reg <= w_data_i[12];
      mem_731_sv2v_reg <= w_data_i[11];
      mem_730_sv2v_reg <= w_data_i[10];
      mem_729_sv2v_reg <= w_data_i[9];
      mem_728_sv2v_reg <= w_data_i[8];
      mem_727_sv2v_reg <= w_data_i[7];
      mem_726_sv2v_reg <= w_data_i[6];
      mem_725_sv2v_reg <= w_data_i[5];
      mem_724_sv2v_reg <= w_data_i[4];
      mem_723_sv2v_reg <= w_data_i[3];
      mem_722_sv2v_reg <= w_data_i[2];
      mem_721_sv2v_reg <= w_data_i[1];
      mem_720_sv2v_reg <= w_data_i[0];
    end 
    if(N185) begin
      mem_719_sv2v_reg <= w_data_i[15];
      mem_718_sv2v_reg <= w_data_i[14];
      mem_717_sv2v_reg <= w_data_i[13];
      mem_716_sv2v_reg <= w_data_i[12];
      mem_715_sv2v_reg <= w_data_i[11];
      mem_714_sv2v_reg <= w_data_i[10];
      mem_713_sv2v_reg <= w_data_i[9];
      mem_712_sv2v_reg <= w_data_i[8];
      mem_711_sv2v_reg <= w_data_i[7];
      mem_710_sv2v_reg <= w_data_i[6];
      mem_709_sv2v_reg <= w_data_i[5];
      mem_708_sv2v_reg <= w_data_i[4];
      mem_707_sv2v_reg <= w_data_i[3];
      mem_706_sv2v_reg <= w_data_i[2];
      mem_705_sv2v_reg <= w_data_i[1];
      mem_704_sv2v_reg <= w_data_i[0];
    end 
    if(N184) begin
      mem_703_sv2v_reg <= w_data_i[15];
      mem_702_sv2v_reg <= w_data_i[14];
      mem_701_sv2v_reg <= w_data_i[13];
      mem_700_sv2v_reg <= w_data_i[12];
      mem_699_sv2v_reg <= w_data_i[11];
      mem_698_sv2v_reg <= w_data_i[10];
      mem_697_sv2v_reg <= w_data_i[9];
      mem_696_sv2v_reg <= w_data_i[8];
      mem_695_sv2v_reg <= w_data_i[7];
      mem_694_sv2v_reg <= w_data_i[6];
      mem_693_sv2v_reg <= w_data_i[5];
      mem_692_sv2v_reg <= w_data_i[4];
      mem_691_sv2v_reg <= w_data_i[3];
      mem_690_sv2v_reg <= w_data_i[2];
      mem_689_sv2v_reg <= w_data_i[1];
      mem_688_sv2v_reg <= w_data_i[0];
    end 
    if(N183) begin
      mem_687_sv2v_reg <= w_data_i[15];
      mem_686_sv2v_reg <= w_data_i[14];
      mem_685_sv2v_reg <= w_data_i[13];
      mem_684_sv2v_reg <= w_data_i[12];
      mem_683_sv2v_reg <= w_data_i[11];
      mem_682_sv2v_reg <= w_data_i[10];
      mem_681_sv2v_reg <= w_data_i[9];
      mem_680_sv2v_reg <= w_data_i[8];
      mem_679_sv2v_reg <= w_data_i[7];
      mem_678_sv2v_reg <= w_data_i[6];
      mem_677_sv2v_reg <= w_data_i[5];
      mem_676_sv2v_reg <= w_data_i[4];
      mem_675_sv2v_reg <= w_data_i[3];
      mem_674_sv2v_reg <= w_data_i[2];
      mem_673_sv2v_reg <= w_data_i[1];
      mem_672_sv2v_reg <= w_data_i[0];
    end 
    if(N182) begin
      mem_671_sv2v_reg <= w_data_i[15];
      mem_670_sv2v_reg <= w_data_i[14];
      mem_669_sv2v_reg <= w_data_i[13];
      mem_668_sv2v_reg <= w_data_i[12];
      mem_667_sv2v_reg <= w_data_i[11];
      mem_666_sv2v_reg <= w_data_i[10];
      mem_665_sv2v_reg <= w_data_i[9];
      mem_664_sv2v_reg <= w_data_i[8];
      mem_663_sv2v_reg <= w_data_i[7];
      mem_662_sv2v_reg <= w_data_i[6];
      mem_661_sv2v_reg <= w_data_i[5];
      mem_660_sv2v_reg <= w_data_i[4];
      mem_659_sv2v_reg <= w_data_i[3];
      mem_658_sv2v_reg <= w_data_i[2];
      mem_657_sv2v_reg <= w_data_i[1];
      mem_656_sv2v_reg <= w_data_i[0];
    end 
    if(N181) begin
      mem_655_sv2v_reg <= w_data_i[15];
      mem_654_sv2v_reg <= w_data_i[14];
      mem_653_sv2v_reg <= w_data_i[13];
      mem_652_sv2v_reg <= w_data_i[12];
      mem_651_sv2v_reg <= w_data_i[11];
      mem_650_sv2v_reg <= w_data_i[10];
      mem_649_sv2v_reg <= w_data_i[9];
      mem_648_sv2v_reg <= w_data_i[8];
      mem_647_sv2v_reg <= w_data_i[7];
      mem_646_sv2v_reg <= w_data_i[6];
      mem_645_sv2v_reg <= w_data_i[5];
      mem_644_sv2v_reg <= w_data_i[4];
      mem_643_sv2v_reg <= w_data_i[3];
      mem_642_sv2v_reg <= w_data_i[2];
      mem_641_sv2v_reg <= w_data_i[1];
      mem_640_sv2v_reg <= w_data_i[0];
    end 
    if(N180) begin
      mem_639_sv2v_reg <= w_data_i[15];
      mem_638_sv2v_reg <= w_data_i[14];
      mem_637_sv2v_reg <= w_data_i[13];
      mem_636_sv2v_reg <= w_data_i[12];
      mem_635_sv2v_reg <= w_data_i[11];
      mem_634_sv2v_reg <= w_data_i[10];
      mem_633_sv2v_reg <= w_data_i[9];
      mem_632_sv2v_reg <= w_data_i[8];
      mem_631_sv2v_reg <= w_data_i[7];
      mem_630_sv2v_reg <= w_data_i[6];
      mem_629_sv2v_reg <= w_data_i[5];
      mem_628_sv2v_reg <= w_data_i[4];
      mem_627_sv2v_reg <= w_data_i[3];
      mem_626_sv2v_reg <= w_data_i[2];
      mem_625_sv2v_reg <= w_data_i[1];
      mem_624_sv2v_reg <= w_data_i[0];
    end 
    if(N179) begin
      mem_623_sv2v_reg <= w_data_i[15];
      mem_622_sv2v_reg <= w_data_i[14];
      mem_621_sv2v_reg <= w_data_i[13];
      mem_620_sv2v_reg <= w_data_i[12];
      mem_619_sv2v_reg <= w_data_i[11];
      mem_618_sv2v_reg <= w_data_i[10];
      mem_617_sv2v_reg <= w_data_i[9];
      mem_616_sv2v_reg <= w_data_i[8];
      mem_615_sv2v_reg <= w_data_i[7];
      mem_614_sv2v_reg <= w_data_i[6];
      mem_613_sv2v_reg <= w_data_i[5];
      mem_612_sv2v_reg <= w_data_i[4];
      mem_611_sv2v_reg <= w_data_i[3];
      mem_610_sv2v_reg <= w_data_i[2];
      mem_609_sv2v_reg <= w_data_i[1];
      mem_608_sv2v_reg <= w_data_i[0];
    end 
    if(N178) begin
      mem_607_sv2v_reg <= w_data_i[15];
      mem_606_sv2v_reg <= w_data_i[14];
      mem_605_sv2v_reg <= w_data_i[13];
      mem_604_sv2v_reg <= w_data_i[12];
      mem_603_sv2v_reg <= w_data_i[11];
      mem_602_sv2v_reg <= w_data_i[10];
      mem_601_sv2v_reg <= w_data_i[9];
      mem_600_sv2v_reg <= w_data_i[8];
      mem_599_sv2v_reg <= w_data_i[7];
      mem_598_sv2v_reg <= w_data_i[6];
      mem_597_sv2v_reg <= w_data_i[5];
      mem_596_sv2v_reg <= w_data_i[4];
      mem_595_sv2v_reg <= w_data_i[3];
      mem_594_sv2v_reg <= w_data_i[2];
      mem_593_sv2v_reg <= w_data_i[1];
      mem_592_sv2v_reg <= w_data_i[0];
    end 
    if(N177) begin
      mem_591_sv2v_reg <= w_data_i[15];
      mem_590_sv2v_reg <= w_data_i[14];
      mem_589_sv2v_reg <= w_data_i[13];
      mem_588_sv2v_reg <= w_data_i[12];
      mem_587_sv2v_reg <= w_data_i[11];
      mem_586_sv2v_reg <= w_data_i[10];
      mem_585_sv2v_reg <= w_data_i[9];
      mem_584_sv2v_reg <= w_data_i[8];
      mem_583_sv2v_reg <= w_data_i[7];
      mem_582_sv2v_reg <= w_data_i[6];
      mem_581_sv2v_reg <= w_data_i[5];
      mem_580_sv2v_reg <= w_data_i[4];
      mem_579_sv2v_reg <= w_data_i[3];
      mem_578_sv2v_reg <= w_data_i[2];
      mem_577_sv2v_reg <= w_data_i[1];
      mem_576_sv2v_reg <= w_data_i[0];
    end 
    if(N176) begin
      mem_575_sv2v_reg <= w_data_i[15];
      mem_574_sv2v_reg <= w_data_i[14];
      mem_573_sv2v_reg <= w_data_i[13];
      mem_572_sv2v_reg <= w_data_i[12];
      mem_571_sv2v_reg <= w_data_i[11];
      mem_570_sv2v_reg <= w_data_i[10];
      mem_569_sv2v_reg <= w_data_i[9];
      mem_568_sv2v_reg <= w_data_i[8];
      mem_567_sv2v_reg <= w_data_i[7];
      mem_566_sv2v_reg <= w_data_i[6];
      mem_565_sv2v_reg <= w_data_i[5];
      mem_564_sv2v_reg <= w_data_i[4];
      mem_563_sv2v_reg <= w_data_i[3];
      mem_562_sv2v_reg <= w_data_i[2];
      mem_561_sv2v_reg <= w_data_i[1];
      mem_560_sv2v_reg <= w_data_i[0];
    end 
    if(N175) begin
      mem_559_sv2v_reg <= w_data_i[15];
      mem_558_sv2v_reg <= w_data_i[14];
      mem_557_sv2v_reg <= w_data_i[13];
      mem_556_sv2v_reg <= w_data_i[12];
      mem_555_sv2v_reg <= w_data_i[11];
      mem_554_sv2v_reg <= w_data_i[10];
      mem_553_sv2v_reg <= w_data_i[9];
      mem_552_sv2v_reg <= w_data_i[8];
      mem_551_sv2v_reg <= w_data_i[7];
      mem_550_sv2v_reg <= w_data_i[6];
      mem_549_sv2v_reg <= w_data_i[5];
      mem_548_sv2v_reg <= w_data_i[4];
      mem_547_sv2v_reg <= w_data_i[3];
      mem_546_sv2v_reg <= w_data_i[2];
      mem_545_sv2v_reg <= w_data_i[1];
      mem_544_sv2v_reg <= w_data_i[0];
    end 
    if(N174) begin
      mem_543_sv2v_reg <= w_data_i[15];
      mem_542_sv2v_reg <= w_data_i[14];
      mem_541_sv2v_reg <= w_data_i[13];
      mem_540_sv2v_reg <= w_data_i[12];
      mem_539_sv2v_reg <= w_data_i[11];
      mem_538_sv2v_reg <= w_data_i[10];
      mem_537_sv2v_reg <= w_data_i[9];
      mem_536_sv2v_reg <= w_data_i[8];
      mem_535_sv2v_reg <= w_data_i[7];
      mem_534_sv2v_reg <= w_data_i[6];
      mem_533_sv2v_reg <= w_data_i[5];
      mem_532_sv2v_reg <= w_data_i[4];
      mem_531_sv2v_reg <= w_data_i[3];
      mem_530_sv2v_reg <= w_data_i[2];
      mem_529_sv2v_reg <= w_data_i[1];
      mem_528_sv2v_reg <= w_data_i[0];
    end 
    if(N173) begin
      mem_527_sv2v_reg <= w_data_i[15];
      mem_526_sv2v_reg <= w_data_i[14];
      mem_525_sv2v_reg <= w_data_i[13];
      mem_524_sv2v_reg <= w_data_i[12];
      mem_523_sv2v_reg <= w_data_i[11];
      mem_522_sv2v_reg <= w_data_i[10];
      mem_521_sv2v_reg <= w_data_i[9];
      mem_520_sv2v_reg <= w_data_i[8];
      mem_519_sv2v_reg <= w_data_i[7];
      mem_518_sv2v_reg <= w_data_i[6];
      mem_517_sv2v_reg <= w_data_i[5];
      mem_516_sv2v_reg <= w_data_i[4];
      mem_515_sv2v_reg <= w_data_i[3];
      mem_514_sv2v_reg <= w_data_i[2];
      mem_513_sv2v_reg <= w_data_i[1];
      mem_512_sv2v_reg <= w_data_i[0];
    end 
    if(N172) begin
      mem_511_sv2v_reg <= w_data_i[15];
      mem_510_sv2v_reg <= w_data_i[14];
      mem_509_sv2v_reg <= w_data_i[13];
      mem_508_sv2v_reg <= w_data_i[12];
      mem_507_sv2v_reg <= w_data_i[11];
      mem_506_sv2v_reg <= w_data_i[10];
      mem_505_sv2v_reg <= w_data_i[9];
      mem_504_sv2v_reg <= w_data_i[8];
      mem_503_sv2v_reg <= w_data_i[7];
      mem_502_sv2v_reg <= w_data_i[6];
      mem_501_sv2v_reg <= w_data_i[5];
      mem_500_sv2v_reg <= w_data_i[4];
      mem_499_sv2v_reg <= w_data_i[3];
      mem_498_sv2v_reg <= w_data_i[2];
      mem_497_sv2v_reg <= w_data_i[1];
      mem_496_sv2v_reg <= w_data_i[0];
    end 
    if(N171) begin
      mem_495_sv2v_reg <= w_data_i[15];
      mem_494_sv2v_reg <= w_data_i[14];
      mem_493_sv2v_reg <= w_data_i[13];
      mem_492_sv2v_reg <= w_data_i[12];
      mem_491_sv2v_reg <= w_data_i[11];
      mem_490_sv2v_reg <= w_data_i[10];
      mem_489_sv2v_reg <= w_data_i[9];
      mem_488_sv2v_reg <= w_data_i[8];
      mem_487_sv2v_reg <= w_data_i[7];
      mem_486_sv2v_reg <= w_data_i[6];
      mem_485_sv2v_reg <= w_data_i[5];
      mem_484_sv2v_reg <= w_data_i[4];
      mem_483_sv2v_reg <= w_data_i[3];
      mem_482_sv2v_reg <= w_data_i[2];
      mem_481_sv2v_reg <= w_data_i[1];
      mem_480_sv2v_reg <= w_data_i[0];
    end 
    if(N170) begin
      mem_479_sv2v_reg <= w_data_i[15];
      mem_478_sv2v_reg <= w_data_i[14];
      mem_477_sv2v_reg <= w_data_i[13];
      mem_476_sv2v_reg <= w_data_i[12];
      mem_475_sv2v_reg <= w_data_i[11];
      mem_474_sv2v_reg <= w_data_i[10];
      mem_473_sv2v_reg <= w_data_i[9];
      mem_472_sv2v_reg <= w_data_i[8];
      mem_471_sv2v_reg <= w_data_i[7];
      mem_470_sv2v_reg <= w_data_i[6];
      mem_469_sv2v_reg <= w_data_i[5];
      mem_468_sv2v_reg <= w_data_i[4];
      mem_467_sv2v_reg <= w_data_i[3];
      mem_466_sv2v_reg <= w_data_i[2];
      mem_465_sv2v_reg <= w_data_i[1];
      mem_464_sv2v_reg <= w_data_i[0];
    end 
    if(N169) begin
      mem_463_sv2v_reg <= w_data_i[15];
      mem_462_sv2v_reg <= w_data_i[14];
      mem_461_sv2v_reg <= w_data_i[13];
      mem_460_sv2v_reg <= w_data_i[12];
      mem_459_sv2v_reg <= w_data_i[11];
      mem_458_sv2v_reg <= w_data_i[10];
      mem_457_sv2v_reg <= w_data_i[9];
      mem_456_sv2v_reg <= w_data_i[8];
      mem_455_sv2v_reg <= w_data_i[7];
      mem_454_sv2v_reg <= w_data_i[6];
      mem_453_sv2v_reg <= w_data_i[5];
      mem_452_sv2v_reg <= w_data_i[4];
      mem_451_sv2v_reg <= w_data_i[3];
      mem_450_sv2v_reg <= w_data_i[2];
      mem_449_sv2v_reg <= w_data_i[1];
      mem_448_sv2v_reg <= w_data_i[0];
    end 
    if(N168) begin
      mem_447_sv2v_reg <= w_data_i[15];
      mem_446_sv2v_reg <= w_data_i[14];
      mem_445_sv2v_reg <= w_data_i[13];
      mem_444_sv2v_reg <= w_data_i[12];
      mem_443_sv2v_reg <= w_data_i[11];
      mem_442_sv2v_reg <= w_data_i[10];
      mem_441_sv2v_reg <= w_data_i[9];
      mem_440_sv2v_reg <= w_data_i[8];
      mem_439_sv2v_reg <= w_data_i[7];
      mem_438_sv2v_reg <= w_data_i[6];
      mem_437_sv2v_reg <= w_data_i[5];
      mem_436_sv2v_reg <= w_data_i[4];
      mem_435_sv2v_reg <= w_data_i[3];
      mem_434_sv2v_reg <= w_data_i[2];
      mem_433_sv2v_reg <= w_data_i[1];
      mem_432_sv2v_reg <= w_data_i[0];
    end 
    if(N167) begin
      mem_431_sv2v_reg <= w_data_i[15];
      mem_430_sv2v_reg <= w_data_i[14];
      mem_429_sv2v_reg <= w_data_i[13];
      mem_428_sv2v_reg <= w_data_i[12];
      mem_427_sv2v_reg <= w_data_i[11];
      mem_426_sv2v_reg <= w_data_i[10];
      mem_425_sv2v_reg <= w_data_i[9];
      mem_424_sv2v_reg <= w_data_i[8];
      mem_423_sv2v_reg <= w_data_i[7];
      mem_422_sv2v_reg <= w_data_i[6];
      mem_421_sv2v_reg <= w_data_i[5];
      mem_420_sv2v_reg <= w_data_i[4];
      mem_419_sv2v_reg <= w_data_i[3];
      mem_418_sv2v_reg <= w_data_i[2];
      mem_417_sv2v_reg <= w_data_i[1];
      mem_416_sv2v_reg <= w_data_i[0];
    end 
    if(N166) begin
      mem_415_sv2v_reg <= w_data_i[15];
      mem_414_sv2v_reg <= w_data_i[14];
      mem_413_sv2v_reg <= w_data_i[13];
      mem_412_sv2v_reg <= w_data_i[12];
      mem_411_sv2v_reg <= w_data_i[11];
      mem_410_sv2v_reg <= w_data_i[10];
      mem_409_sv2v_reg <= w_data_i[9];
      mem_408_sv2v_reg <= w_data_i[8];
      mem_407_sv2v_reg <= w_data_i[7];
      mem_406_sv2v_reg <= w_data_i[6];
      mem_405_sv2v_reg <= w_data_i[5];
      mem_404_sv2v_reg <= w_data_i[4];
      mem_403_sv2v_reg <= w_data_i[3];
      mem_402_sv2v_reg <= w_data_i[2];
      mem_401_sv2v_reg <= w_data_i[1];
      mem_400_sv2v_reg <= w_data_i[0];
    end 
    if(N165) begin
      mem_399_sv2v_reg <= w_data_i[15];
      mem_398_sv2v_reg <= w_data_i[14];
      mem_397_sv2v_reg <= w_data_i[13];
      mem_396_sv2v_reg <= w_data_i[12];
      mem_395_sv2v_reg <= w_data_i[11];
      mem_394_sv2v_reg <= w_data_i[10];
      mem_393_sv2v_reg <= w_data_i[9];
      mem_392_sv2v_reg <= w_data_i[8];
      mem_391_sv2v_reg <= w_data_i[7];
      mem_390_sv2v_reg <= w_data_i[6];
      mem_389_sv2v_reg <= w_data_i[5];
      mem_388_sv2v_reg <= w_data_i[4];
      mem_387_sv2v_reg <= w_data_i[3];
      mem_386_sv2v_reg <= w_data_i[2];
      mem_385_sv2v_reg <= w_data_i[1];
      mem_384_sv2v_reg <= w_data_i[0];
    end 
    if(N164) begin
      mem_383_sv2v_reg <= w_data_i[15];
      mem_382_sv2v_reg <= w_data_i[14];
      mem_381_sv2v_reg <= w_data_i[13];
      mem_380_sv2v_reg <= w_data_i[12];
      mem_379_sv2v_reg <= w_data_i[11];
      mem_378_sv2v_reg <= w_data_i[10];
      mem_377_sv2v_reg <= w_data_i[9];
      mem_376_sv2v_reg <= w_data_i[8];
      mem_375_sv2v_reg <= w_data_i[7];
      mem_374_sv2v_reg <= w_data_i[6];
      mem_373_sv2v_reg <= w_data_i[5];
      mem_372_sv2v_reg <= w_data_i[4];
      mem_371_sv2v_reg <= w_data_i[3];
      mem_370_sv2v_reg <= w_data_i[2];
      mem_369_sv2v_reg <= w_data_i[1];
      mem_368_sv2v_reg <= w_data_i[0];
    end 
    if(N163) begin
      mem_367_sv2v_reg <= w_data_i[15];
      mem_366_sv2v_reg <= w_data_i[14];
      mem_365_sv2v_reg <= w_data_i[13];
      mem_364_sv2v_reg <= w_data_i[12];
      mem_363_sv2v_reg <= w_data_i[11];
      mem_362_sv2v_reg <= w_data_i[10];
      mem_361_sv2v_reg <= w_data_i[9];
      mem_360_sv2v_reg <= w_data_i[8];
      mem_359_sv2v_reg <= w_data_i[7];
      mem_358_sv2v_reg <= w_data_i[6];
      mem_357_sv2v_reg <= w_data_i[5];
      mem_356_sv2v_reg <= w_data_i[4];
      mem_355_sv2v_reg <= w_data_i[3];
      mem_354_sv2v_reg <= w_data_i[2];
      mem_353_sv2v_reg <= w_data_i[1];
      mem_352_sv2v_reg <= w_data_i[0];
    end 
    if(N162) begin
      mem_351_sv2v_reg <= w_data_i[15];
      mem_350_sv2v_reg <= w_data_i[14];
      mem_349_sv2v_reg <= w_data_i[13];
      mem_348_sv2v_reg <= w_data_i[12];
      mem_347_sv2v_reg <= w_data_i[11];
      mem_346_sv2v_reg <= w_data_i[10];
      mem_345_sv2v_reg <= w_data_i[9];
      mem_344_sv2v_reg <= w_data_i[8];
      mem_343_sv2v_reg <= w_data_i[7];
      mem_342_sv2v_reg <= w_data_i[6];
      mem_341_sv2v_reg <= w_data_i[5];
      mem_340_sv2v_reg <= w_data_i[4];
      mem_339_sv2v_reg <= w_data_i[3];
      mem_338_sv2v_reg <= w_data_i[2];
      mem_337_sv2v_reg <= w_data_i[1];
      mem_336_sv2v_reg <= w_data_i[0];
    end 
    if(N161) begin
      mem_335_sv2v_reg <= w_data_i[15];
      mem_334_sv2v_reg <= w_data_i[14];
      mem_333_sv2v_reg <= w_data_i[13];
      mem_332_sv2v_reg <= w_data_i[12];
      mem_331_sv2v_reg <= w_data_i[11];
      mem_330_sv2v_reg <= w_data_i[10];
      mem_329_sv2v_reg <= w_data_i[9];
      mem_328_sv2v_reg <= w_data_i[8];
      mem_327_sv2v_reg <= w_data_i[7];
      mem_326_sv2v_reg <= w_data_i[6];
      mem_325_sv2v_reg <= w_data_i[5];
      mem_324_sv2v_reg <= w_data_i[4];
      mem_323_sv2v_reg <= w_data_i[3];
      mem_322_sv2v_reg <= w_data_i[2];
      mem_321_sv2v_reg <= w_data_i[1];
      mem_320_sv2v_reg <= w_data_i[0];
    end 
    if(N160) begin
      mem_319_sv2v_reg <= w_data_i[15];
      mem_318_sv2v_reg <= w_data_i[14];
      mem_317_sv2v_reg <= w_data_i[13];
      mem_316_sv2v_reg <= w_data_i[12];
      mem_315_sv2v_reg <= w_data_i[11];
      mem_314_sv2v_reg <= w_data_i[10];
      mem_313_sv2v_reg <= w_data_i[9];
      mem_312_sv2v_reg <= w_data_i[8];
      mem_311_sv2v_reg <= w_data_i[7];
      mem_310_sv2v_reg <= w_data_i[6];
      mem_309_sv2v_reg <= w_data_i[5];
      mem_308_sv2v_reg <= w_data_i[4];
      mem_307_sv2v_reg <= w_data_i[3];
      mem_306_sv2v_reg <= w_data_i[2];
      mem_305_sv2v_reg <= w_data_i[1];
      mem_304_sv2v_reg <= w_data_i[0];
    end 
    if(N159) begin
      mem_303_sv2v_reg <= w_data_i[15];
      mem_302_sv2v_reg <= w_data_i[14];
      mem_301_sv2v_reg <= w_data_i[13];
      mem_300_sv2v_reg <= w_data_i[12];
      mem_299_sv2v_reg <= w_data_i[11];
      mem_298_sv2v_reg <= w_data_i[10];
      mem_297_sv2v_reg <= w_data_i[9];
      mem_296_sv2v_reg <= w_data_i[8];
      mem_295_sv2v_reg <= w_data_i[7];
      mem_294_sv2v_reg <= w_data_i[6];
      mem_293_sv2v_reg <= w_data_i[5];
      mem_292_sv2v_reg <= w_data_i[4];
      mem_291_sv2v_reg <= w_data_i[3];
      mem_290_sv2v_reg <= w_data_i[2];
      mem_289_sv2v_reg <= w_data_i[1];
      mem_288_sv2v_reg <= w_data_i[0];
    end 
    if(N158) begin
      mem_287_sv2v_reg <= w_data_i[15];
      mem_286_sv2v_reg <= w_data_i[14];
      mem_285_sv2v_reg <= w_data_i[13];
      mem_284_sv2v_reg <= w_data_i[12];
      mem_283_sv2v_reg <= w_data_i[11];
      mem_282_sv2v_reg <= w_data_i[10];
      mem_281_sv2v_reg <= w_data_i[9];
      mem_280_sv2v_reg <= w_data_i[8];
      mem_279_sv2v_reg <= w_data_i[7];
      mem_278_sv2v_reg <= w_data_i[6];
      mem_277_sv2v_reg <= w_data_i[5];
      mem_276_sv2v_reg <= w_data_i[4];
      mem_275_sv2v_reg <= w_data_i[3];
      mem_274_sv2v_reg <= w_data_i[2];
      mem_273_sv2v_reg <= w_data_i[1];
      mem_272_sv2v_reg <= w_data_i[0];
    end 
    if(N157) begin
      mem_271_sv2v_reg <= w_data_i[15];
      mem_270_sv2v_reg <= w_data_i[14];
      mem_269_sv2v_reg <= w_data_i[13];
      mem_268_sv2v_reg <= w_data_i[12];
      mem_267_sv2v_reg <= w_data_i[11];
      mem_266_sv2v_reg <= w_data_i[10];
      mem_265_sv2v_reg <= w_data_i[9];
      mem_264_sv2v_reg <= w_data_i[8];
      mem_263_sv2v_reg <= w_data_i[7];
      mem_262_sv2v_reg <= w_data_i[6];
      mem_261_sv2v_reg <= w_data_i[5];
      mem_260_sv2v_reg <= w_data_i[4];
      mem_259_sv2v_reg <= w_data_i[3];
      mem_258_sv2v_reg <= w_data_i[2];
      mem_257_sv2v_reg <= w_data_i[1];
      mem_256_sv2v_reg <= w_data_i[0];
    end 
    if(N156) begin
      mem_255_sv2v_reg <= w_data_i[15];
      mem_254_sv2v_reg <= w_data_i[14];
      mem_253_sv2v_reg <= w_data_i[13];
      mem_252_sv2v_reg <= w_data_i[12];
      mem_251_sv2v_reg <= w_data_i[11];
      mem_250_sv2v_reg <= w_data_i[10];
      mem_249_sv2v_reg <= w_data_i[9];
      mem_248_sv2v_reg <= w_data_i[8];
      mem_247_sv2v_reg <= w_data_i[7];
      mem_246_sv2v_reg <= w_data_i[6];
      mem_245_sv2v_reg <= w_data_i[5];
      mem_244_sv2v_reg <= w_data_i[4];
      mem_243_sv2v_reg <= w_data_i[3];
      mem_242_sv2v_reg <= w_data_i[2];
      mem_241_sv2v_reg <= w_data_i[1];
      mem_240_sv2v_reg <= w_data_i[0];
    end 
    if(N155) begin
      mem_239_sv2v_reg <= w_data_i[15];
      mem_238_sv2v_reg <= w_data_i[14];
      mem_237_sv2v_reg <= w_data_i[13];
      mem_236_sv2v_reg <= w_data_i[12];
      mem_235_sv2v_reg <= w_data_i[11];
      mem_234_sv2v_reg <= w_data_i[10];
      mem_233_sv2v_reg <= w_data_i[9];
      mem_232_sv2v_reg <= w_data_i[8];
      mem_231_sv2v_reg <= w_data_i[7];
      mem_230_sv2v_reg <= w_data_i[6];
      mem_229_sv2v_reg <= w_data_i[5];
      mem_228_sv2v_reg <= w_data_i[4];
      mem_227_sv2v_reg <= w_data_i[3];
      mem_226_sv2v_reg <= w_data_i[2];
      mem_225_sv2v_reg <= w_data_i[1];
      mem_224_sv2v_reg <= w_data_i[0];
    end 
    if(N154) begin
      mem_223_sv2v_reg <= w_data_i[15];
      mem_222_sv2v_reg <= w_data_i[14];
      mem_221_sv2v_reg <= w_data_i[13];
      mem_220_sv2v_reg <= w_data_i[12];
      mem_219_sv2v_reg <= w_data_i[11];
      mem_218_sv2v_reg <= w_data_i[10];
      mem_217_sv2v_reg <= w_data_i[9];
      mem_216_sv2v_reg <= w_data_i[8];
      mem_215_sv2v_reg <= w_data_i[7];
      mem_214_sv2v_reg <= w_data_i[6];
      mem_213_sv2v_reg <= w_data_i[5];
      mem_212_sv2v_reg <= w_data_i[4];
      mem_211_sv2v_reg <= w_data_i[3];
      mem_210_sv2v_reg <= w_data_i[2];
      mem_209_sv2v_reg <= w_data_i[1];
      mem_208_sv2v_reg <= w_data_i[0];
    end 
    if(N153) begin
      mem_207_sv2v_reg <= w_data_i[15];
      mem_206_sv2v_reg <= w_data_i[14];
      mem_205_sv2v_reg <= w_data_i[13];
      mem_204_sv2v_reg <= w_data_i[12];
      mem_203_sv2v_reg <= w_data_i[11];
      mem_202_sv2v_reg <= w_data_i[10];
      mem_201_sv2v_reg <= w_data_i[9];
      mem_200_sv2v_reg <= w_data_i[8];
      mem_199_sv2v_reg <= w_data_i[7];
      mem_198_sv2v_reg <= w_data_i[6];
      mem_197_sv2v_reg <= w_data_i[5];
      mem_196_sv2v_reg <= w_data_i[4];
      mem_195_sv2v_reg <= w_data_i[3];
      mem_194_sv2v_reg <= w_data_i[2];
      mem_193_sv2v_reg <= w_data_i[1];
      mem_192_sv2v_reg <= w_data_i[0];
    end 
    if(N152) begin
      mem_191_sv2v_reg <= w_data_i[15];
      mem_190_sv2v_reg <= w_data_i[14];
      mem_189_sv2v_reg <= w_data_i[13];
      mem_188_sv2v_reg <= w_data_i[12];
      mem_187_sv2v_reg <= w_data_i[11];
      mem_186_sv2v_reg <= w_data_i[10];
      mem_185_sv2v_reg <= w_data_i[9];
      mem_184_sv2v_reg <= w_data_i[8];
      mem_183_sv2v_reg <= w_data_i[7];
      mem_182_sv2v_reg <= w_data_i[6];
      mem_181_sv2v_reg <= w_data_i[5];
      mem_180_sv2v_reg <= w_data_i[4];
      mem_179_sv2v_reg <= w_data_i[3];
      mem_178_sv2v_reg <= w_data_i[2];
      mem_177_sv2v_reg <= w_data_i[1];
      mem_176_sv2v_reg <= w_data_i[0];
    end 
    if(N151) begin
      mem_175_sv2v_reg <= w_data_i[15];
      mem_174_sv2v_reg <= w_data_i[14];
      mem_173_sv2v_reg <= w_data_i[13];
      mem_172_sv2v_reg <= w_data_i[12];
      mem_171_sv2v_reg <= w_data_i[11];
      mem_170_sv2v_reg <= w_data_i[10];
      mem_169_sv2v_reg <= w_data_i[9];
      mem_168_sv2v_reg <= w_data_i[8];
      mem_167_sv2v_reg <= w_data_i[7];
      mem_166_sv2v_reg <= w_data_i[6];
      mem_165_sv2v_reg <= w_data_i[5];
      mem_164_sv2v_reg <= w_data_i[4];
      mem_163_sv2v_reg <= w_data_i[3];
      mem_162_sv2v_reg <= w_data_i[2];
      mem_161_sv2v_reg <= w_data_i[1];
      mem_160_sv2v_reg <= w_data_i[0];
    end 
    if(N150) begin
      mem_159_sv2v_reg <= w_data_i[15];
      mem_158_sv2v_reg <= w_data_i[14];
      mem_157_sv2v_reg <= w_data_i[13];
      mem_156_sv2v_reg <= w_data_i[12];
      mem_155_sv2v_reg <= w_data_i[11];
      mem_154_sv2v_reg <= w_data_i[10];
      mem_153_sv2v_reg <= w_data_i[9];
      mem_152_sv2v_reg <= w_data_i[8];
      mem_151_sv2v_reg <= w_data_i[7];
      mem_150_sv2v_reg <= w_data_i[6];
      mem_149_sv2v_reg <= w_data_i[5];
      mem_148_sv2v_reg <= w_data_i[4];
      mem_147_sv2v_reg <= w_data_i[3];
      mem_146_sv2v_reg <= w_data_i[2];
      mem_145_sv2v_reg <= w_data_i[1];
      mem_144_sv2v_reg <= w_data_i[0];
    end 
    if(N149) begin
      mem_143_sv2v_reg <= w_data_i[15];
      mem_142_sv2v_reg <= w_data_i[14];
      mem_141_sv2v_reg <= w_data_i[13];
      mem_140_sv2v_reg <= w_data_i[12];
      mem_139_sv2v_reg <= w_data_i[11];
      mem_138_sv2v_reg <= w_data_i[10];
      mem_137_sv2v_reg <= w_data_i[9];
      mem_136_sv2v_reg <= w_data_i[8];
      mem_135_sv2v_reg <= w_data_i[7];
      mem_134_sv2v_reg <= w_data_i[6];
      mem_133_sv2v_reg <= w_data_i[5];
      mem_132_sv2v_reg <= w_data_i[4];
      mem_131_sv2v_reg <= w_data_i[3];
      mem_130_sv2v_reg <= w_data_i[2];
      mem_129_sv2v_reg <= w_data_i[1];
      mem_128_sv2v_reg <= w_data_i[0];
    end 
    if(N148) begin
      mem_127_sv2v_reg <= w_data_i[15];
      mem_126_sv2v_reg <= w_data_i[14];
      mem_125_sv2v_reg <= w_data_i[13];
      mem_124_sv2v_reg <= w_data_i[12];
      mem_123_sv2v_reg <= w_data_i[11];
      mem_122_sv2v_reg <= w_data_i[10];
      mem_121_sv2v_reg <= w_data_i[9];
      mem_120_sv2v_reg <= w_data_i[8];
      mem_119_sv2v_reg <= w_data_i[7];
      mem_118_sv2v_reg <= w_data_i[6];
      mem_117_sv2v_reg <= w_data_i[5];
      mem_116_sv2v_reg <= w_data_i[4];
      mem_115_sv2v_reg <= w_data_i[3];
      mem_114_sv2v_reg <= w_data_i[2];
      mem_113_sv2v_reg <= w_data_i[1];
      mem_112_sv2v_reg <= w_data_i[0];
    end 
    if(N147) begin
      mem_111_sv2v_reg <= w_data_i[15];
      mem_110_sv2v_reg <= w_data_i[14];
      mem_109_sv2v_reg <= w_data_i[13];
      mem_108_sv2v_reg <= w_data_i[12];
      mem_107_sv2v_reg <= w_data_i[11];
      mem_106_sv2v_reg <= w_data_i[10];
      mem_105_sv2v_reg <= w_data_i[9];
      mem_104_sv2v_reg <= w_data_i[8];
      mem_103_sv2v_reg <= w_data_i[7];
      mem_102_sv2v_reg <= w_data_i[6];
      mem_101_sv2v_reg <= w_data_i[5];
      mem_100_sv2v_reg <= w_data_i[4];
      mem_99_sv2v_reg <= w_data_i[3];
      mem_98_sv2v_reg <= w_data_i[2];
      mem_97_sv2v_reg <= w_data_i[1];
      mem_96_sv2v_reg <= w_data_i[0];
    end 
    if(N146) begin
      mem_95_sv2v_reg <= w_data_i[15];
      mem_94_sv2v_reg <= w_data_i[14];
      mem_93_sv2v_reg <= w_data_i[13];
      mem_92_sv2v_reg <= w_data_i[12];
      mem_91_sv2v_reg <= w_data_i[11];
      mem_90_sv2v_reg <= w_data_i[10];
      mem_89_sv2v_reg <= w_data_i[9];
      mem_88_sv2v_reg <= w_data_i[8];
      mem_87_sv2v_reg <= w_data_i[7];
      mem_86_sv2v_reg <= w_data_i[6];
      mem_85_sv2v_reg <= w_data_i[5];
      mem_84_sv2v_reg <= w_data_i[4];
      mem_83_sv2v_reg <= w_data_i[3];
      mem_82_sv2v_reg <= w_data_i[2];
      mem_81_sv2v_reg <= w_data_i[1];
      mem_80_sv2v_reg <= w_data_i[0];
    end 
    if(N145) begin
      mem_79_sv2v_reg <= w_data_i[15];
      mem_78_sv2v_reg <= w_data_i[14];
      mem_77_sv2v_reg <= w_data_i[13];
      mem_76_sv2v_reg <= w_data_i[12];
      mem_75_sv2v_reg <= w_data_i[11];
      mem_74_sv2v_reg <= w_data_i[10];
      mem_73_sv2v_reg <= w_data_i[9];
      mem_72_sv2v_reg <= w_data_i[8];
      mem_71_sv2v_reg <= w_data_i[7];
      mem_70_sv2v_reg <= w_data_i[6];
      mem_69_sv2v_reg <= w_data_i[5];
      mem_68_sv2v_reg <= w_data_i[4];
      mem_67_sv2v_reg <= w_data_i[3];
      mem_66_sv2v_reg <= w_data_i[2];
      mem_65_sv2v_reg <= w_data_i[1];
      mem_64_sv2v_reg <= w_data_i[0];
    end 
    if(N144) begin
      mem_63_sv2v_reg <= w_data_i[15];
      mem_62_sv2v_reg <= w_data_i[14];
      mem_61_sv2v_reg <= w_data_i[13];
      mem_60_sv2v_reg <= w_data_i[12];
      mem_59_sv2v_reg <= w_data_i[11];
      mem_58_sv2v_reg <= w_data_i[10];
      mem_57_sv2v_reg <= w_data_i[9];
      mem_56_sv2v_reg <= w_data_i[8];
      mem_55_sv2v_reg <= w_data_i[7];
      mem_54_sv2v_reg <= w_data_i[6];
      mem_53_sv2v_reg <= w_data_i[5];
      mem_52_sv2v_reg <= w_data_i[4];
      mem_51_sv2v_reg <= w_data_i[3];
      mem_50_sv2v_reg <= w_data_i[2];
      mem_49_sv2v_reg <= w_data_i[1];
      mem_48_sv2v_reg <= w_data_i[0];
    end 
    if(N143) begin
      mem_47_sv2v_reg <= w_data_i[15];
      mem_46_sv2v_reg <= w_data_i[14];
      mem_45_sv2v_reg <= w_data_i[13];
      mem_44_sv2v_reg <= w_data_i[12];
      mem_43_sv2v_reg <= w_data_i[11];
      mem_42_sv2v_reg <= w_data_i[10];
      mem_41_sv2v_reg <= w_data_i[9];
      mem_40_sv2v_reg <= w_data_i[8];
      mem_39_sv2v_reg <= w_data_i[7];
      mem_38_sv2v_reg <= w_data_i[6];
      mem_37_sv2v_reg <= w_data_i[5];
      mem_36_sv2v_reg <= w_data_i[4];
      mem_35_sv2v_reg <= w_data_i[3];
      mem_34_sv2v_reg <= w_data_i[2];
      mem_33_sv2v_reg <= w_data_i[1];
      mem_32_sv2v_reg <= w_data_i[0];
    end 
    if(N142) begin
      mem_31_sv2v_reg <= w_data_i[15];
      mem_30_sv2v_reg <= w_data_i[14];
      mem_29_sv2v_reg <= w_data_i[13];
      mem_28_sv2v_reg <= w_data_i[12];
      mem_27_sv2v_reg <= w_data_i[11];
      mem_26_sv2v_reg <= w_data_i[10];
      mem_25_sv2v_reg <= w_data_i[9];
      mem_24_sv2v_reg <= w_data_i[8];
      mem_23_sv2v_reg <= w_data_i[7];
      mem_22_sv2v_reg <= w_data_i[6];
      mem_21_sv2v_reg <= w_data_i[5];
      mem_20_sv2v_reg <= w_data_i[4];
      mem_19_sv2v_reg <= w_data_i[3];
      mem_18_sv2v_reg <= w_data_i[2];
      mem_17_sv2v_reg <= w_data_i[1];
      mem_16_sv2v_reg <= w_data_i[0];
    end 
    if(N141) begin
      mem_15_sv2v_reg <= w_data_i[15];
      mem_14_sv2v_reg <= w_data_i[14];
      mem_13_sv2v_reg <= w_data_i[13];
      mem_12_sv2v_reg <= w_data_i[12];
      mem_11_sv2v_reg <= w_data_i[11];
      mem_10_sv2v_reg <= w_data_i[10];
      mem_9_sv2v_reg <= w_data_i[9];
      mem_8_sv2v_reg <= w_data_i[8];
      mem_7_sv2v_reg <= w_data_i[7];
      mem_6_sv2v_reg <= w_data_i[6];
      mem_5_sv2v_reg <= w_data_i[5];
      mem_4_sv2v_reg <= w_data_i[4];
      mem_3_sv2v_reg <= w_data_i[3];
      mem_2_sv2v_reg <= w_data_i[2];
      mem_1_sv2v_reg <= w_data_i[1];
      mem_0_sv2v_reg <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p16_els_p64_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [5:0] w_addr_i;
  input [15:0] w_data_i;
  input [5:0] r_addr_i;
  output [15:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [15:0] r_data_o;

  bsg_mem_1r1w_synth_width_p16_els_p64_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_launch_sync_sync_posedge_7_unit
(
  iclk_i,
  iclk_reset_i,
  oclk_i,
  iclk_data_i,
  iclk_data_o,
  oclk_data_o
);

  input [6:0] iclk_data_i;
  output [6:0] iclk_data_o;
  output [6:0] oclk_data_o;
  input iclk_i;
  input iclk_reset_i;
  input oclk_i;
  wire [6:0] iclk_data_o,oclk_data_o,bsg_SYNC_1_r;
  reg iclk_data_o_6_sv2v_reg,iclk_data_o_5_sv2v_reg,iclk_data_o_4_sv2v_reg,
  iclk_data_o_3_sv2v_reg,iclk_data_o_2_sv2v_reg,iclk_data_o_1_sv2v_reg,
  iclk_data_o_0_sv2v_reg,bsg_SYNC_1_r_6_sv2v_reg,bsg_SYNC_1_r_5_sv2v_reg,bsg_SYNC_1_r_4_sv2v_reg,
  bsg_SYNC_1_r_3_sv2v_reg,bsg_SYNC_1_r_2_sv2v_reg,bsg_SYNC_1_r_1_sv2v_reg,
  bsg_SYNC_1_r_0_sv2v_reg,oclk_data_o_6_sv2v_reg,oclk_data_o_5_sv2v_reg,oclk_data_o_4_sv2v_reg,
  oclk_data_o_3_sv2v_reg,oclk_data_o_2_sv2v_reg,oclk_data_o_1_sv2v_reg,
  oclk_data_o_0_sv2v_reg;
  assign iclk_data_o[6] = iclk_data_o_6_sv2v_reg;
  assign iclk_data_o[5] = iclk_data_o_5_sv2v_reg;
  assign iclk_data_o[4] = iclk_data_o_4_sv2v_reg;
  assign iclk_data_o[3] = iclk_data_o_3_sv2v_reg;
  assign iclk_data_o[2] = iclk_data_o_2_sv2v_reg;
  assign iclk_data_o[1] = iclk_data_o_1_sv2v_reg;
  assign iclk_data_o[0] = iclk_data_o_0_sv2v_reg;
  assign bsg_SYNC_1_r[6] = bsg_SYNC_1_r_6_sv2v_reg;
  assign bsg_SYNC_1_r[5] = bsg_SYNC_1_r_5_sv2v_reg;
  assign bsg_SYNC_1_r[4] = bsg_SYNC_1_r_4_sv2v_reg;
  assign bsg_SYNC_1_r[3] = bsg_SYNC_1_r_3_sv2v_reg;
  assign bsg_SYNC_1_r[2] = bsg_SYNC_1_r_2_sv2v_reg;
  assign bsg_SYNC_1_r[1] = bsg_SYNC_1_r_1_sv2v_reg;
  assign bsg_SYNC_1_r[0] = bsg_SYNC_1_r_0_sv2v_reg;
  assign oclk_data_o[6] = oclk_data_o_6_sv2v_reg;
  assign oclk_data_o[5] = oclk_data_o_5_sv2v_reg;
  assign oclk_data_o[4] = oclk_data_o_4_sv2v_reg;
  assign oclk_data_o[3] = oclk_data_o_3_sv2v_reg;
  assign oclk_data_o[2] = oclk_data_o_2_sv2v_reg;
  assign oclk_data_o[1] = oclk_data_o_1_sv2v_reg;
  assign oclk_data_o[0] = oclk_data_o_0_sv2v_reg;

  always @(posedge iclk_i) begin
    if(iclk_reset_i) begin
      iclk_data_o_6_sv2v_reg <= 1'b0;
      iclk_data_o_5_sv2v_reg <= 1'b0;
      iclk_data_o_4_sv2v_reg <= 1'b0;
      iclk_data_o_3_sv2v_reg <= 1'b0;
      iclk_data_o_2_sv2v_reg <= 1'b0;
      iclk_data_o_1_sv2v_reg <= 1'b0;
      iclk_data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      iclk_data_o_6_sv2v_reg <= iclk_data_i[6];
      iclk_data_o_5_sv2v_reg <= iclk_data_i[5];
      iclk_data_o_4_sv2v_reg <= iclk_data_i[4];
      iclk_data_o_3_sv2v_reg <= iclk_data_i[3];
      iclk_data_o_2_sv2v_reg <= iclk_data_i[2];
      iclk_data_o_1_sv2v_reg <= iclk_data_i[1];
      iclk_data_o_0_sv2v_reg <= iclk_data_i[0];
    end 
  end


  always @(posedge oclk_i) begin
    if(1'b1) begin
      bsg_SYNC_1_r_6_sv2v_reg <= iclk_data_o[6];
      bsg_SYNC_1_r_5_sv2v_reg <= iclk_data_o[5];
      bsg_SYNC_1_r_4_sv2v_reg <= iclk_data_o[4];
      bsg_SYNC_1_r_3_sv2v_reg <= iclk_data_o[3];
      bsg_SYNC_1_r_2_sv2v_reg <= iclk_data_o[2];
      bsg_SYNC_1_r_1_sv2v_reg <= iclk_data_o[1];
      bsg_SYNC_1_r_0_sv2v_reg <= iclk_data_o[0];
      oclk_data_o_6_sv2v_reg <= bsg_SYNC_1_r[6];
      oclk_data_o_5_sv2v_reg <= bsg_SYNC_1_r[5];
      oclk_data_o_4_sv2v_reg <= bsg_SYNC_1_r[4];
      oclk_data_o_3_sv2v_reg <= bsg_SYNC_1_r[3];
      oclk_data_o_2_sv2v_reg <= bsg_SYNC_1_r[2];
      oclk_data_o_1_sv2v_reg <= bsg_SYNC_1_r[1];
      oclk_data_o_0_sv2v_reg <= bsg_SYNC_1_r[0];
    end 
  end


endmodule



module bsg_launch_sync_sync_width_p7_use_negedge_for_launch_p0_use_async_reset_p0
(
  iclk_i,
  iclk_reset_i,
  oclk_i,
  iclk_data_i,
  iclk_data_o,
  oclk_data_o
);

  input [6:0] iclk_data_i;
  output [6:0] iclk_data_o;
  output [6:0] oclk_data_o;
  input iclk_i;
  input iclk_reset_i;
  input oclk_i;
  wire [6:0] iclk_data_o,oclk_data_o;

  bsg_launch_sync_sync_posedge_7_unit
  sync_p_z_blss 
  (
    .iclk_i(iclk_i),
    .iclk_reset_i(iclk_reset_i),
    .oclk_i(oclk_i),
    .iclk_data_i(iclk_data_i),
    .iclk_data_o(iclk_data_o),
    .oclk_data_o(oclk_data_o)
  );


endmodule



module bsg_async_ptr_gray_lg_size_p7
(
  w_clk_i,
  w_reset_i,
  w_inc_i,
  r_clk_i,
  w_ptr_binary_r_o,
  w_ptr_gray_r_o,
  w_ptr_gray_r_rsync_o
);

  output [6:0] w_ptr_binary_r_o;
  output [6:0] w_ptr_gray_r_o;
  output [6:0] w_ptr_gray_r_rsync_o;
  input w_clk_i;
  input w_reset_i;
  input w_inc_i;
  input r_clk_i;
  wire [6:0] w_ptr_binary_r_o,w_ptr_gray_r_o,w_ptr_gray_r_rsync_o,w_ptr_p1_r,w_ptr_p2,
  w_ptr_n,w_ptr_p1_n,w_ptr_gray_n;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8;
  reg w_ptr_p1_r_6_sv2v_reg,w_ptr_p1_r_5_sv2v_reg,w_ptr_p1_r_4_sv2v_reg,
  w_ptr_p1_r_3_sv2v_reg,w_ptr_p1_r_2_sv2v_reg,w_ptr_p1_r_1_sv2v_reg,w_ptr_p1_r_0_sv2v_reg,
  w_ptr_binary_r_o_6_sv2v_reg,w_ptr_binary_r_o_5_sv2v_reg,w_ptr_binary_r_o_4_sv2v_reg,
  w_ptr_binary_r_o_3_sv2v_reg,w_ptr_binary_r_o_2_sv2v_reg,
  w_ptr_binary_r_o_1_sv2v_reg,w_ptr_binary_r_o_0_sv2v_reg;
  assign w_ptr_p1_r[6] = w_ptr_p1_r_6_sv2v_reg;
  assign w_ptr_p1_r[5] = w_ptr_p1_r_5_sv2v_reg;
  assign w_ptr_p1_r[4] = w_ptr_p1_r_4_sv2v_reg;
  assign w_ptr_p1_r[3] = w_ptr_p1_r_3_sv2v_reg;
  assign w_ptr_p1_r[2] = w_ptr_p1_r_2_sv2v_reg;
  assign w_ptr_p1_r[1] = w_ptr_p1_r_1_sv2v_reg;
  assign w_ptr_p1_r[0] = w_ptr_p1_r_0_sv2v_reg;
  assign w_ptr_binary_r_o[6] = w_ptr_binary_r_o_6_sv2v_reg;
  assign w_ptr_binary_r_o[5] = w_ptr_binary_r_o_5_sv2v_reg;
  assign w_ptr_binary_r_o[4] = w_ptr_binary_r_o_4_sv2v_reg;
  assign w_ptr_binary_r_o[3] = w_ptr_binary_r_o_3_sv2v_reg;
  assign w_ptr_binary_r_o[2] = w_ptr_binary_r_o_2_sv2v_reg;
  assign w_ptr_binary_r_o[1] = w_ptr_binary_r_o_1_sv2v_reg;
  assign w_ptr_binary_r_o[0] = w_ptr_binary_r_o_0_sv2v_reg;

  bsg_launch_sync_sync_width_p7_use_negedge_for_launch_p0_use_async_reset_p0
  ptr_sync
  (
    .iclk_i(w_clk_i),
    .iclk_reset_i(w_reset_i),
    .oclk_i(r_clk_i),
    .iclk_data_i(w_ptr_gray_n),
    .iclk_data_o(w_ptr_gray_r_o),
    .oclk_data_o(w_ptr_gray_r_rsync_o)
  );

  assign w_ptr_p2 = w_ptr_p1_r + 1'b1;
  assign w_ptr_n = (N0)? w_ptr_p1_r : 
                   (N1)? w_ptr_binary_r_o : 1'b0;
  assign N0 = w_inc_i;
  assign N1 = N2;
  assign w_ptr_p1_n = (N0)? w_ptr_p2 : 
                      (N1)? w_ptr_p1_r : 1'b0;
  assign w_ptr_gray_n = (N0)? { w_ptr_p1_r[6:6], N3, N4, N5, N6, N7, N8 } : 
                        (N1)? w_ptr_gray_r_o : 1'b0;
  assign N2 = ~w_inc_i;
  assign N3 = w_ptr_p1_r[6] ^ w_ptr_p1_r[5];
  assign N4 = w_ptr_p1_r[5] ^ w_ptr_p1_r[4];
  assign N5 = w_ptr_p1_r[4] ^ w_ptr_p1_r[3];
  assign N6 = w_ptr_p1_r[3] ^ w_ptr_p1_r[2];
  assign N7 = w_ptr_p1_r[2] ^ w_ptr_p1_r[1];
  assign N8 = w_ptr_p1_r[1] ^ w_ptr_p1_r[0];

  always @(posedge w_clk_i) begin
    if(w_reset_i) begin
      w_ptr_p1_r_6_sv2v_reg <= 1'b0;
      w_ptr_p1_r_5_sv2v_reg <= 1'b0;
      w_ptr_p1_r_4_sv2v_reg <= 1'b0;
      w_ptr_p1_r_3_sv2v_reg <= 1'b0;
      w_ptr_p1_r_2_sv2v_reg <= 1'b0;
      w_ptr_p1_r_1_sv2v_reg <= 1'b0;
      w_ptr_p1_r_0_sv2v_reg <= 1'b1;
      w_ptr_binary_r_o_6_sv2v_reg <= 1'b0;
      w_ptr_binary_r_o_5_sv2v_reg <= 1'b0;
      w_ptr_binary_r_o_4_sv2v_reg <= 1'b0;
      w_ptr_binary_r_o_3_sv2v_reg <= 1'b0;
      w_ptr_binary_r_o_2_sv2v_reg <= 1'b0;
      w_ptr_binary_r_o_1_sv2v_reg <= 1'b0;
      w_ptr_binary_r_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      w_ptr_p1_r_6_sv2v_reg <= w_ptr_p1_n[6];
      w_ptr_p1_r_5_sv2v_reg <= w_ptr_p1_n[5];
      w_ptr_p1_r_4_sv2v_reg <= w_ptr_p1_n[4];
      w_ptr_p1_r_3_sv2v_reg <= w_ptr_p1_n[3];
      w_ptr_p1_r_2_sv2v_reg <= w_ptr_p1_n[2];
      w_ptr_p1_r_1_sv2v_reg <= w_ptr_p1_n[1];
      w_ptr_p1_r_0_sv2v_reg <= w_ptr_p1_n[0];
      w_ptr_binary_r_o_6_sv2v_reg <= w_ptr_n[6];
      w_ptr_binary_r_o_5_sv2v_reg <= w_ptr_n[5];
      w_ptr_binary_r_o_4_sv2v_reg <= w_ptr_n[4];
      w_ptr_binary_r_o_3_sv2v_reg <= w_ptr_n[3];
      w_ptr_binary_r_o_2_sv2v_reg <= w_ptr_n[2];
      w_ptr_binary_r_o_1_sv2v_reg <= w_ptr_n[1];
      w_ptr_binary_r_o_0_sv2v_reg <= w_ptr_n[0];
    end 
  end


endmodule



module bsg_scan_width_p7_xor_p1
(
  i,
  o
);

  input [6:0] i;
  output [6:0] o;
  wire [6:0] o;
  wire t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__6_,t_1__5_,t_1__4_,
  t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__6_ = i[6] ^ 1'b0;
  assign t_1__5_ = i[5] ^ i[6];
  assign t_1__4_ = i[4] ^ i[5];
  assign t_1__3_ = i[3] ^ i[4];
  assign t_1__2_ = i[2] ^ i[3];
  assign t_1__1_ = i[1] ^ i[2];
  assign t_1__0_ = i[0] ^ i[1];
  assign t_2__6_ = t_1__6_ ^ 1'b0;
  assign t_2__5_ = t_1__5_ ^ 1'b0;
  assign t_2__4_ = t_1__4_ ^ t_1__6_;
  assign t_2__3_ = t_1__3_ ^ t_1__5_;
  assign t_2__2_ = t_1__2_ ^ t_1__4_;
  assign t_2__1_ = t_1__1_ ^ t_1__3_;
  assign t_2__0_ = t_1__0_ ^ t_1__2_;
  assign o[6] = t_2__6_ ^ 1'b0;
  assign o[5] = t_2__5_ ^ 1'b0;
  assign o[4] = t_2__4_ ^ 1'b0;
  assign o[3] = t_2__3_ ^ 1'b0;
  assign o[2] = t_2__2_ ^ t_2__6_;
  assign o[1] = t_2__1_ ^ t_2__5_;
  assign o[0] = t_2__0_ ^ t_2__4_;

endmodule



module bsg_gray_to_binary_width_p7
(
  gray_i,
  binary_o
);

  input [6:0] gray_i;
  output [6:0] binary_o;
  wire [6:0] binary_o;

  bsg_scan_width_p7_xor_p1
  scan_xor
  (
    .i(gray_i),
    .o(binary_o)
  );


endmodule



module bsg_async_fifo_lg_size_p6_width_p16
(
  w_clk_i,
  w_reset_i,
  w_enq_i,
  w_data_i,
  w_full_o,
  r_clk_i,
  r_reset_i,
  r_deq_i,
  r_data_o,
  r_valid_o
);

  input [15:0] w_data_i;
  output [15:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_enq_i;
  input r_clk_i;
  input r_reset_i;
  input r_deq_i;
  output w_full_o;
  output r_valid_o;
  wire [15:0] r_data_o;
  wire w_full_o,r_valid_o,N0,N1;
  wire [6:0] w_ptr_binary_r,r_ptr_binary_r,w_ptr_gray_r,w_ptr_gray_r_rsync,r_ptr_gray_r,
  r_ptr_gray_r_wsync,w_ptr_binary_r_rsync;

  bsg_mem_1r1w_width_p16_els_p64_read_write_same_addr_p0
  MSYNC_1r1w
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_enq_i),
    .w_addr_i(w_ptr_binary_r[5:0]),
    .w_data_i(w_data_i),
    .r_v_i(r_valid_o),
    .r_addr_i(r_ptr_binary_r[5:0]),
    .r_data_o(r_data_o)
  );


  bsg_async_ptr_gray_lg_size_p7
  bapg_wr
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_inc_i(w_enq_i),
    .r_clk_i(r_clk_i),
    .w_ptr_binary_r_o(w_ptr_binary_r),
    .w_ptr_gray_r_o(w_ptr_gray_r),
    .w_ptr_gray_r_rsync_o(w_ptr_gray_r_rsync)
  );


  bsg_async_ptr_gray_lg_size_p7
  bapg_rd
  (
    .w_clk_i(r_clk_i),
    .w_reset_i(r_reset_i),
    .w_inc_i(r_deq_i),
    .r_clk_i(w_clk_i),
    .w_ptr_binary_r_o(r_ptr_binary_r),
    .w_ptr_gray_r_o(r_ptr_gray_r),
    .w_ptr_gray_r_rsync_o(r_ptr_gray_r_wsync)
  );

  assign r_valid_o = r_ptr_gray_r != w_ptr_gray_r_rsync;
  assign w_full_o = w_ptr_gray_r == { N0, N1, r_ptr_gray_r_wsync[4:0] };

  bsg_gray_to_binary_width_p7
  bsg_g2b
  (
    .gray_i(w_ptr_gray_r_rsync),
    .binary_o(w_ptr_binary_r_rsync)
  );

  assign N0 = ~r_ptr_gray_r_wsync[6];
  assign N1 = ~r_ptr_gray_r_wsync[5];

endmodule



module bsg_mem_1r1w_synth_width_p16_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [15:0] w_data_i;
  input [0:0] r_addr_i;
  output [15:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [15:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7;
  wire [31:0] mem;
  reg mem_31_sv2v_reg,mem_30_sv2v_reg,mem_29_sv2v_reg,mem_28_sv2v_reg,mem_27_sv2v_reg,
  mem_26_sv2v_reg,mem_25_sv2v_reg,mem_24_sv2v_reg,mem_23_sv2v_reg,mem_22_sv2v_reg,
  mem_21_sv2v_reg,mem_20_sv2v_reg,mem_19_sv2v_reg,mem_18_sv2v_reg,mem_17_sv2v_reg,
  mem_16_sv2v_reg,mem_15_sv2v_reg,mem_14_sv2v_reg,mem_13_sv2v_reg,mem_12_sv2v_reg,
  mem_11_sv2v_reg,mem_10_sv2v_reg,mem_9_sv2v_reg,mem_8_sv2v_reg,mem_7_sv2v_reg,
  mem_6_sv2v_reg,mem_5_sv2v_reg,mem_4_sv2v_reg,mem_3_sv2v_reg,mem_2_sv2v_reg,
  mem_1_sv2v_reg,mem_0_sv2v_reg;
  assign mem[31] = mem_31_sv2v_reg;
  assign mem[30] = mem_30_sv2v_reg;
  assign mem[29] = mem_29_sv2v_reg;
  assign mem[28] = mem_28_sv2v_reg;
  assign mem[27] = mem_27_sv2v_reg;
  assign mem[26] = mem_26_sv2v_reg;
  assign mem[25] = mem_25_sv2v_reg;
  assign mem[24] = mem_24_sv2v_reg;
  assign mem[23] = mem_23_sv2v_reg;
  assign mem[22] = mem_22_sv2v_reg;
  assign mem[21] = mem_21_sv2v_reg;
  assign mem[20] = mem_20_sv2v_reg;
  assign mem[19] = mem_19_sv2v_reg;
  assign mem[18] = mem_18_sv2v_reg;
  assign mem[17] = mem_17_sv2v_reg;
  assign mem[16] = mem_16_sv2v_reg;
  assign mem[15] = mem_15_sv2v_reg;
  assign mem[14] = mem_14_sv2v_reg;
  assign mem[13] = mem_13_sv2v_reg;
  assign mem[12] = mem_12_sv2v_reg;
  assign mem[11] = mem_11_sv2v_reg;
  assign mem[10] = mem_10_sv2v_reg;
  assign mem[9] = mem_9_sv2v_reg;
  assign mem[8] = mem_8_sv2v_reg;
  assign mem[7] = mem_7_sv2v_reg;
  assign mem[6] = mem_6_sv2v_reg;
  assign mem[5] = mem_5_sv2v_reg;
  assign mem[4] = mem_4_sv2v_reg;
  assign mem[3] = mem_3_sv2v_reg;
  assign mem[2] = mem_2_sv2v_reg;
  assign mem[1] = mem_1_sv2v_reg;
  assign mem[0] = mem_0_sv2v_reg;
  assign r_data_o[15] = (N3)? mem[15] : 
                        (N0)? mem[31] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[14] = (N3)? mem[14] : 
                        (N0)? mem[30] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] : 
                        (N0)? mem[29] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] : 
                        (N0)? mem[28] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] : 
                        (N0)? mem[27] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] : 
                        (N0)? mem[26] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] : 
                       (N0)? mem[25] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] : 
                       (N0)? mem[24] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] : 
                       (N0)? mem[23] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] : 
                       (N0)? mem[22] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[21] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[20] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[19] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[18] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[17] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[16] : 1'b0;
  assign N7 = ~w_addr_i[0];
  assign { N6, N5 } = (N1)? { w_addr_i[0:0], N7 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N6) begin
      mem_31_sv2v_reg <= w_data_i[15];
      mem_30_sv2v_reg <= w_data_i[14];
      mem_29_sv2v_reg <= w_data_i[13];
      mem_28_sv2v_reg <= w_data_i[12];
      mem_27_sv2v_reg <= w_data_i[11];
      mem_26_sv2v_reg <= w_data_i[10];
      mem_25_sv2v_reg <= w_data_i[9];
      mem_24_sv2v_reg <= w_data_i[8];
      mem_23_sv2v_reg <= w_data_i[7];
      mem_22_sv2v_reg <= w_data_i[6];
      mem_21_sv2v_reg <= w_data_i[5];
      mem_20_sv2v_reg <= w_data_i[4];
      mem_19_sv2v_reg <= w_data_i[3];
      mem_18_sv2v_reg <= w_data_i[2];
      mem_17_sv2v_reg <= w_data_i[1];
      mem_16_sv2v_reg <= w_data_i[0];
    end 
    if(N5) begin
      mem_15_sv2v_reg <= w_data_i[15];
      mem_14_sv2v_reg <= w_data_i[14];
      mem_13_sv2v_reg <= w_data_i[13];
      mem_12_sv2v_reg <= w_data_i[12];
      mem_11_sv2v_reg <= w_data_i[11];
      mem_10_sv2v_reg <= w_data_i[10];
      mem_9_sv2v_reg <= w_data_i[9];
      mem_8_sv2v_reg <= w_data_i[8];
      mem_7_sv2v_reg <= w_data_i[7];
      mem_6_sv2v_reg <= w_data_i[6];
      mem_5_sv2v_reg <= w_data_i[5];
      mem_4_sv2v_reg <= w_data_i[4];
      mem_3_sv2v_reg <= w_data_i[3];
      mem_2_sv2v_reg <= w_data_i[2];
      mem_1_sv2v_reg <= w_data_i[1];
      mem_0_sv2v_reg <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p16_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [15:0] w_data_i;
  input [0:0] r_addr_i;
  output [15:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [15:0] r_data_o;

  bsg_mem_1r1w_synth_width_p16_els_p2_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p16
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [15:0] data_i;
  output [15:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [15:0] data_o;
  wire ready_o,v_o,enq_i,tail_r,_0_net_,head_r,empty_r,full_r,N0,N1,N2,N3,N4,N5,N6,N7,
  N8,N9,N10,N11,N12,N13,N14;
  reg full_r_sv2v_reg,tail_r_sv2v_reg,head_r_sv2v_reg,empty_r_sv2v_reg;
  assign full_r = full_r_sv2v_reg;
  assign tail_r = tail_r_sv2v_reg;
  assign head_r = head_r_sv2v_reg;
  assign empty_r = empty_r_sv2v_reg;

  bsg_mem_1r1w_width_p16_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign _0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N5;
  assign N5 = ~full_r;
  assign N1 = enq_i;
  assign N0 = ~tail_r;
  assign N2 = ~head_r;
  assign N3 = N7 | N9;
  assign N7 = empty_r & N6;
  assign N6 = ~enq_i;
  assign N9 = N8 & N6;
  assign N8 = N5 & yumi_i;
  assign N4 = N13 | N14;
  assign N13 = N11 & N12;
  assign N11 = N10 & enq_i;
  assign N10 = ~empty_r;
  assign N12 = ~yumi_i;
  assign N14 = full_r & N12;

  always @(posedge clk_i) begin
    if(reset_i) begin
      full_r_sv2v_reg <= 1'b0;
      empty_r_sv2v_reg <= 1'b1;
    end else if(1'b1) begin
      full_r_sv2v_reg <= N4;
      empty_r_sv2v_reg <= N3;
    end 
    if(reset_i) begin
      tail_r_sv2v_reg <= 1'b0;
    end else if(N1) begin
      tail_r_sv2v_reg <= N0;
    end 
    if(reset_i) begin
      head_r_sv2v_reg <= 1'b0;
    end else if(yumi_i) begin
      head_r_sv2v_reg <= N2;
    end 
  end


endmodule



module bsg_counter_clear_up_f_0_1
(
  clk_i,
  reset_i,
  clear_i,
  up_i,
  count_o
);

  output [3:0] count_o;
  input clk_i;
  input reset_i;
  input clear_i;
  input up_i;
  wire [3:0] count_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10;
  reg count_o_3_sv2v_reg,count_o_2_sv2v_reg,count_o_1_sv2v_reg,count_o_0_sv2v_reg;
  assign count_o[3] = count_o_3_sv2v_reg;
  assign count_o[2] = count_o_2_sv2v_reg;
  assign count_o[1] = count_o_1_sv2v_reg;
  assign count_o[0] = count_o_0_sv2v_reg;
  assign N10 = reset_i | clear_i;
  assign { N8, N7, N6, N5 } = count_o + up_i;
  assign N9 = (N0)? up_i : 
              (N1)? N5 : 1'b0;
  assign N0 = clear_i;
  assign N1 = N4;
  assign N2 = ~reset_i;
  assign N3 = N2;
  assign N4 = ~clear_i;

  always @(posedge clk_i) begin
    if(N10) begin
      count_o_3_sv2v_reg <= 1'b0;
      count_o_2_sv2v_reg <= 1'b0;
      count_o_1_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      count_o_3_sv2v_reg <= N8;
      count_o_2_sv2v_reg <= N7;
      count_o_1_sv2v_reg <= N6;
    end 
    if(reset_i) begin
      count_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      count_o_0_sv2v_reg <= N9;
    end 
  end


endmodule



module bsg_link_source_sync_downstream_channel_width_p16_lg_fifo_depth_p6_lg_credit_to_token_decimation_p3
(
  core_clk_i,
  core_link_reset_i,
  io_link_reset_i,
  io_clk_i,
  io_data_i,
  io_valid_i,
  core_token_r_o,
  core_data_o,
  core_valid_o,
  core_yumi_i
);

  input [15:0] io_data_i;
  output [15:0] core_data_o;
  input core_clk_i;
  input core_link_reset_i;
  input io_link_reset_i;
  input io_clk_i;
  input io_valid_i;
  input core_yumi_i;
  output core_token_r_o;
  output core_valid_o;
  wire [15:0] core_data_o,core_async_fifo_data_lo;
  reg  [15:0] data_commit;
  wire core_token_r_o,core_valid_o,io_async_fifo_full,core_async_fifo_deque,
  core_async_fifo_valid_lo,core_async_fifo_ready_li;
  wire [2:0] core_credits_sent_r;

  always @(posedge core_clk_i) begin
    if(core_async_fifo_deque)
      data_commit <= core_async_fifo_data_lo;
  end 

  bsg_async_fifo_lg_size_p6_width_p16
  baf
  (
    .w_clk_i(io_clk_i),
    .w_reset_i(io_link_reset_i),
    .w_enq_i(io_valid_i),
    .w_data_i(io_data_i),
    .w_full_o(io_async_fifo_full),
    .r_clk_i(core_clk_i),
    .r_reset_i(core_link_reset_i),
    .r_deq_i(core_async_fifo_deque),
    .r_data_o(core_async_fifo_data_lo),
    .r_valid_o(core_async_fifo_valid_lo)
  );


  bsg_two_fifo_width_p16
  twofer
  (
    .clk_i(core_clk_i),
    .reset_i(core_link_reset_i),
    .ready_o(core_async_fifo_ready_li),
    .data_i(core_async_fifo_data_lo),
    .v_i(core_async_fifo_valid_lo),
    .v_o(core_valid_o),
    .data_o(core_data_o),
    .yumi_i(core_yumi_i)
  );


  bsg_counter_clear_up_f_0_1
  token_counter
  (
    .clk_i(core_clk_i),
    .reset_i(core_link_reset_i),
    .clear_i(1'b0),
    .up_i(core_async_fifo_deque),
    .count_o({ core_token_r_o, core_credits_sent_r })
  );

  assign core_async_fifo_deque = core_async_fifo_valid_lo & core_async_fifo_ready_li;

endmodule



module bsg_circular_ptr_slots_p2_max_add_p1
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [0:0] add_i;
  output [0:0] o;
  output [0:0] n_o;
  input clk;
  input reset_i;
  wire [0:0] o,n_o,\genblk1.genblk1.ptr_r_p1 ;
  wire N0,N1,N2;
  reg o_0_sv2v_reg;
  assign o[0] = o_0_sv2v_reg;
  assign \genblk1.genblk1.ptr_r_p1 [0] = o[0] ^ 1'b1;
  assign n_o[0] = (N0)? \genblk1.genblk1.ptr_r_p1 [0] : 
                  (N1)? o[0] : 1'b0;
  assign N0 = add_i[0];
  assign N1 = N2;
  assign N2 = ~add_i[0];

  always @(posedge clk) begin
    if(reset_i) begin
      o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      o_0_sv2v_reg <= n_o[0];
    end 
  end


endmodule



module bsg_round_robin_1_to_n_width_p32_num_out_p2
(
  clk_i,
  reset_i,
  valid_i,
  ready_o,
  valid_o,
  ready_i
);

  output [1:0] valid_o;
  input [1:0] ready_i;
  input clk_i;
  input reset_i;
  input valid_i;
  output ready_o;
  wire [1:0] valid_o;
  wire ready_o,N0,\one_to_n.yumi_i ,N1,sv2v_dc_1;
  wire [0:0] \one_to_n.ptr_r ;

  bsg_circular_ptr_slots_p2_max_add_p1
  one_to_n_circular_ptr 
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(\one_to_n.yumi_i ),
    .o(\one_to_n.ptr_r [0]),
    .n_o(sv2v_dc_1)
  );

  assign valid_o = { 1'b0, valid_i } << \one_to_n.ptr_r [0];
  assign ready_o = (N1)? ready_i[0] : 
                   (N0)? ready_i[1] : 1'b0;
  assign N0 = \one_to_n.ptr_r [0];
  assign \one_to_n.yumi_i  = valid_i & ready_o;
  assign N1 = ~\one_to_n.ptr_r [0];

endmodule



module bsg_mem_1r1w_synth_width_p32_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [31:0] w_data_i;
  input [0:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7;
  wire [63:0] mem;
  reg mem_63_sv2v_reg,mem_62_sv2v_reg,mem_61_sv2v_reg,mem_60_sv2v_reg,mem_59_sv2v_reg,
  mem_58_sv2v_reg,mem_57_sv2v_reg,mem_56_sv2v_reg,mem_55_sv2v_reg,mem_54_sv2v_reg,
  mem_53_sv2v_reg,mem_52_sv2v_reg,mem_51_sv2v_reg,mem_50_sv2v_reg,mem_49_sv2v_reg,
  mem_48_sv2v_reg,mem_47_sv2v_reg,mem_46_sv2v_reg,mem_45_sv2v_reg,mem_44_sv2v_reg,
  mem_43_sv2v_reg,mem_42_sv2v_reg,mem_41_sv2v_reg,mem_40_sv2v_reg,mem_39_sv2v_reg,
  mem_38_sv2v_reg,mem_37_sv2v_reg,mem_36_sv2v_reg,mem_35_sv2v_reg,mem_34_sv2v_reg,
  mem_33_sv2v_reg,mem_32_sv2v_reg,mem_31_sv2v_reg,mem_30_sv2v_reg,mem_29_sv2v_reg,
  mem_28_sv2v_reg,mem_27_sv2v_reg,mem_26_sv2v_reg,mem_25_sv2v_reg,mem_24_sv2v_reg,
  mem_23_sv2v_reg,mem_22_sv2v_reg,mem_21_sv2v_reg,mem_20_sv2v_reg,mem_19_sv2v_reg,
  mem_18_sv2v_reg,mem_17_sv2v_reg,mem_16_sv2v_reg,mem_15_sv2v_reg,mem_14_sv2v_reg,
  mem_13_sv2v_reg,mem_12_sv2v_reg,mem_11_sv2v_reg,mem_10_sv2v_reg,mem_9_sv2v_reg,
  mem_8_sv2v_reg,mem_7_sv2v_reg,mem_6_sv2v_reg,mem_5_sv2v_reg,mem_4_sv2v_reg,
  mem_3_sv2v_reg,mem_2_sv2v_reg,mem_1_sv2v_reg,mem_0_sv2v_reg;
  assign mem[63] = mem_63_sv2v_reg;
  assign mem[62] = mem_62_sv2v_reg;
  assign mem[61] = mem_61_sv2v_reg;
  assign mem[60] = mem_60_sv2v_reg;
  assign mem[59] = mem_59_sv2v_reg;
  assign mem[58] = mem_58_sv2v_reg;
  assign mem[57] = mem_57_sv2v_reg;
  assign mem[56] = mem_56_sv2v_reg;
  assign mem[55] = mem_55_sv2v_reg;
  assign mem[54] = mem_54_sv2v_reg;
  assign mem[53] = mem_53_sv2v_reg;
  assign mem[52] = mem_52_sv2v_reg;
  assign mem[51] = mem_51_sv2v_reg;
  assign mem[50] = mem_50_sv2v_reg;
  assign mem[49] = mem_49_sv2v_reg;
  assign mem[48] = mem_48_sv2v_reg;
  assign mem[47] = mem_47_sv2v_reg;
  assign mem[46] = mem_46_sv2v_reg;
  assign mem[45] = mem_45_sv2v_reg;
  assign mem[44] = mem_44_sv2v_reg;
  assign mem[43] = mem_43_sv2v_reg;
  assign mem[42] = mem_42_sv2v_reg;
  assign mem[41] = mem_41_sv2v_reg;
  assign mem[40] = mem_40_sv2v_reg;
  assign mem[39] = mem_39_sv2v_reg;
  assign mem[38] = mem_38_sv2v_reg;
  assign mem[37] = mem_37_sv2v_reg;
  assign mem[36] = mem_36_sv2v_reg;
  assign mem[35] = mem_35_sv2v_reg;
  assign mem[34] = mem_34_sv2v_reg;
  assign mem[33] = mem_33_sv2v_reg;
  assign mem[32] = mem_32_sv2v_reg;
  assign mem[31] = mem_31_sv2v_reg;
  assign mem[30] = mem_30_sv2v_reg;
  assign mem[29] = mem_29_sv2v_reg;
  assign mem[28] = mem_28_sv2v_reg;
  assign mem[27] = mem_27_sv2v_reg;
  assign mem[26] = mem_26_sv2v_reg;
  assign mem[25] = mem_25_sv2v_reg;
  assign mem[24] = mem_24_sv2v_reg;
  assign mem[23] = mem_23_sv2v_reg;
  assign mem[22] = mem_22_sv2v_reg;
  assign mem[21] = mem_21_sv2v_reg;
  assign mem[20] = mem_20_sv2v_reg;
  assign mem[19] = mem_19_sv2v_reg;
  assign mem[18] = mem_18_sv2v_reg;
  assign mem[17] = mem_17_sv2v_reg;
  assign mem[16] = mem_16_sv2v_reg;
  assign mem[15] = mem_15_sv2v_reg;
  assign mem[14] = mem_14_sv2v_reg;
  assign mem[13] = mem_13_sv2v_reg;
  assign mem[12] = mem_12_sv2v_reg;
  assign mem[11] = mem_11_sv2v_reg;
  assign mem[10] = mem_10_sv2v_reg;
  assign mem[9] = mem_9_sv2v_reg;
  assign mem[8] = mem_8_sv2v_reg;
  assign mem[7] = mem_7_sv2v_reg;
  assign mem[6] = mem_6_sv2v_reg;
  assign mem[5] = mem_5_sv2v_reg;
  assign mem[4] = mem_4_sv2v_reg;
  assign mem[3] = mem_3_sv2v_reg;
  assign mem[2] = mem_2_sv2v_reg;
  assign mem[1] = mem_1_sv2v_reg;
  assign mem[0] = mem_0_sv2v_reg;
  assign r_data_o[31] = (N3)? mem[31] : 
                        (N0)? mem[63] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[30] = (N3)? mem[30] : 
                        (N0)? mem[62] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] : 
                        (N0)? mem[61] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] : 
                        (N0)? mem[60] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] : 
                        (N0)? mem[59] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] : 
                        (N0)? mem[58] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] : 
                        (N0)? mem[57] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] : 
                        (N0)? mem[56] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] : 
                        (N0)? mem[55] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] : 
                        (N0)? mem[54] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] : 
                        (N0)? mem[53] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] : 
                        (N0)? mem[52] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] : 
                        (N0)? mem[51] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] : 
                        (N0)? mem[50] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] : 
                        (N0)? mem[49] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] : 
                        (N0)? mem[48] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] : 
                        (N0)? mem[47] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] : 
                        (N0)? mem[46] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] : 
                        (N0)? mem[45] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] : 
                        (N0)? mem[44] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] : 
                        (N0)? mem[43] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] : 
                        (N0)? mem[42] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] : 
                       (N0)? mem[41] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] : 
                       (N0)? mem[40] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] : 
                       (N0)? mem[39] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] : 
                       (N0)? mem[38] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[37] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[36] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[35] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[34] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[33] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[32] : 1'b0;
  assign N7 = ~w_addr_i[0];
  assign { N6, N5 } = (N1)? { w_addr_i[0:0], N7 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N6) begin
      mem_63_sv2v_reg <= w_data_i[31];
      mem_62_sv2v_reg <= w_data_i[30];
      mem_61_sv2v_reg <= w_data_i[29];
      mem_60_sv2v_reg <= w_data_i[28];
      mem_59_sv2v_reg <= w_data_i[27];
      mem_58_sv2v_reg <= w_data_i[26];
      mem_57_sv2v_reg <= w_data_i[25];
      mem_56_sv2v_reg <= w_data_i[24];
      mem_55_sv2v_reg <= w_data_i[23];
      mem_54_sv2v_reg <= w_data_i[22];
      mem_53_sv2v_reg <= w_data_i[21];
      mem_52_sv2v_reg <= w_data_i[20];
      mem_51_sv2v_reg <= w_data_i[19];
      mem_50_sv2v_reg <= w_data_i[18];
      mem_49_sv2v_reg <= w_data_i[17];
      mem_48_sv2v_reg <= w_data_i[16];
      mem_47_sv2v_reg <= w_data_i[15];
      mem_46_sv2v_reg <= w_data_i[14];
      mem_45_sv2v_reg <= w_data_i[13];
      mem_44_sv2v_reg <= w_data_i[12];
      mem_43_sv2v_reg <= w_data_i[11];
      mem_42_sv2v_reg <= w_data_i[10];
      mem_41_sv2v_reg <= w_data_i[9];
      mem_40_sv2v_reg <= w_data_i[8];
      mem_39_sv2v_reg <= w_data_i[7];
      mem_38_sv2v_reg <= w_data_i[6];
      mem_37_sv2v_reg <= w_data_i[5];
      mem_36_sv2v_reg <= w_data_i[4];
      mem_35_sv2v_reg <= w_data_i[3];
      mem_34_sv2v_reg <= w_data_i[2];
      mem_33_sv2v_reg <= w_data_i[1];
      mem_32_sv2v_reg <= w_data_i[0];
    end 
    if(N5) begin
      mem_31_sv2v_reg <= w_data_i[31];
      mem_30_sv2v_reg <= w_data_i[30];
      mem_29_sv2v_reg <= w_data_i[29];
      mem_28_sv2v_reg <= w_data_i[28];
      mem_27_sv2v_reg <= w_data_i[27];
      mem_26_sv2v_reg <= w_data_i[26];
      mem_25_sv2v_reg <= w_data_i[25];
      mem_24_sv2v_reg <= w_data_i[24];
      mem_23_sv2v_reg <= w_data_i[23];
      mem_22_sv2v_reg <= w_data_i[22];
      mem_21_sv2v_reg <= w_data_i[21];
      mem_20_sv2v_reg <= w_data_i[20];
      mem_19_sv2v_reg <= w_data_i[19];
      mem_18_sv2v_reg <= w_data_i[18];
      mem_17_sv2v_reg <= w_data_i[17];
      mem_16_sv2v_reg <= w_data_i[16];
      mem_15_sv2v_reg <= w_data_i[15];
      mem_14_sv2v_reg <= w_data_i[14];
      mem_13_sv2v_reg <= w_data_i[13];
      mem_12_sv2v_reg <= w_data_i[12];
      mem_11_sv2v_reg <= w_data_i[11];
      mem_10_sv2v_reg <= w_data_i[10];
      mem_9_sv2v_reg <= w_data_i[9];
      mem_8_sv2v_reg <= w_data_i[8];
      mem_7_sv2v_reg <= w_data_i[7];
      mem_6_sv2v_reg <= w_data_i[6];
      mem_5_sv2v_reg <= w_data_i[5];
      mem_4_sv2v_reg <= w_data_i[4];
      mem_3_sv2v_reg <= w_data_i[3];
      mem_2_sv2v_reg <= w_data_i[2];
      mem_1_sv2v_reg <= w_data_i[1];
      mem_0_sv2v_reg <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p32_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [31:0] w_data_i;
  input [0:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;

  bsg_mem_1r1w_synth_width_p32_els_p2_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p32
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,enq_i,tail_r,_0_net_,head_r,empty_r,full_r,N0,N1,N2,N3,N4,N5,N6,N7,
  N8,N9,N10,N11,N12,N13,N14;
  reg full_r_sv2v_reg,tail_r_sv2v_reg,head_r_sv2v_reg,empty_r_sv2v_reg;
  assign full_r = full_r_sv2v_reg;
  assign tail_r = tail_r_sv2v_reg;
  assign head_r = head_r_sv2v_reg;
  assign empty_r = empty_r_sv2v_reg;

  bsg_mem_1r1w_width_p32_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign _0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N5;
  assign N5 = ~full_r;
  assign N1 = enq_i;
  assign N0 = ~tail_r;
  assign N2 = ~head_r;
  assign N3 = N7 | N9;
  assign N7 = empty_r & N6;
  assign N6 = ~enq_i;
  assign N9 = N8 & N6;
  assign N8 = N5 & yumi_i;
  assign N4 = N13 | N14;
  assign N13 = N11 & N12;
  assign N11 = N10 & enq_i;
  assign N10 = ~empty_r;
  assign N12 = ~yumi_i;
  assign N14 = full_r & N12;

  always @(posedge clk_i) begin
    if(reset_i) begin
      full_r_sv2v_reg <= 1'b0;
      empty_r_sv2v_reg <= 1'b1;
    end else if(1'b1) begin
      full_r_sv2v_reg <= N4;
      empty_r_sv2v_reg <= N3;
    end 
    if(reset_i) begin
      tail_r_sv2v_reg <= 1'b0;
    end else if(N1) begin
      tail_r_sv2v_reg <= N0;
    end 
    if(reset_i) begin
      head_r_sv2v_reg <= 1'b0;
    end else if(yumi_i) begin
      head_r_sv2v_reg <= N2;
    end 
  end


endmodule



module bsg_dff_reset_width_p1
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  input reset_i;
  wire [0:0] data_o;
  reg data_o_0_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_width_p32_harden_p0
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input en_i;
  wire [31:0] data_o;
  reg data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,
  data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,
  data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,
  data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,
  data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_one_fifo_width_p32
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,N0,N1,_0_net_,N2,N3,_1_net_;

  bsg_dff_reset_width_p1
  dff_full
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(_0_net_),
    .data_o(v_o)
  );


  bsg_dff_en_width_p32_harden_p0
  dff
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .en_i(_1_net_),
    .data_o(data_o)
  );

  assign _0_net_ = (N0)? N3 : 
                   (N1)? v_i : 1'b0;
  assign N0 = v_o;
  assign N1 = N2;
  assign ready_o = ~v_o;
  assign N2 = ~v_o;
  assign N3 = ~yumi_i;
  assign _1_net_ = v_i & ready_o;

endmodule



module bsg_serial_in_parallel_out_full_width_p32_els_p2
(
  clk_i,
  reset_i,
  v_i,
  ready_o,
  data_i,
  data_o,
  v_o,
  yumi_i
);

  input [31:0] data_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [63:0] data_o;
  wire ready_o,v_o;
  wire [1:0] fifo_valid_lo,fifo_valid_li,fifo_ready_lo;

  bsg_round_robin_1_to_n_width_p32_num_out_p2
  brr
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .valid_i(v_i),
    .ready_o(ready_o),
    .valid_o(fifo_valid_li),
    .ready_i(fifo_ready_lo)
  );


  bsg_two_fifo_width_p32
  fifos_0_twofifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(fifo_ready_lo[0]),
    .data_i(data_i),
    .v_i(fifo_valid_li[0]),
    .v_o(fifo_valid_lo[0]),
    .data_o(data_o[31:0]),
    .yumi_i(yumi_i)
  );


  bsg_one_fifo_width_p32
  fifos_1_onefifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(fifo_ready_lo[1]),
    .data_i(data_i),
    .v_i(fifo_valid_li[1]),
    .v_o(fifo_valid_lo[1]),
    .data_o(data_o[63:32]),
    .yumi_i(yumi_i)
  );

  assign v_o = fifo_valid_lo[1] & fifo_valid_lo[0];

endmodule



module bsg_link_ddr_downstream
(
  core_clk_i,
  core_link_reset_i,
  io_link_reset_i,
  core_data_o,
  core_valid_o,
  core_yumi_i,
  io_clk_i,
  io_data_i,
  io_valid_i,
  core_token_r_o
);

  input io_link_reset_i;
  output [63:0] core_data_o;
  input io_clk_i;
  input [15:0] io_data_i;
  input io_valid_i;
  output [1:0] core_token_r_o;
  input core_clk_i;
  input core_link_reset_i;
  input core_yumi_i;
  output core_valid_o;
  wire [63:0] core_data_o;
  wire [1:0] core_token_r_o,core_sipo_valid_li;
  wire core_valid_o,core_sipo_ready_lo,core_sipo_yumi_lo,\ch_0_.io_iddr_v_lo ,
  \ch_1_.io_iddr_v_lo ,_6_net_,N0;
  wire [8:0] \ch_0_.io_iddr_data_top ,\ch_1_.io_iddr_data_top ;
  wire [7:0] \ch_0_.io_iddr_data_bottom ,\ch_1_.io_iddr_data_bottom ;
  wire [31:0] core_sipo_data_li;

  bsg_link_iddr_phy_width_p9
  ch_0_iddr_data 
  (
    .clk_i(io_clk_i),
    .data_i({ io_valid_i, io_data_i[7:0] }),
    .data_r_o({ \ch_0_.io_iddr_data_top , \ch_0_.io_iddr_v_lo , \ch_0_.io_iddr_data_bottom  }),
    .rst(io_link_reset_i)
  );


  bsg_link_source_sync_downstream_channel_width_p16_lg_fifo_depth_p6_lg_credit_to_token_decimation_p3
  ch_0_downstream 
  (
    .core_clk_i(core_clk_i),
    .core_link_reset_i(core_link_reset_i),
    .io_link_reset_i(io_link_reset_i),
    .io_clk_i(io_clk_i),
    .io_data_i({ \ch_0_.io_iddr_data_top [7:0], \ch_0_.io_iddr_data_bottom  }),
    .io_valid_i(\ch_0_.io_iddr_v_lo ),
    .core_token_r_o(core_token_r_o[0]),
    .core_data_o(core_sipo_data_li[15:0]),
    .core_valid_o(core_sipo_valid_li[0]),
    .core_yumi_i(core_sipo_yumi_lo)
  );


  bsg_link_iddr_phy_width_p9
  ch_1_iddr_data 
  (
    .clk_i(io_clk_i),
    .data_i({ io_valid_i, io_data_i[15:8] }),
    .data_r_o({ \ch_1_.io_iddr_data_top , \ch_1_.io_iddr_v_lo , \ch_1_.io_iddr_data_bottom  }),
    .rst(io_link_reset_i)
  );


  bsg_link_source_sync_downstream_channel_width_p16_lg_fifo_depth_p6_lg_credit_to_token_decimation_p3
  ch_1_downstream 
  (
    .core_clk_i(core_clk_i),
    .core_link_reset_i(core_link_reset_i),
    .io_link_reset_i(io_link_reset_i),
    .io_clk_i(io_clk_i),
    .io_data_i({ \ch_1_.io_iddr_data_top [7:0], \ch_1_.io_iddr_data_bottom  }),
    .io_valid_i(\ch_1_.io_iddr_v_lo ),
    .core_token_r_o(core_token_r_o[1]),
    .core_data_o(core_sipo_data_li[31:16]),
    .core_valid_o(core_sipo_valid_li[1]),
    .core_yumi_i(core_sipo_yumi_lo)
  );


  bsg_serial_in_parallel_out_full_width_p32_els_p2
  in_sipof
  (
    .clk_i(core_clk_i),
    .reset_i(core_link_reset_i),
    .v_i(_6_net_),
    .ready_o(core_sipo_ready_lo),
    .data_i(core_sipo_data_li),
    .data_o(core_data_o),
    .v_o(core_valid_o),
    .yumi_i(core_yumi_i)
  );


  assign core_sipo_yumi_lo = N0 & core_sipo_ready_lo;
  assign N0 = core_sipo_valid_li[1] & core_sipo_valid_li[0];
  assign _6_net_ = core_sipo_valid_li[1] & core_sipo_valid_li[0];

endmodule
