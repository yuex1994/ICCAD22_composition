
//------> ./PECore_ccs_conn_in_wait_v1.v 
module PECore_ccs_conn_in_wait_v1 (
  vld, rdy, dat, idat, irdy, ivld, clk, en, arst, srst
);

  parameter integer width = 32;
  parameter integer ph_clk  = 1;
  parameter integer ph_en   = 1;
  parameter integer ph_arst = 1;
  parameter integer ph_srst = 1;
  //parameter         has_en  = 1'b1;
  input [width-1:0] dat;
  input vld;
  output rdy;
  output [width-1:0] idat;
  input irdy;
  output ivld;
  input clk;
  input en;
  input arst;
  input srst;

  localparam stallOff = 0;
  wire                  stall_ctrl;
  assign stall_ctrl = stallOff;

  assign idat = dat;
  assign rdy = irdy && !stall_ctrl;
  assign ivld = vld && !stall_ctrl;
endmodule




//------> ./PECore_ccs_conn_out_wait_v1.v 
module PECore_ccs_conn_out_wait_v1 (
  vld, rdy, dat, idat, ivld, irdy,
      clk, en, arst, srst
);
  parameter integer width = 32;
  parameter integer ph_clk  = 1;
  parameter integer ph_en  = 1;
  parameter integer ph_arst = 1;
  parameter integer ph_srst = 1;
  //parameter         has_en  = 1'b1;
  output [width-1:0] dat;
  output vld;
  input rdy;
  input [width-1:0] idat;
  input ivld;
  output irdy;
  input clk;
  input en;
  input arst;
  input srst;

  localparam stallOff = 0;
  wire stall_ctrl;
  assign stall_ctrl = stallOff;

  assign dat = idat;
  assign vld = ivld && !stall_ctrl;
  assign irdy = rdy && !stall_ctrl;

endmodule




//------> ./PECore_ProductSum_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_ProductSum_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_ProductSum_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_ProductSum_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./PECore_ProductSum_mgc_shift_l_beh_v5.v 
module PECore_ProductSum_mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./PECore_ProductSum_ACC_16i25_1o29_6c39adcf8fa7ac08d026ec7c525fe9f9e6.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.6a/933210 Production Release
//  HLS Date:       Mon Apr 12 07:56:29 PDT 2021
//
//  Generated date: Wed Mar 30 23:27:46 2022
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    ACC_16i25_1o29_6c39adcf8fa7ac08d026ec7c525fe9f9e6
// ------------------------------------------------------------------


module PECore_ProductSum_ACC_16i25_1o29_6c39adcf8fa7ac08d026ec7c525fe9f9e6 (
  I_1, I_2, I_3, I_4, I_5, I_6, I_7, I_8, I_9, I_10, I_11, I_12, I_13, I_14, I_15,
      I_16, O_1
);
  input [24:0] I_1;
  input [24:0] I_2;
  input [24:0] I_3;
  input [24:0] I_4;
  input [24:0] I_5;
  input [24:0] I_6;
  input [24:0] I_7;
  input [24:0] I_8;
  input [24:0] I_9;
  input [24:0] I_10;
  input [24:0] I_11;
  input [24:0] I_12;
  input [24:0] I_13;
  input [24:0] I_14;
  input [24:0] I_15;
  input [24:0] I_16;
  output [28:0] O_1;
  wire [32:0] nl_O_1;



  // Interconnect Declarations for Component Instantiations
  assign nl_O_1 = conv_s2s_25_29(I_4) + conv_s2s_25_29(I_5) + conv_s2s_25_29(I_6)
      + conv_s2s_25_29(I_7) + conv_s2s_25_29(I_8) + conv_s2s_25_29(I_9) + conv_s2s_25_29(I_10)
      + conv_s2s_25_29(I_11) + conv_s2s_25_29(I_12) + conv_s2s_25_29(I_1) + conv_s2s_25_29(I_2)
      + conv_s2s_25_29(I_3) + conv_s2s_25_29(I_13) + conv_s2s_25_29(I_14) + conv_s2s_25_29(I_15)
      + conv_s2s_25_29(I_16);
  assign O_1 = nl_O_1[28:0];

  function automatic [28:0] conv_s2s_25_29 ;
    input [24:0]  vector ;
  begin
    conv_s2s_25_29 = {{4{vector[24]}}, vector};
  end
  endfunction

endmodule




//------> ./PECore_ProductSum.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.6a/933210 Production Release
//  HLS Date:       Mon Apr 12 07:56:29 PDT 2021
//
//  Generated date: Wed Mar 30 23:29:06 2022
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    ProductSum_ProductSum_core
// ------------------------------------------------------------------


module PECore_ProductSum_ProductSum_core (
  in_1_data_rsc_dat, in_2_data_rsc_dat, out_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_arst, ccs_ccore_en
);
  input [127:0] in_1_data_rsc_dat;
  input [127:0] in_2_data_rsc_dat;
  output [31:0] out_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [127:0] in_1_data_rsci_idat;
  wire [127:0] in_2_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [28:0] out_rsci_d_28_0;
  wire [24:0] for_10_adpfloat_mul_template_8U_3U_32U_lshift_itm;
  wire [24:0] for_11_adpfloat_mul_template_8U_3U_32U_lshift_itm;
  wire [24:0] for_12_adpfloat_mul_template_8U_3U_32U_lshift_itm;
  wire [24:0] for_13_adpfloat_mul_template_8U_3U_32U_lshift_itm;
  wire [24:0] for_14_adpfloat_mul_template_8U_3U_32U_lshift_itm;
  wire [24:0] for_15_adpfloat_mul_template_8U_3U_32U_lshift_itm;
  wire [24:0] for_16_adpfloat_mul_template_8U_3U_32U_lshift_itm;
  wire [24:0] for_1_adpfloat_mul_template_8U_3U_32U_lshift_itm;
  wire [24:0] for_2_adpfloat_mul_template_8U_3U_32U_lshift_itm;
  wire [24:0] for_3_adpfloat_mul_template_8U_3U_32U_lshift_itm;
  wire [24:0] for_4_adpfloat_mul_template_8U_3U_32U_lshift_itm;
  wire [24:0] for_5_adpfloat_mul_template_8U_3U_32U_lshift_itm;
  wire [24:0] for_6_adpfloat_mul_template_8U_3U_32U_lshift_itm;
  wire [24:0] for_7_adpfloat_mul_template_8U_3U_32U_lshift_itm;
  wire [24:0] for_8_adpfloat_mul_template_8U_3U_32U_lshift_itm;
  wire [24:0] for_9_adpfloat_mul_template_8U_3U_32U_lshift_itm;
  wire [10:0] adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_1_sva_1;
  wire [11:0] nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_1_sva_1;
  wire [9:0] adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_1_sva_1;
  wire [10:0] adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_2_sva_1;
  wire [11:0] nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_2_sva_1;
  wire [9:0] adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_2_sva_1;
  wire [10:0] adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_3_sva_1;
  wire [11:0] nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_3_sva_1;
  wire [9:0] adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_3_sva_1;
  wire [10:0] adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_4_sva_1;
  wire [11:0] nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_4_sva_1;
  wire [9:0] adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_4_sva_1;
  wire [10:0] adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_5_sva_1;
  wire [11:0] nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_5_sva_1;
  wire [9:0] adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_5_sva_1;
  wire [10:0] adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_6_sva_1;
  wire [11:0] nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_6_sva_1;
  wire [9:0] adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_6_sva_1;
  wire [10:0] adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_7_sva_1;
  wire [11:0] nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_7_sva_1;
  wire [9:0] adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_7_sva_1;
  wire [10:0] adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_8_sva_1;
  wire [11:0] nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_8_sva_1;
  wire [9:0] adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_8_sva_1;
  wire [10:0] adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_9_sva_1;
  wire [11:0] nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_9_sva_1;
  wire [9:0] adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_9_sva_1;
  wire [10:0] adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_10_sva_1;
  wire [11:0] nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_10_sva_1;
  wire [9:0] adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_10_sva_1;
  wire [10:0] adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_11_sva_1;
  wire [11:0] nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_11_sva_1;
  wire [9:0] adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_11_sva_1;
  wire [10:0] adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_12_sva_1;
  wire [11:0] nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_12_sva_1;
  wire [9:0] adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_12_sva_1;
  wire [10:0] adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_13_sva_1;
  wire [11:0] nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_13_sva_1;
  wire [9:0] adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_13_sva_1;
  wire [10:0] adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_14_sva_1;
  wire [11:0] nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_14_sva_1;
  wire [9:0] adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_14_sva_1;
  wire [10:0] adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_15_sva_1;
  wire [11:0] nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_15_sva_1;
  wire [9:0] adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_15_sva_1;
  wire [10:0] adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_sva_1;
  wire [11:0] nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_sva_1;
  wire [9:0] adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_sva_1;
  wire for_10_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  wire for_11_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  wire for_12_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  wire for_13_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  wire for_14_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  wire for_15_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  wire for_16_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  wire for_1_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  wire for_2_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  wire for_3_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  wire for_4_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  wire for_5_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  wire for_6_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  wire for_7_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  wire for_8_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  wire for_9_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  wire [28:0] ACC_16i25_1o29_c7aa682b5659f7f20224ec66be5b70f85d_1;

  wire for_1_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl;
  wire for_1_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl;
  wire for_2_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl;
  wire for_2_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl;
  wire for_3_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl;
  wire for_3_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl;
  wire for_4_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl;
  wire for_4_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl;
  wire for_5_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl;
  wire for_5_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl;
  wire for_6_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl;
  wire for_6_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl;
  wire for_7_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl;
  wire for_7_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl;
  wire for_8_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl;
  wire for_8_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl;
  wire for_9_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl;
  wire for_9_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl;
  wire for_10_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl;
  wire for_10_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl;
  wire for_11_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl;
  wire for_11_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl;
  wire for_12_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl;
  wire for_12_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl;
  wire for_13_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl;
  wire for_13_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl;
  wire for_14_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl;
  wire for_14_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl;
  wire for_15_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl;
  wire for_15_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl;
  wire for_16_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl;
  wire for_16_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl;

  // Interconnect Declarations for Component Instantiations
  wire [31:0] nl_out_rsci_d;
  assign nl_out_rsci_d = {{3{out_rsci_d_28_0[28]}}, out_rsci_d_28_0};
  wire adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_9_nl;
  wire[9:0] adpfloat_mul_template_8U_3U_32U_mux_29_nl;
  wire [10:0] nl_for_10_adpfloat_mul_template_8U_3U_32U_lshift_rg_a;
  assign adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_9_nl
      = (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_10_sva_1[10]) & for_10_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  assign adpfloat_mul_template_8U_3U_32U_mux_29_nl = MUX_v_10_2_2(adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_10_sva_1,
      (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_10_sva_1[9:0]), for_10_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1);
  assign nl_for_10_adpfloat_mul_template_8U_3U_32U_lshift_rg_a = {adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_9_nl
      , adpfloat_mul_template_8U_3U_32U_mux_29_nl};
  wire [3:0] nl_for_10_adpfloat_mul_template_8U_3U_32U_lshift_rg_s;
  assign nl_for_10_adpfloat_mul_template_8U_3U_32U_lshift_rg_s = conv_u2u_3_4(in_1_data_rsci_idat[78:76])
      + conv_u2u_3_4(in_2_data_rsci_idat[78:76]);
  wire adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_10_nl;
  wire[9:0] adpfloat_mul_template_8U_3U_32U_mux_32_nl;
  wire [10:0] nl_for_11_adpfloat_mul_template_8U_3U_32U_lshift_rg_a;
  assign adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_10_nl
      = (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_11_sva_1[10]) & for_11_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  assign adpfloat_mul_template_8U_3U_32U_mux_32_nl = MUX_v_10_2_2(adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_11_sva_1,
      (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_11_sva_1[9:0]), for_11_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1);
  assign nl_for_11_adpfloat_mul_template_8U_3U_32U_lshift_rg_a = {adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_10_nl
      , adpfloat_mul_template_8U_3U_32U_mux_32_nl};
  wire [3:0] nl_for_11_adpfloat_mul_template_8U_3U_32U_lshift_rg_s;
  assign nl_for_11_adpfloat_mul_template_8U_3U_32U_lshift_rg_s = conv_u2u_3_4(in_1_data_rsci_idat[86:84])
      + conv_u2u_3_4(in_2_data_rsci_idat[86:84]);
  wire adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_11_nl;
  wire[9:0] adpfloat_mul_template_8U_3U_32U_mux_35_nl;
  wire [10:0] nl_for_12_adpfloat_mul_template_8U_3U_32U_lshift_rg_a;
  assign adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_11_nl
      = (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_12_sva_1[10]) & for_12_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  assign adpfloat_mul_template_8U_3U_32U_mux_35_nl = MUX_v_10_2_2(adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_12_sva_1,
      (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_12_sva_1[9:0]), for_12_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1);
  assign nl_for_12_adpfloat_mul_template_8U_3U_32U_lshift_rg_a = {adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_11_nl
      , adpfloat_mul_template_8U_3U_32U_mux_35_nl};
  wire [3:0] nl_for_12_adpfloat_mul_template_8U_3U_32U_lshift_rg_s;
  assign nl_for_12_adpfloat_mul_template_8U_3U_32U_lshift_rg_s = conv_u2u_3_4(in_1_data_rsci_idat[94:92])
      + conv_u2u_3_4(in_2_data_rsci_idat[94:92]);
  wire adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_12_nl;
  wire[9:0] adpfloat_mul_template_8U_3U_32U_mux_38_nl;
  wire [10:0] nl_for_13_adpfloat_mul_template_8U_3U_32U_lshift_rg_a;
  assign adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_12_nl
      = (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_13_sva_1[10]) & for_13_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  assign adpfloat_mul_template_8U_3U_32U_mux_38_nl = MUX_v_10_2_2(adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_13_sva_1,
      (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_13_sva_1[9:0]), for_13_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1);
  assign nl_for_13_adpfloat_mul_template_8U_3U_32U_lshift_rg_a = {adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_12_nl
      , adpfloat_mul_template_8U_3U_32U_mux_38_nl};
  wire [3:0] nl_for_13_adpfloat_mul_template_8U_3U_32U_lshift_rg_s;
  assign nl_for_13_adpfloat_mul_template_8U_3U_32U_lshift_rg_s = conv_u2u_3_4(in_1_data_rsci_idat[102:100])
      + conv_u2u_3_4(in_2_data_rsci_idat[102:100]);
  wire adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_13_nl;
  wire[9:0] adpfloat_mul_template_8U_3U_32U_mux_41_nl;
  wire [10:0] nl_for_14_adpfloat_mul_template_8U_3U_32U_lshift_rg_a;
  assign adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_13_nl
      = (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_14_sva_1[10]) & for_14_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  assign adpfloat_mul_template_8U_3U_32U_mux_41_nl = MUX_v_10_2_2(adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_14_sva_1,
      (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_14_sva_1[9:0]), for_14_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1);
  assign nl_for_14_adpfloat_mul_template_8U_3U_32U_lshift_rg_a = {adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_13_nl
      , adpfloat_mul_template_8U_3U_32U_mux_41_nl};
  wire [3:0] nl_for_14_adpfloat_mul_template_8U_3U_32U_lshift_rg_s;
  assign nl_for_14_adpfloat_mul_template_8U_3U_32U_lshift_rg_s = conv_u2u_3_4(in_1_data_rsci_idat[110:108])
      + conv_u2u_3_4(in_2_data_rsci_idat[110:108]);
  wire adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_14_nl;
  wire[9:0] adpfloat_mul_template_8U_3U_32U_mux_44_nl;
  wire [10:0] nl_for_15_adpfloat_mul_template_8U_3U_32U_lshift_rg_a;
  assign adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_14_nl
      = (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_15_sva_1[10]) & for_15_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  assign adpfloat_mul_template_8U_3U_32U_mux_44_nl = MUX_v_10_2_2(adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_15_sva_1,
      (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_15_sva_1[9:0]), for_15_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1);
  assign nl_for_15_adpfloat_mul_template_8U_3U_32U_lshift_rg_a = {adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_14_nl
      , adpfloat_mul_template_8U_3U_32U_mux_44_nl};
  wire [3:0] nl_for_15_adpfloat_mul_template_8U_3U_32U_lshift_rg_s;
  assign nl_for_15_adpfloat_mul_template_8U_3U_32U_lshift_rg_s = conv_u2u_3_4(in_1_data_rsci_idat[118:116])
      + conv_u2u_3_4(in_2_data_rsci_idat[118:116]);
  wire adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_15_nl;
  wire[9:0] adpfloat_mul_template_8U_3U_32U_mux_47_nl;
  wire [10:0] nl_for_16_adpfloat_mul_template_8U_3U_32U_lshift_rg_a;
  assign adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_15_nl
      = (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_sva_1[10]) & for_16_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  assign adpfloat_mul_template_8U_3U_32U_mux_47_nl = MUX_v_10_2_2(adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_sva_1,
      (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_sva_1[9:0]), for_16_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1);
  assign nl_for_16_adpfloat_mul_template_8U_3U_32U_lshift_rg_a = {adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_15_nl
      , adpfloat_mul_template_8U_3U_32U_mux_47_nl};
  wire [3:0] nl_for_16_adpfloat_mul_template_8U_3U_32U_lshift_rg_s;
  assign nl_for_16_adpfloat_mul_template_8U_3U_32U_lshift_rg_s = conv_u2u_3_4(in_1_data_rsci_idat[126:124])
      + conv_u2u_3_4(in_2_data_rsci_idat[126:124]);
  wire adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_nl;
  wire[9:0] adpfloat_mul_template_8U_3U_32U_mux_2_nl;
  wire [10:0] nl_for_1_adpfloat_mul_template_8U_3U_32U_lshift_rg_a;
  assign adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_nl =
      (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_1_sva_1[10]) & for_1_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  assign adpfloat_mul_template_8U_3U_32U_mux_2_nl = MUX_v_10_2_2(adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_1_sva_1,
      (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_1_sva_1[9:0]), for_1_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1);
  assign nl_for_1_adpfloat_mul_template_8U_3U_32U_lshift_rg_a = {adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_nl
      , adpfloat_mul_template_8U_3U_32U_mux_2_nl};
  wire [3:0] nl_for_1_adpfloat_mul_template_8U_3U_32U_lshift_rg_s;
  assign nl_for_1_adpfloat_mul_template_8U_3U_32U_lshift_rg_s = conv_u2u_3_4(in_1_data_rsci_idat[6:4])
      + conv_u2u_3_4(in_2_data_rsci_idat[6:4]);
  wire adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_1_nl;
  wire[9:0] adpfloat_mul_template_8U_3U_32U_mux_5_nl;
  wire [10:0] nl_for_2_adpfloat_mul_template_8U_3U_32U_lshift_rg_a;
  assign adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_1_nl
      = (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_2_sva_1[10]) & for_2_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  assign adpfloat_mul_template_8U_3U_32U_mux_5_nl = MUX_v_10_2_2(adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_2_sva_1,
      (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_2_sva_1[9:0]), for_2_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1);
  assign nl_for_2_adpfloat_mul_template_8U_3U_32U_lshift_rg_a = {adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_1_nl
      , adpfloat_mul_template_8U_3U_32U_mux_5_nl};
  wire [3:0] nl_for_2_adpfloat_mul_template_8U_3U_32U_lshift_rg_s;
  assign nl_for_2_adpfloat_mul_template_8U_3U_32U_lshift_rg_s = conv_u2u_3_4(in_1_data_rsci_idat[14:12])
      + conv_u2u_3_4(in_2_data_rsci_idat[14:12]);
  wire adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_2_nl;
  wire[9:0] adpfloat_mul_template_8U_3U_32U_mux_8_nl;
  wire [10:0] nl_for_3_adpfloat_mul_template_8U_3U_32U_lshift_rg_a;
  assign adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_2_nl
      = (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_3_sva_1[10]) & for_3_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  assign adpfloat_mul_template_8U_3U_32U_mux_8_nl = MUX_v_10_2_2(adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_3_sva_1,
      (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_3_sva_1[9:0]), for_3_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1);
  assign nl_for_3_adpfloat_mul_template_8U_3U_32U_lshift_rg_a = {adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_2_nl
      , adpfloat_mul_template_8U_3U_32U_mux_8_nl};
  wire [3:0] nl_for_3_adpfloat_mul_template_8U_3U_32U_lshift_rg_s;
  assign nl_for_3_adpfloat_mul_template_8U_3U_32U_lshift_rg_s = conv_u2u_3_4(in_1_data_rsci_idat[22:20])
      + conv_u2u_3_4(in_2_data_rsci_idat[22:20]);
  wire adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_3_nl;
  wire[9:0] adpfloat_mul_template_8U_3U_32U_mux_11_nl;
  wire [10:0] nl_for_4_adpfloat_mul_template_8U_3U_32U_lshift_rg_a;
  assign adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_3_nl
      = (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_4_sva_1[10]) & for_4_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  assign adpfloat_mul_template_8U_3U_32U_mux_11_nl = MUX_v_10_2_2(adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_4_sva_1,
      (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_4_sva_1[9:0]), for_4_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1);
  assign nl_for_4_adpfloat_mul_template_8U_3U_32U_lshift_rg_a = {adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_3_nl
      , adpfloat_mul_template_8U_3U_32U_mux_11_nl};
  wire [3:0] nl_for_4_adpfloat_mul_template_8U_3U_32U_lshift_rg_s;
  assign nl_for_4_adpfloat_mul_template_8U_3U_32U_lshift_rg_s = conv_u2u_3_4(in_1_data_rsci_idat[30:28])
      + conv_u2u_3_4(in_2_data_rsci_idat[30:28]);
  wire adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_4_nl;
  wire[9:0] adpfloat_mul_template_8U_3U_32U_mux_14_nl;
  wire [10:0] nl_for_5_adpfloat_mul_template_8U_3U_32U_lshift_rg_a;
  assign adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_4_nl
      = (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_5_sva_1[10]) & for_5_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  assign adpfloat_mul_template_8U_3U_32U_mux_14_nl = MUX_v_10_2_2(adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_5_sva_1,
      (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_5_sva_1[9:0]), for_5_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1);
  assign nl_for_5_adpfloat_mul_template_8U_3U_32U_lshift_rg_a = {adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_4_nl
      , adpfloat_mul_template_8U_3U_32U_mux_14_nl};
  wire [3:0] nl_for_5_adpfloat_mul_template_8U_3U_32U_lshift_rg_s;
  assign nl_for_5_adpfloat_mul_template_8U_3U_32U_lshift_rg_s = conv_u2u_3_4(in_1_data_rsci_idat[38:36])
      + conv_u2u_3_4(in_2_data_rsci_idat[38:36]);
  wire adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_5_nl;
  wire[9:0] adpfloat_mul_template_8U_3U_32U_mux_17_nl;
  wire [10:0] nl_for_6_adpfloat_mul_template_8U_3U_32U_lshift_rg_a;
  assign adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_5_nl
      = (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_6_sva_1[10]) & for_6_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  assign adpfloat_mul_template_8U_3U_32U_mux_17_nl = MUX_v_10_2_2(adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_6_sva_1,
      (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_6_sva_1[9:0]), for_6_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1);
  assign nl_for_6_adpfloat_mul_template_8U_3U_32U_lshift_rg_a = {adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_5_nl
      , adpfloat_mul_template_8U_3U_32U_mux_17_nl};
  wire [3:0] nl_for_6_adpfloat_mul_template_8U_3U_32U_lshift_rg_s;
  assign nl_for_6_adpfloat_mul_template_8U_3U_32U_lshift_rg_s = conv_u2u_3_4(in_1_data_rsci_idat[46:44])
      + conv_u2u_3_4(in_2_data_rsci_idat[46:44]);
  wire adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_6_nl;
  wire[9:0] adpfloat_mul_template_8U_3U_32U_mux_20_nl;
  wire [10:0] nl_for_7_adpfloat_mul_template_8U_3U_32U_lshift_rg_a;
  assign adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_6_nl
      = (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_7_sva_1[10]) & for_7_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  assign adpfloat_mul_template_8U_3U_32U_mux_20_nl = MUX_v_10_2_2(adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_7_sva_1,
      (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_7_sva_1[9:0]), for_7_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1);
  assign nl_for_7_adpfloat_mul_template_8U_3U_32U_lshift_rg_a = {adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_6_nl
      , adpfloat_mul_template_8U_3U_32U_mux_20_nl};
  wire [3:0] nl_for_7_adpfloat_mul_template_8U_3U_32U_lshift_rg_s;
  assign nl_for_7_adpfloat_mul_template_8U_3U_32U_lshift_rg_s = conv_u2u_3_4(in_1_data_rsci_idat[54:52])
      + conv_u2u_3_4(in_2_data_rsci_idat[54:52]);
  wire adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_7_nl;
  wire[9:0] adpfloat_mul_template_8U_3U_32U_mux_23_nl;
  wire [10:0] nl_for_8_adpfloat_mul_template_8U_3U_32U_lshift_rg_a;
  assign adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_7_nl
      = (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_8_sva_1[10]) & for_8_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  assign adpfloat_mul_template_8U_3U_32U_mux_23_nl = MUX_v_10_2_2(adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_8_sva_1,
      (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_8_sva_1[9:0]), for_8_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1);
  assign nl_for_8_adpfloat_mul_template_8U_3U_32U_lshift_rg_a = {adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_7_nl
      , adpfloat_mul_template_8U_3U_32U_mux_23_nl};
  wire [3:0] nl_for_8_adpfloat_mul_template_8U_3U_32U_lshift_rg_s;
  assign nl_for_8_adpfloat_mul_template_8U_3U_32U_lshift_rg_s = conv_u2u_3_4(in_1_data_rsci_idat[62:60])
      + conv_u2u_3_4(in_2_data_rsci_idat[62:60]);
  wire adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_8_nl;
  wire[9:0] adpfloat_mul_template_8U_3U_32U_mux_26_nl;
  wire [10:0] nl_for_9_adpfloat_mul_template_8U_3U_32U_lshift_rg_a;
  assign adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_8_nl
      = (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_9_sva_1[10]) & for_9_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1;
  assign adpfloat_mul_template_8U_3U_32U_mux_26_nl = MUX_v_10_2_2(adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_9_sva_1,
      (adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_9_sva_1[9:0]), for_9_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1);
  assign nl_for_9_adpfloat_mul_template_8U_3U_32U_lshift_rg_a = {adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_and_8_nl
      , adpfloat_mul_template_8U_3U_32U_mux_26_nl};
  wire [3:0] nl_for_9_adpfloat_mul_template_8U_3U_32U_lshift_rg_s;
  assign nl_for_9_adpfloat_mul_template_8U_3U_32U_lshift_rg_s = conv_u2u_3_4(in_1_data_rsci_idat[70:68])
      + conv_u2u_3_4(in_2_data_rsci_idat[70:68]);
  PECore_ProductSum_ccs_in_v1 #(.rscid(32'sd13),
  .width(32'sd128)) in_1_data_rsci (
      .dat(in_1_data_rsc_dat),
      .idat(in_1_data_rsci_idat)
    );
  PECore_ProductSum_ccs_in_v1 #(.rscid(32'sd14),
  .width(32'sd128)) in_2_data_rsci (
      .dat(in_2_data_rsc_dat),
      .idat(in_2_data_rsci_idat)
    );
  PECore_ProductSum_mgc_out_dreg_v2 #(.rscid(32'sd15),
  .width(32'sd32)) out_rsci (
      .d(nl_out_rsci_d[31:0]),
      .z(out_rsc_z)
    );
  PECore_ProductSum_ccs_in_v1 #(.rscid(32'sd148),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  PECore_ProductSum_mgc_shift_l_v5 #(.width_a(32'sd11),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd25)) for_10_adpfloat_mul_template_8U_3U_32U_lshift_rg (
      .a(nl_for_10_adpfloat_mul_template_8U_3U_32U_lshift_rg_a[10:0]),
      .s(nl_for_10_adpfloat_mul_template_8U_3U_32U_lshift_rg_s[3:0]),
      .z(for_10_adpfloat_mul_template_8U_3U_32U_lshift_itm)
    );
  PECore_ProductSum_mgc_shift_l_v5 #(.width_a(32'sd11),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd25)) for_11_adpfloat_mul_template_8U_3U_32U_lshift_rg (
      .a(nl_for_11_adpfloat_mul_template_8U_3U_32U_lshift_rg_a[10:0]),
      .s(nl_for_11_adpfloat_mul_template_8U_3U_32U_lshift_rg_s[3:0]),
      .z(for_11_adpfloat_mul_template_8U_3U_32U_lshift_itm)
    );
  PECore_ProductSum_mgc_shift_l_v5 #(.width_a(32'sd11),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd25)) for_12_adpfloat_mul_template_8U_3U_32U_lshift_rg (
      .a(nl_for_12_adpfloat_mul_template_8U_3U_32U_lshift_rg_a[10:0]),
      .s(nl_for_12_adpfloat_mul_template_8U_3U_32U_lshift_rg_s[3:0]),
      .z(for_12_adpfloat_mul_template_8U_3U_32U_lshift_itm)
    );
  PECore_ProductSum_mgc_shift_l_v5 #(.width_a(32'sd11),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd25)) for_13_adpfloat_mul_template_8U_3U_32U_lshift_rg (
      .a(nl_for_13_adpfloat_mul_template_8U_3U_32U_lshift_rg_a[10:0]),
      .s(nl_for_13_adpfloat_mul_template_8U_3U_32U_lshift_rg_s[3:0]),
      .z(for_13_adpfloat_mul_template_8U_3U_32U_lshift_itm)
    );
  PECore_ProductSum_mgc_shift_l_v5 #(.width_a(32'sd11),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd25)) for_14_adpfloat_mul_template_8U_3U_32U_lshift_rg (
      .a(nl_for_14_adpfloat_mul_template_8U_3U_32U_lshift_rg_a[10:0]),
      .s(nl_for_14_adpfloat_mul_template_8U_3U_32U_lshift_rg_s[3:0]),
      .z(for_14_adpfloat_mul_template_8U_3U_32U_lshift_itm)
    );
  PECore_ProductSum_mgc_shift_l_v5 #(.width_a(32'sd11),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd25)) for_15_adpfloat_mul_template_8U_3U_32U_lshift_rg (
      .a(nl_for_15_adpfloat_mul_template_8U_3U_32U_lshift_rg_a[10:0]),
      .s(nl_for_15_adpfloat_mul_template_8U_3U_32U_lshift_rg_s[3:0]),
      .z(for_15_adpfloat_mul_template_8U_3U_32U_lshift_itm)
    );
  PECore_ProductSum_mgc_shift_l_v5 #(.width_a(32'sd11),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd25)) for_16_adpfloat_mul_template_8U_3U_32U_lshift_rg (
      .a(nl_for_16_adpfloat_mul_template_8U_3U_32U_lshift_rg_a[10:0]),
      .s(nl_for_16_adpfloat_mul_template_8U_3U_32U_lshift_rg_s[3:0]),
      .z(for_16_adpfloat_mul_template_8U_3U_32U_lshift_itm)
    );
  PECore_ProductSum_mgc_shift_l_v5 #(.width_a(32'sd11),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd25)) for_1_adpfloat_mul_template_8U_3U_32U_lshift_rg (
      .a(nl_for_1_adpfloat_mul_template_8U_3U_32U_lshift_rg_a[10:0]),
      .s(nl_for_1_adpfloat_mul_template_8U_3U_32U_lshift_rg_s[3:0]),
      .z(for_1_adpfloat_mul_template_8U_3U_32U_lshift_itm)
    );
  PECore_ProductSum_mgc_shift_l_v5 #(.width_a(32'sd11),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd25)) for_2_adpfloat_mul_template_8U_3U_32U_lshift_rg (
      .a(nl_for_2_adpfloat_mul_template_8U_3U_32U_lshift_rg_a[10:0]),
      .s(nl_for_2_adpfloat_mul_template_8U_3U_32U_lshift_rg_s[3:0]),
      .z(for_2_adpfloat_mul_template_8U_3U_32U_lshift_itm)
    );
  PECore_ProductSum_mgc_shift_l_v5 #(.width_a(32'sd11),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd25)) for_3_adpfloat_mul_template_8U_3U_32U_lshift_rg (
      .a(nl_for_3_adpfloat_mul_template_8U_3U_32U_lshift_rg_a[10:0]),
      .s(nl_for_3_adpfloat_mul_template_8U_3U_32U_lshift_rg_s[3:0]),
      .z(for_3_adpfloat_mul_template_8U_3U_32U_lshift_itm)
    );
  PECore_ProductSum_mgc_shift_l_v5 #(.width_a(32'sd11),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd25)) for_4_adpfloat_mul_template_8U_3U_32U_lshift_rg (
      .a(nl_for_4_adpfloat_mul_template_8U_3U_32U_lshift_rg_a[10:0]),
      .s(nl_for_4_adpfloat_mul_template_8U_3U_32U_lshift_rg_s[3:0]),
      .z(for_4_adpfloat_mul_template_8U_3U_32U_lshift_itm)
    );
  PECore_ProductSum_mgc_shift_l_v5 #(.width_a(32'sd11),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd25)) for_5_adpfloat_mul_template_8U_3U_32U_lshift_rg (
      .a(nl_for_5_adpfloat_mul_template_8U_3U_32U_lshift_rg_a[10:0]),
      .s(nl_for_5_adpfloat_mul_template_8U_3U_32U_lshift_rg_s[3:0]),
      .z(for_5_adpfloat_mul_template_8U_3U_32U_lshift_itm)
    );
  PECore_ProductSum_mgc_shift_l_v5 #(.width_a(32'sd11),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd25)) for_6_adpfloat_mul_template_8U_3U_32U_lshift_rg (
      .a(nl_for_6_adpfloat_mul_template_8U_3U_32U_lshift_rg_a[10:0]),
      .s(nl_for_6_adpfloat_mul_template_8U_3U_32U_lshift_rg_s[3:0]),
      .z(for_6_adpfloat_mul_template_8U_3U_32U_lshift_itm)
    );
  PECore_ProductSum_mgc_shift_l_v5 #(.width_a(32'sd11),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd25)) for_7_adpfloat_mul_template_8U_3U_32U_lshift_rg (
      .a(nl_for_7_adpfloat_mul_template_8U_3U_32U_lshift_rg_a[10:0]),
      .s(nl_for_7_adpfloat_mul_template_8U_3U_32U_lshift_rg_s[3:0]),
      .z(for_7_adpfloat_mul_template_8U_3U_32U_lshift_itm)
    );
  PECore_ProductSum_mgc_shift_l_v5 #(.width_a(32'sd11),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd25)) for_8_adpfloat_mul_template_8U_3U_32U_lshift_rg (
      .a(nl_for_8_adpfloat_mul_template_8U_3U_32U_lshift_rg_a[10:0]),
      .s(nl_for_8_adpfloat_mul_template_8U_3U_32U_lshift_rg_s[3:0]),
      .z(for_8_adpfloat_mul_template_8U_3U_32U_lshift_itm)
    );
  PECore_ProductSum_mgc_shift_l_v5 #(.width_a(32'sd11),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd25)) for_9_adpfloat_mul_template_8U_3U_32U_lshift_rg (
      .a(nl_for_9_adpfloat_mul_template_8U_3U_32U_lshift_rg_a[10:0]),
      .s(nl_for_9_adpfloat_mul_template_8U_3U_32U_lshift_rg_s[3:0]),
      .z(for_9_adpfloat_mul_template_8U_3U_32U_lshift_itm)
    );
  PECore_ProductSum_ACC_16i25_1o29_6c39adcf8fa7ac08d026ec7c525fe9f9e6  U_ACC_16i25_1o29_c7aa682b5659f7f20224ec66be5b70f85d_rg
      (
      .I_1(for_10_adpfloat_mul_template_8U_3U_32U_lshift_itm),
      .I_2(for_11_adpfloat_mul_template_8U_3U_32U_lshift_itm),
      .I_3(for_12_adpfloat_mul_template_8U_3U_32U_lshift_itm),
      .I_4(for_13_adpfloat_mul_template_8U_3U_32U_lshift_itm),
      .I_5(for_14_adpfloat_mul_template_8U_3U_32U_lshift_itm),
      .I_6(for_15_adpfloat_mul_template_8U_3U_32U_lshift_itm),
      .I_7(for_16_adpfloat_mul_template_8U_3U_32U_lshift_itm),
      .I_8(for_1_adpfloat_mul_template_8U_3U_32U_lshift_itm),
      .I_9(for_2_adpfloat_mul_template_8U_3U_32U_lshift_itm),
      .I_10(for_3_adpfloat_mul_template_8U_3U_32U_lshift_itm),
      .I_11(for_4_adpfloat_mul_template_8U_3U_32U_lshift_itm),
      .I_12(for_5_adpfloat_mul_template_8U_3U_32U_lshift_itm),
      .I_13(for_6_adpfloat_mul_template_8U_3U_32U_lshift_itm),
      .I_14(for_7_adpfloat_mul_template_8U_3U_32U_lshift_itm),
      .I_15(for_8_adpfloat_mul_template_8U_3U_32U_lshift_itm),
      .I_16(for_9_adpfloat_mul_template_8U_3U_32U_lshift_itm),
      .O_1(ACC_16i25_1o29_c7aa682b5659f7f20224ec66be5b70f85d_1)
    );
  assign nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_1_sva_1 = ({1'b1 ,
      (~ adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_1_sva_1)}) + 11'b00000000001;
  assign adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_1_sva_1 = nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_1_sva_1[10:0];
  assign for_1_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      = (in_1_data_rsci_idat[6:0]!=7'b0000000);
  assign for_1_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      = (in_2_data_rsci_idat[6:0]!=7'b0000000);
  assign adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_1_sva_1 = conv_u2u_10_10(({for_1_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      , (in_1_data_rsci_idat[3:0])}) * ({for_1_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      , (in_2_data_rsci_idat[3:0])}));
  assign nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_2_sva_1 = ({1'b1 ,
      (~ adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_2_sva_1)}) + 11'b00000000001;
  assign adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_2_sva_1 = nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_2_sva_1[10:0];
  assign for_2_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      = (in_1_data_rsci_idat[14:8]!=7'b0000000);
  assign for_2_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      = (in_2_data_rsci_idat[14:8]!=7'b0000000);
  assign adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_2_sva_1 = conv_u2u_10_10(({for_2_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      , (in_1_data_rsci_idat[11:8])}) * ({for_2_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      , (in_2_data_rsci_idat[11:8])}));
  assign nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_3_sva_1 = ({1'b1 ,
      (~ adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_3_sva_1)}) + 11'b00000000001;
  assign adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_3_sva_1 = nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_3_sva_1[10:0];
  assign for_3_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      = (in_1_data_rsci_idat[22:16]!=7'b0000000);
  assign for_3_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      = (in_2_data_rsci_idat[22:16]!=7'b0000000);
  assign adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_3_sva_1 = conv_u2u_10_10(({for_3_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      , (in_1_data_rsci_idat[19:16])}) * ({for_3_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      , (in_2_data_rsci_idat[19:16])}));
  assign nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_4_sva_1 = ({1'b1 ,
      (~ adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_4_sva_1)}) + 11'b00000000001;
  assign adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_4_sva_1 = nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_4_sva_1[10:0];
  assign for_4_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      = (in_1_data_rsci_idat[30:24]!=7'b0000000);
  assign for_4_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      = (in_2_data_rsci_idat[30:24]!=7'b0000000);
  assign adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_4_sva_1 = conv_u2u_10_10(({for_4_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      , (in_1_data_rsci_idat[27:24])}) * ({for_4_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      , (in_2_data_rsci_idat[27:24])}));
  assign nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_5_sva_1 = ({1'b1 ,
      (~ adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_5_sva_1)}) + 11'b00000000001;
  assign adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_5_sva_1 = nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_5_sva_1[10:0];
  assign for_5_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      = (in_1_data_rsci_idat[38:32]!=7'b0000000);
  assign for_5_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      = (in_2_data_rsci_idat[38:32]!=7'b0000000);
  assign adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_5_sva_1 = conv_u2u_10_10(({for_5_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      , (in_1_data_rsci_idat[35:32])}) * ({for_5_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      , (in_2_data_rsci_idat[35:32])}));
  assign nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_6_sva_1 = ({1'b1 ,
      (~ adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_6_sva_1)}) + 11'b00000000001;
  assign adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_6_sva_1 = nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_6_sva_1[10:0];
  assign for_6_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      = (in_1_data_rsci_idat[46:40]!=7'b0000000);
  assign for_6_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      = (in_2_data_rsci_idat[46:40]!=7'b0000000);
  assign adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_6_sva_1 = conv_u2u_10_10(({for_6_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      , (in_1_data_rsci_idat[43:40])}) * ({for_6_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      , (in_2_data_rsci_idat[43:40])}));
  assign nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_7_sva_1 = ({1'b1 ,
      (~ adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_7_sva_1)}) + 11'b00000000001;
  assign adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_7_sva_1 = nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_7_sva_1[10:0];
  assign for_7_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      = (in_1_data_rsci_idat[54:48]!=7'b0000000);
  assign for_7_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      = (in_2_data_rsci_idat[54:48]!=7'b0000000);
  assign adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_7_sva_1 = conv_u2u_10_10(({for_7_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      , (in_1_data_rsci_idat[51:48])}) * ({for_7_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      , (in_2_data_rsci_idat[51:48])}));
  assign nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_8_sva_1 = ({1'b1 ,
      (~ adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_8_sva_1)}) + 11'b00000000001;
  assign adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_8_sva_1 = nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_8_sva_1[10:0];
  assign for_8_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      = (in_1_data_rsci_idat[62:56]!=7'b0000000);
  assign for_8_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      = (in_2_data_rsci_idat[62:56]!=7'b0000000);
  assign adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_8_sva_1 = conv_u2u_10_10(({for_8_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      , (in_1_data_rsci_idat[59:56])}) * ({for_8_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      , (in_2_data_rsci_idat[59:56])}));
  assign nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_9_sva_1 = ({1'b1 ,
      (~ adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_9_sva_1)}) + 11'b00000000001;
  assign adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_9_sva_1 = nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_9_sva_1[10:0];
  assign for_9_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      = (in_1_data_rsci_idat[70:64]!=7'b0000000);
  assign for_9_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      = (in_2_data_rsci_idat[70:64]!=7'b0000000);
  assign adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_9_sva_1 = conv_u2u_10_10(({for_9_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      , (in_1_data_rsci_idat[67:64])}) * ({for_9_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      , (in_2_data_rsci_idat[67:64])}));
  assign nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_10_sva_1 = ({1'b1 ,
      (~ adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_10_sva_1)}) + 11'b00000000001;
  assign adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_10_sva_1 = nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_10_sva_1[10:0];
  assign for_10_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      = (in_1_data_rsci_idat[78:72]!=7'b0000000);
  assign for_10_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      = (in_2_data_rsci_idat[78:72]!=7'b0000000);
  assign adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_10_sva_1 = conv_u2u_10_10(({for_10_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      , (in_1_data_rsci_idat[75:72])}) * ({for_10_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      , (in_2_data_rsci_idat[75:72])}));
  assign nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_11_sva_1 = ({1'b1 ,
      (~ adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_11_sva_1)}) + 11'b00000000001;
  assign adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_11_sva_1 = nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_11_sva_1[10:0];
  assign for_11_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      = (in_1_data_rsci_idat[86:80]!=7'b0000000);
  assign for_11_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      = (in_2_data_rsci_idat[86:80]!=7'b0000000);
  assign adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_11_sva_1 = conv_u2u_10_10(({for_11_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      , (in_1_data_rsci_idat[83:80])}) * ({for_11_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      , (in_2_data_rsci_idat[83:80])}));
  assign nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_12_sva_1 = ({1'b1 ,
      (~ adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_12_sva_1)}) + 11'b00000000001;
  assign adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_12_sva_1 = nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_12_sva_1[10:0];
  assign for_12_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      = (in_1_data_rsci_idat[94:88]!=7'b0000000);
  assign for_12_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      = (in_2_data_rsci_idat[94:88]!=7'b0000000);
  assign adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_12_sva_1 = conv_u2u_10_10(({for_12_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      , (in_1_data_rsci_idat[91:88])}) * ({for_12_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      , (in_2_data_rsci_idat[91:88])}));
  assign nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_13_sva_1 = ({1'b1 ,
      (~ adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_13_sva_1)}) + 11'b00000000001;
  assign adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_13_sva_1 = nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_13_sva_1[10:0];
  assign for_13_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      = (in_1_data_rsci_idat[102:96]!=7'b0000000);
  assign for_13_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      = (in_2_data_rsci_idat[102:96]!=7'b0000000);
  assign adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_13_sva_1 = conv_u2u_10_10(({for_13_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      , (in_1_data_rsci_idat[99:96])}) * ({for_13_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      , (in_2_data_rsci_idat[99:96])}));
  assign nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_14_sva_1 = ({1'b1 ,
      (~ adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_14_sva_1)}) + 11'b00000000001;
  assign adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_14_sva_1 = nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_14_sva_1[10:0];
  assign for_14_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      = (in_1_data_rsci_idat[110:104]!=7'b0000000);
  assign for_14_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      = (in_2_data_rsci_idat[110:104]!=7'b0000000);
  assign adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_14_sva_1 = conv_u2u_10_10(({for_14_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      , (in_1_data_rsci_idat[107:104])}) * ({for_14_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      , (in_2_data_rsci_idat[107:104])}));
  assign nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_15_sva_1 = ({1'b1 ,
      (~ adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_15_sva_1)}) + 11'b00000000001;
  assign adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_15_sva_1 = nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_15_sva_1[10:0];
  assign for_15_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      = (in_1_data_rsci_idat[118:112]!=7'b0000000);
  assign for_15_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      = (in_2_data_rsci_idat[118:112]!=7'b0000000);
  assign adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_15_sva_1 = conv_u2u_10_10(({for_15_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      , (in_1_data_rsci_idat[115:112])}) * ({for_15_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      , (in_2_data_rsci_idat[115:112])}));
  assign nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_sva_1 = ({1'b1 , (~
      adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_sva_1)}) + 11'b00000000001;
  assign adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_sva_1 = nl_adpfloat_mul_template_8U_3U_32U_if_2_ac_int_cctor_sva_1[10:0];
  assign for_16_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      = (in_1_data_rsci_idat[126:120]!=7'b0000000);
  assign for_16_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      = (in_2_data_rsci_idat[126:120]!=7'b0000000);
  assign adpfloat_mul_template_8U_3U_32U_ac_int_cctor_2_9_0_sva_1 = conv_u2u_10_10(({for_16_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_in_a_is_zero_out_in_a_is_zero_if_or_nl
      , (in_1_data_rsci_idat[123:120])}) * ({for_16_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_1_in_b_is_zero_out_in_b_is_zero_if_or_nl
      , (in_2_data_rsci_idat[123:120])}));
  assign for_10_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1
      = (in_1_data_rsci_idat[79]) ^ (in_2_data_rsci_idat[79]);
  assign for_11_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1
      = (in_1_data_rsci_idat[87]) ^ (in_2_data_rsci_idat[87]);
  assign for_12_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1
      = (in_1_data_rsci_idat[95]) ^ (in_2_data_rsci_idat[95]);
  assign for_13_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1
      = (in_1_data_rsci_idat[103]) ^ (in_2_data_rsci_idat[103]);
  assign for_14_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1
      = (in_1_data_rsci_idat[111]) ^ (in_2_data_rsci_idat[111]);
  assign for_15_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1
      = (in_1_data_rsci_idat[119]) ^ (in_2_data_rsci_idat[119]);
  assign for_16_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1
      = (in_1_data_rsci_idat[127]) ^ (in_2_data_rsci_idat[127]);
  assign for_1_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1
      = (in_1_data_rsci_idat[7]) ^ (in_2_data_rsci_idat[7]);
  assign for_2_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1
      = (in_1_data_rsci_idat[15]) ^ (in_2_data_rsci_idat[15]);
  assign for_3_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1
      = (in_1_data_rsci_idat[23]) ^ (in_2_data_rsci_idat[23]);
  assign for_4_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1
      = (in_1_data_rsci_idat[31]) ^ (in_2_data_rsci_idat[31]);
  assign for_5_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1
      = (in_1_data_rsci_idat[39]) ^ (in_2_data_rsci_idat[39]);
  assign for_6_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1
      = (in_1_data_rsci_idat[47]) ^ (in_2_data_rsci_idat[47]);
  assign for_7_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1
      = (in_1_data_rsci_idat[55]) ^ (in_2_data_rsci_idat[55]);
  assign for_8_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1
      = (in_1_data_rsci_idat[63]) ^ (in_2_data_rsci_idat[63]);
  assign for_9_adpfloat_mul_template_8U_3U_32U_adpfloat_mul_template_8U_3U_32U_if_2_xor_svs_1
      = (in_1_data_rsci_idat[71]) ^ (in_2_data_rsci_idat[71]);
  always @(posedge ccs_ccore_clk) begin
    if ( ~ ccs_ccore_arst ) begin
      out_rsci_d_28_0 <= 29'b00000000000000000000000000000;
    end
    else if ( ccs_ccore_en & ccs_ccore_start_rsci_idat ) begin
      out_rsci_d_28_0 <= ACC_16i25_1o29_c7aa682b5659f7f20224ec66be5b70f85d_1;
    end
  end

  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input  sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_10_10 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_10 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ProductSum
// ------------------------------------------------------------------


module PECore_ProductSum (
  in_1_data_rsc_dat, in_2_data_rsc_dat, out_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_arst, ccs_ccore_en
);
  input [127:0] in_1_data_rsc_dat;
  input [127:0] in_2_data_rsc_dat;
  output [31:0] out_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations
  PECore_ProductSum_ProductSum_core ProductSum_core_inst (
      .in_1_data_rsc_dat(in_1_data_rsc_dat),
      .in_2_data_rsc_dat(in_2_data_rsc_dat),
      .out_rsc_z(out_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ./PECore_mgc_muladd1_beh.v 
//muladd1
module PECore_mgc_muladd1(a,b,c,cst,d,z);
  // operation is z = a * (b + d) + c + cst
  parameter width_a = 0;
  parameter signd_a = 0;
  parameter width_b = 0;
  parameter signd_b = 0;
  parameter width_c = 0;
  parameter signd_c = 0;
  parameter width_cst = 0;
  parameter signd_cst = 0;
  parameter width_d = 0;
  parameter signd_d = 0;
  parameter width_z = 0;
  parameter add_axb = 1;
  parameter add_c = 1;
  parameter add_d = 1;
  parameter use_const = 1;
  input  [width_a-1:0] a;
  input  [width_b-1:0] b;
  input  [width_c-1:0] c;
  input  [width_cst-1:0] cst;
  input  [width_d-1:0] d;
  output [width_z-1:0] z;

  reg [width_a-signd_a:0] aa;
  reg [width_b-signd_b:0] bb;
  reg [width_c-signd_c:0] cc;
  reg [width_d-signd_d:0] dd;
  reg [width_cst-signd_cst:0] cstin;

  localparam width_bd = (width_d) ? 1+ ((width_b-signd_b>width_d-signd_d) ? width_b - signd_b
                                                                          : width_d - signd_d)
                                  : width_b - signd_b;
  reg [width_bd:0] bd;

  // make all inputs signed
  always @(*) aa = signd_a ? a : {1'b0, a};
  always @(*) bb = signd_b ? b : {1'b0, b};
  generate if (width_c) begin
    always @(*) cc = signd_c ? c : {1'b0, c};
  end endgenerate
  generate if (width_d) begin
    always @(*) dd = signd_d ? d : {1'b0, d};
  end endgenerate
  always @(*) cstin = signd_cst ? cst : {1'b0, cst};

  // perform pre-adder
  generate
    if (width_d) begin
      if (add_d) begin always @(*)  bd = $signed(bb) + $signed(dd); end
      else       begin always @(*)  bd = $signed(bb) - $signed(dd); end
    end else     begin always @(*)  bd = $signed(bb); end
  endgenerate

  // perform muladd1
  wire [width_z-1:0]  zz;

  generate
    if (use_const) begin
      if ( add_axb &&  add_c && width_c) begin assign zz = ($signed(aa) * $signed(bd)) + $signed(cc) + $signed(cstin); end else
      if ( add_axb && !add_c && width_c) begin assign zz = ($signed(aa) * $signed(bd)) - $signed(cc) + $signed(cstin); end else
      if (!add_axb &&  add_c && width_c) begin assign zz = $signed(cc) - ($signed(aa) * $signed(bd)) + $signed(cstin); end else
      if (!add_axb && !add_c && width_c) begin assign zz = $signed(cstin) - ($signed(aa) * $signed(bd)) - $signed(cc); end else
      if ( add_axb )                     begin assign zz = ($signed(aa) * $signed(bd)) + $signed(cstin); end else
                                         begin assign zz = $signed(cstin) - ($signed(aa) * $signed(bd)); end
    end  else begin
      if ( add_axb &&  add_c && width_c) begin assign zz = ($signed(aa) * $signed(bd)) + $signed(cc); end else
      if ( add_axb && !add_c && width_c) begin assign zz = ($signed(aa) * $signed(bd)) - $signed(cc); end else
      if (!add_axb &&  add_c && width_c) begin assign zz = $signed(cc) - ($signed(aa) * $signed(bd)); end else
      if (!add_axb && !add_c && width_c) begin assign zz = -($signed(aa) * $signed(bd)) - $signed(cc); end else
      if ( add_axb )                     begin assign zz = ($signed(aa) * $signed(bd)); end else
                                         begin assign zz = -($signed(aa) * $signed(bd)); end
    end
  endgenerate

  // adjust output
  assign z = zz;
endmodule // mgc_muladd1

//------> ./PECore_mgc_shift_l_beh_v5.v 
module PECore_mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./PECore_mgc_shift_r_beh_v5.v 
module PECore_mgc_shift_r_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SGNED
       assign z = fshr_u(a,s,a[width_a-1]);
     end
     else
     begin: UNSGNED
       assign z = fshr_u(a,s,1'b0);
     end
   endgenerate

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

endmodule

//------> ./PECore_mgc_shift_bl_beh_v5.v 
module PECore_mgc_shift_bl_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate if ( signd_a )
   begin: SGNED
     assign z = fshl_s(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
     assign z = fshl_s(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift left - signed shift argument
   function [width_z-1:0] fshl_s;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      reg [width_a:0] sbit_arg1;
      begin
        // Ignoring the possibility that arg2[width_s-1] could be X
        // because of customer complaints regarding X'es in simulation results
        if ( arg2[width_s-1] == 1'b0 )
        begin
          sbit_arg1[width_a:0] = {(width_a+1){1'b0}};
          fshl_s = fshl_u(arg1, arg2, sbit);
        end
        else
        begin
          sbit_arg1[width_a] = sbit;
          sbit_arg1[width_a-1:0] = arg1;
          fshl_s = fshr_u(sbit_arg1[width_a:1], ~arg2, sbit);
        end
      end
   endfunction

endmodule

//------> /usr/licensed/MentorGraphics2021/Catapult_Synthesis_10.6a/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Memory Type:            BLOCK
// Operating Mode:         Simple Dual Port (2-Port)
// Clock Mode:             Single Clock
// 
// RTL Code RW Resolution: RBW
// Catapult RW Resolution: RBW
// 
// HDL Work Library:       Xilinx_RAMS_lib
// Component Name:         BLOCK_1R1W_RBW
// Latency = 1:            RAM with no registers on inputs or outputs
//         = 2:            adds embedded register on RAM output
//         = 3:            adds fabric registers to non-clock input RAM pins
//         = 4:            adds fabric register to output (driven by embedded register from latency=2)

module BLOCK_1R1W_RBW #(
  parameter addr_width = 8 ,
  parameter data_width = 7 ,
  parameter depth = 256 ,
  parameter latency = 1 
  
)( clk,clken,d,q,radr,wadr,we);

  input  clk;
  input  clken;
  input [data_width-1:0] d;
  output [data_width-1:0] q;
  input [addr_width-1:0] radr;
  input [addr_width-1:0] wadr;
  input  we;
  
  (* ram_style = "block" *)
  reg [data_width-1:0] mem [depth-1:0];// synthesis syn_ramstyle="block"
  
  reg [data_width-1:0] ramq;
  
  // Port Map
  // readA :: CLOCK clk ENABLE clken DATA_OUT q ADDRESS radr
  // writeA :: CLOCK clk ENABLE clken DATA_IN d ADDRESS wadr WRITE_ENABLE we

  generate
    // Register all non-clock inputs (latency < 3)
    if (latency > 2 ) begin
      reg [addr_width-1:0] radr_reg;
      reg [data_width-1:0] d_reg;
      reg [addr_width-1:0] wadr_reg;
      reg we_reg;
      
      always @(posedge clk) begin
        if (clken) begin
          radr_reg <= radr;
        end
      end
      always @(posedge clk) begin
        if (clken) begin
          d_reg <= d;
          wadr_reg <= wadr;
          we_reg <= we;
        end
      end
      
    // Access memory with registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr_reg];
            if (we_reg) begin
              mem[wadr_reg] <= d_reg;
            end
        end
      end
      
    end // END register inputs

    else begin
    // latency = 1||2: Access memory with non-registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr];
            if (we) begin
              mem[wadr] <= d;
            end
        end
      end
      
    end
  endgenerate //END input port generate 

  generate
    // latency=1: sequential RAM outputs drive module outputs
    if (latency == 1) begin
      assign q = ramq;
      
    end

    else if (latency == 2 || latency == 3) begin
    // latency=2: sequential (RAM output => tmp register => module output)
      reg [data_width-1:0] tmpq;
      
      always @(posedge clk) begin
        if (clken) begin
          tmpq <= ramq;
        end
      end
      
      assign q = tmpq;
      
    end
    else if (latency == 4) begin
    // latency=4: (RAM => tmp1 register => tmp2 fabric register => module output)
      reg [data_width-1:0] tmp1q;
      
      reg [data_width-1:0] tmp2q;
      
      always @(posedge clk) begin
        if (clken) begin
          tmp1q <= ramq;
        end
      end
      
      always @(posedge clk) begin
        if (clken) begin
          tmp2q <= tmp1q;
        end
      end
      
      assign q = tmp2q;
      
    end
    else begin
      //Add error check if latency > 4 or add N-pipeline regs
    end
  endgenerate //END output port generate

endmodule

//------> ./PECore.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.6a/933210 Production Release
//  HLS Date:       Mon Apr 12 07:56:29 PDT 2021
// 
//  Generated date: Mon Apr  4 22:46:53 2022
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_125_8_128_256_256_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_125_8_128_256_256_128_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output [7:0] radr;
  output we;
  output [127:0] d;
  output [7:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [7:0] radr_d;
  input [7:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_123_12_128_4096_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_123_12_128_4096_4096_128_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_122_12_128_4096_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_122_12_128_4096_4096_128_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_121_12_128_4096_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_121_12_128_4096_4096_128_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_120_12_128_4096_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_120_12_128_4096_4096_128_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_119_12_128_4096_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_119_12_128_4096_4096_128_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_118_12_128_4096_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_118_12_128_4096_4096_128_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_117_12_128_4096_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_117_12_128_4096_4096_128_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_116_12_128_4096_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_116_12_128_4096_4096_128_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_115_12_128_4096_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_115_12_128_4096_4096_128_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_114_12_128_4096_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_114_12_128_4096_4096_128_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_113_12_128_4096_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_113_12_128_4096_4096_128_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_112_12_128_4096_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_112_12_128_4096_4096_128_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_111_12_128_4096_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_111_12_128_4096_4096_128_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_110_12_128_4096_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_110_12_128_4096_4096_128_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_109_12_128_4096_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_109_12_128_4096_4096_128_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_108_12_128_4096_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_108_12_128_4096_4096_128_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_PECoreRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_PECoreRun_fsm (
  clk, rst, PECoreRun_wen, fsm_output
);
  input clk;
  input rst;
  input PECoreRun_wen;
  output [4:0] fsm_output;
  reg [4:0] fsm_output;


  // FSM State Type Declaration for PECore_PECore_PECoreRun_PECoreRun_fsm_1
  parameter
    PECoreRun_rlp_C_0 = 3'd0,
    while_C_0 = 3'd1,
    while_C_1 = 3'd2,
    while_C_2 = 3'd3,
    while_C_3 = 3'd4;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : PECore_PECore_PECoreRun_PECoreRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 5'b00010;
        state_var_NS = while_C_1;
      end
      while_C_1 : begin
        fsm_output = 5'b00100;
        state_var_NS = while_C_2;
      end
      while_C_2 : begin
        fsm_output = 5'b01000;
        state_var_NS = while_C_3;
      end
      while_C_3 : begin
        fsm_output = 5'b10000;
        state_var_NS = while_C_0;
      end
      // PECoreRun_rlp_C_0
      default : begin
        fsm_output = 5'b00001;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk ) begin
    if ( ~ rst ) begin
      state_var <= PECoreRun_rlp_C_0;
    end
    else if ( PECoreRun_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_staller
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_staller (
  clk, rst, PECoreRun_wen, PECoreRun_wten, act_port_Push_mioi_wen_comp, rva_out_Push_mioi_wen_comp
);
  input clk;
  input rst;
  output PECoreRun_wen;
  output PECoreRun_wten;
  reg PECoreRun_wten;
  input act_port_Push_mioi_wen_comp;
  input rva_out_Push_mioi_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign PECoreRun_wen = act_port_Push_mioi_wen_comp & rva_out_Push_mioi_wen_comp;
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      PECoreRun_wten <= 1'b0;
    end
    else begin
      PECoreRun_wten <= ~ PECoreRun_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp (
  clk, rst, start_PopNB_mioi_idat_mxwt, start_PopNB_mioi_ivld_mxwt, start_PopNB_mioi_biwt,
      start_PopNB_mioi_bdwt, start_PopNB_mioi_idat, start_PopNB_mioi_ivld
);
  input clk;
  input rst;
  output start_PopNB_mioi_idat_mxwt;
  output start_PopNB_mioi_ivld_mxwt;
  input start_PopNB_mioi_biwt;
  input start_PopNB_mioi_bdwt;
  input start_PopNB_mioi_idat;
  input start_PopNB_mioi_ivld;


  // Interconnect Declarations
  reg start_PopNB_mioi_bcwt;
  reg start_PopNB_mioi_idat_bfwt;
  reg start_PopNB_mioi_ivld_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_idat_mxwt = MUX_s_1_2_2(start_PopNB_mioi_idat, start_PopNB_mioi_idat_bfwt,
      start_PopNB_mioi_bcwt);
  assign start_PopNB_mioi_ivld_mxwt = MUX_s_1_2_2(start_PopNB_mioi_ivld, start_PopNB_mioi_ivld_bfwt,
      start_PopNB_mioi_bcwt);
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      start_PopNB_mioi_bcwt <= ~((~(start_PopNB_mioi_bcwt | start_PopNB_mioi_biwt))
          | start_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_idat_bfwt <= 1'b0;
      start_PopNB_mioi_ivld_bfwt <= 1'b0;
    end
    else if ( start_PopNB_mioi_biwt ) begin
      start_PopNB_mioi_idat_bfwt <= start_PopNB_mioi_idat;
      start_PopNB_mioi_ivld_bfwt <= start_PopNB_mioi_ivld;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl (
  PECoreRun_wen, PECoreRun_wten, start_PopNB_mioi_oswt, start_PopNB_mioi_biwt, start_PopNB_mioi_bdwt
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_biwt;
  output start_PopNB_mioi_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_bdwt = start_PopNB_mioi_oswt & PECoreRun_wen;
  assign start_PopNB_mioi_biwt = (~ PECoreRun_wten) & start_PopNB_mioi_oswt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp (
  clk, rst, rva_out_Push_mioi_oswt, rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_biwt,
      rva_out_Push_mioi_bdwt, rva_out_Push_mioi_bcwt
);
  input clk;
  input rst;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input rva_out_Push_mioi_biwt;
  input rva_out_Push_mioi_bdwt;
  output rva_out_Push_mioi_bcwt;
  reg rva_out_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_wen_comp = (~ rva_out_Push_mioi_oswt) | rva_out_Push_mioi_biwt
      | rva_out_Push_mioi_bcwt;
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_out_Push_mioi_bcwt <= ~((~(rva_out_Push_mioi_bcwt | rva_out_Push_mioi_biwt))
          | rva_out_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl (
  PECoreRun_wen, rva_out_Push_mioi_oswt, rva_out_Push_mioi_biwt, rva_out_Push_mioi_bdwt,
      rva_out_Push_mioi_bcwt, rva_out_Push_mioi_ivld_PECoreRun_sct, rva_out_Push_mioi_irdy
);
  input PECoreRun_wen;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_biwt;
  output rva_out_Push_mioi_bdwt;
  input rva_out_Push_mioi_bcwt;
  output rva_out_Push_mioi_ivld_PECoreRun_sct;
  input rva_out_Push_mioi_irdy;


  // Interconnect Declarations
  wire rva_out_Push_mioi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_bdwt = rva_out_Push_mioi_oswt & PECoreRun_wen;
  assign rva_out_Push_mioi_biwt = rva_out_Push_mioi_ogwt & rva_out_Push_mioi_irdy;
  assign rva_out_Push_mioi_ogwt = rva_out_Push_mioi_oswt & (~ rva_out_Push_mioi_bcwt);
  assign rva_out_Push_mioi_ivld_PECoreRun_sct = rva_out_Push_mioi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp (
  clk, rst, act_port_Push_mioi_oswt, act_port_Push_mioi_wen_comp, act_port_Push_mioi_biwt,
      act_port_Push_mioi_bdwt, act_port_Push_mioi_bcwt
);
  input clk;
  input rst;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_wen_comp;
  input act_port_Push_mioi_biwt;
  input act_port_Push_mioi_bdwt;
  output act_port_Push_mioi_bcwt;
  reg act_port_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign act_port_Push_mioi_wen_comp = (~ act_port_Push_mioi_oswt) | act_port_Push_mioi_biwt
      | act_port_Push_mioi_bcwt;
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      act_port_Push_mioi_bcwt <= ~((~(act_port_Push_mioi_bcwt | act_port_Push_mioi_biwt))
          | act_port_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl (
  PECoreRun_wen, act_port_Push_mioi_oswt, act_port_Push_mioi_biwt, act_port_Push_mioi_bdwt,
      act_port_Push_mioi_bcwt, act_port_Push_mioi_ivld_PECoreRun_sct, act_port_Push_mioi_irdy
);
  input PECoreRun_wen;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_biwt;
  output act_port_Push_mioi_bdwt;
  input act_port_Push_mioi_bcwt;
  output act_port_Push_mioi_ivld_PECoreRun_sct;
  input act_port_Push_mioi_irdy;


  // Interconnect Declarations
  wire act_port_Push_mioi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign act_port_Push_mioi_bdwt = act_port_Push_mioi_oswt & PECoreRun_wen;
  assign act_port_Push_mioi_biwt = act_port_Push_mioi_ogwt & act_port_Push_mioi_irdy;
  assign act_port_Push_mioi_ogwt = act_port_Push_mioi_oswt & (~ act_port_Push_mioi_bcwt);
  assign act_port_Push_mioi_ivld_PECoreRun_sct = act_port_Push_mioi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp (
  clk, rst, rva_in_PopNB_mioi_idat_mxwt, rva_in_PopNB_mioi_ivld_mxwt, rva_in_PopNB_mioi_biwt,
      rva_in_PopNB_mioi_bdwt, rva_in_PopNB_mioi_idat, rva_in_PopNB_mioi_ivld
);
  input clk;
  input rst;
  output [168:0] rva_in_PopNB_mioi_idat_mxwt;
  output rva_in_PopNB_mioi_ivld_mxwt;
  input rva_in_PopNB_mioi_biwt;
  input rva_in_PopNB_mioi_bdwt;
  input [168:0] rva_in_PopNB_mioi_idat;
  input rva_in_PopNB_mioi_ivld;


  // Interconnect Declarations
  reg rva_in_PopNB_mioi_bcwt;
  reg [168:0] rva_in_PopNB_mioi_idat_bfwt;
  reg rva_in_PopNB_mioi_ivld_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_idat_mxwt = MUX_v_169_2_2(rva_in_PopNB_mioi_idat, rva_in_PopNB_mioi_idat_bfwt,
      rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_ivld_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_ivld, rva_in_PopNB_mioi_ivld_bfwt,
      rva_in_PopNB_mioi_bcwt);
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_in_PopNB_mioi_bcwt <= ~((~(rva_in_PopNB_mioi_bcwt | rva_in_PopNB_mioi_biwt))
          | rva_in_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_idat_bfwt <= 169'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      rva_in_PopNB_mioi_ivld_bfwt <= 1'b0;
    end
    else if ( rva_in_PopNB_mioi_biwt ) begin
      rva_in_PopNB_mioi_idat_bfwt <= rva_in_PopNB_mioi_idat;
      rva_in_PopNB_mioi_ivld_bfwt <= rva_in_PopNB_mioi_ivld;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [168:0] MUX_v_169_2_2;
    input [168:0] input_0;
    input [168:0] input_1;
    input  sel;
    reg [168:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_169_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl (
  PECoreRun_wen, PECoreRun_wten, rva_in_PopNB_mioi_oswt, rva_in_PopNB_mioi_biwt,
      rva_in_PopNB_mioi_bdwt
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output rva_in_PopNB_mioi_biwt;
  output rva_in_PopNB_mioi_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_bdwt = rva_in_PopNB_mioi_oswt & PECoreRun_wen;
  assign rva_in_PopNB_mioi_biwt = (~ PECoreRun_wten) & rva_in_PopNB_mioi_oswt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_wait_dp (
  weight_mem_banks_bank_array_impl_data0_rsci_clken_d, weight_mem_banks_bank_array_impl_data1_rsci_clken_d,
      weight_mem_banks_bank_array_impl_data2_rsci_clken_d, weight_mem_banks_bank_array_impl_data3_rsci_clken_d,
      weight_mem_banks_bank_array_impl_data4_rsci_clken_d, weight_mem_banks_bank_array_impl_data5_rsci_clken_d,
      weight_mem_banks_bank_array_impl_data6_rsci_clken_d, weight_mem_banks_bank_array_impl_data7_rsci_clken_d,
      weight_mem_banks_bank_array_impl_data8_rsci_clken_d, weight_mem_banks_bank_array_impl_data9_rsci_clken_d,
      weight_mem_banks_bank_array_impl_data10_rsci_clken_d, weight_mem_banks_bank_array_impl_data11_rsci_clken_d,
      weight_mem_banks_bank_array_impl_data12_rsci_clken_d, weight_mem_banks_bank_array_impl_data13_rsci_clken_d,
      weight_mem_banks_bank_array_impl_data14_rsci_clken_d, weight_mem_banks_bank_array_impl_data15_rsci_clken_d,
      input_mem_banks_bank_array_impl_data0_rsci_clken_d, PECoreRun_wen, weight_mem_banks_bank_array_impl_data0_rsci_cgo,
      weight_mem_banks_bank_array_impl_data0_rsci_cgo_ir_unreg, weight_mem_banks_bank_array_impl_data1_rsci_cgo,
      weight_mem_banks_bank_array_impl_data1_rsci_cgo_ir_unreg, weight_mem_banks_bank_array_impl_data2_rsci_cgo,
      weight_mem_banks_bank_array_impl_data2_rsci_cgo_ir_unreg, weight_mem_banks_bank_array_impl_data3_rsci_cgo,
      weight_mem_banks_bank_array_impl_data3_rsci_cgo_ir_unreg, weight_mem_banks_bank_array_impl_data4_rsci_cgo,
      weight_mem_banks_bank_array_impl_data4_rsci_cgo_ir_unreg, weight_mem_banks_bank_array_impl_data5_rsci_cgo,
      weight_mem_banks_bank_array_impl_data5_rsci_cgo_ir_unreg, weight_mem_banks_bank_array_impl_data6_rsci_cgo,
      weight_mem_banks_bank_array_impl_data6_rsci_cgo_ir_unreg, weight_mem_banks_bank_array_impl_data7_rsci_cgo,
      weight_mem_banks_bank_array_impl_data7_rsci_cgo_ir_unreg, weight_mem_banks_bank_array_impl_data8_rsci_cgo,
      weight_mem_banks_bank_array_impl_data8_rsci_cgo_ir_unreg, weight_mem_banks_bank_array_impl_data9_rsci_cgo,
      weight_mem_banks_bank_array_impl_data9_rsci_cgo_ir_unreg, weight_mem_banks_bank_array_impl_data10_rsci_cgo,
      weight_mem_banks_bank_array_impl_data10_rsci_cgo_ir_unreg, weight_mem_banks_bank_array_impl_data11_rsci_cgo,
      weight_mem_banks_bank_array_impl_data11_rsci_cgo_ir_unreg, weight_mem_banks_bank_array_impl_data12_rsci_cgo,
      weight_mem_banks_bank_array_impl_data12_rsci_cgo_ir_unreg, weight_mem_banks_bank_array_impl_data13_rsci_cgo,
      weight_mem_banks_bank_array_impl_data13_rsci_cgo_ir_unreg, weight_mem_banks_bank_array_impl_data14_rsci_cgo,
      weight_mem_banks_bank_array_impl_data14_rsci_cgo_ir_unreg, weight_mem_banks_bank_array_impl_data15_rsci_cgo,
      weight_mem_banks_bank_array_impl_data15_rsci_cgo_ir_unreg, input_mem_banks_bank_array_impl_data0_rsci_cgo,
      input_mem_banks_bank_array_impl_data0_rsci_cgo_ir_unreg, Datapath_for_1_ProductSum_cmp_cgo,
      Datapath_for_1_ProductSum_cmp_cgo_ir_unreg, Datapath_for_1_ProductSum_cmp_ccs_ccore_en
);
  output weight_mem_banks_bank_array_impl_data0_rsci_clken_d;
  output weight_mem_banks_bank_array_impl_data1_rsci_clken_d;
  output weight_mem_banks_bank_array_impl_data2_rsci_clken_d;
  output weight_mem_banks_bank_array_impl_data3_rsci_clken_d;
  output weight_mem_banks_bank_array_impl_data4_rsci_clken_d;
  output weight_mem_banks_bank_array_impl_data5_rsci_clken_d;
  output weight_mem_banks_bank_array_impl_data6_rsci_clken_d;
  output weight_mem_banks_bank_array_impl_data7_rsci_clken_d;
  output weight_mem_banks_bank_array_impl_data8_rsci_clken_d;
  output weight_mem_banks_bank_array_impl_data9_rsci_clken_d;
  output weight_mem_banks_bank_array_impl_data10_rsci_clken_d;
  output weight_mem_banks_bank_array_impl_data11_rsci_clken_d;
  output weight_mem_banks_bank_array_impl_data12_rsci_clken_d;
  output weight_mem_banks_bank_array_impl_data13_rsci_clken_d;
  output weight_mem_banks_bank_array_impl_data14_rsci_clken_d;
  output weight_mem_banks_bank_array_impl_data15_rsci_clken_d;
  output input_mem_banks_bank_array_impl_data0_rsci_clken_d;
  input PECoreRun_wen;
  input weight_mem_banks_bank_array_impl_data0_rsci_cgo;
  input weight_mem_banks_bank_array_impl_data0_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_array_impl_data1_rsci_cgo;
  input weight_mem_banks_bank_array_impl_data1_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_array_impl_data2_rsci_cgo;
  input weight_mem_banks_bank_array_impl_data2_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_array_impl_data3_rsci_cgo;
  input weight_mem_banks_bank_array_impl_data3_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_array_impl_data4_rsci_cgo;
  input weight_mem_banks_bank_array_impl_data4_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_array_impl_data5_rsci_cgo;
  input weight_mem_banks_bank_array_impl_data5_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_array_impl_data6_rsci_cgo;
  input weight_mem_banks_bank_array_impl_data6_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_array_impl_data7_rsci_cgo;
  input weight_mem_banks_bank_array_impl_data7_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_array_impl_data8_rsci_cgo;
  input weight_mem_banks_bank_array_impl_data8_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_array_impl_data9_rsci_cgo;
  input weight_mem_banks_bank_array_impl_data9_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_array_impl_data10_rsci_cgo;
  input weight_mem_banks_bank_array_impl_data10_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_array_impl_data11_rsci_cgo;
  input weight_mem_banks_bank_array_impl_data11_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_array_impl_data12_rsci_cgo;
  input weight_mem_banks_bank_array_impl_data12_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_array_impl_data13_rsci_cgo;
  input weight_mem_banks_bank_array_impl_data13_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_array_impl_data14_rsci_cgo;
  input weight_mem_banks_bank_array_impl_data14_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_array_impl_data15_rsci_cgo;
  input weight_mem_banks_bank_array_impl_data15_rsci_cgo_ir_unreg;
  input input_mem_banks_bank_array_impl_data0_rsci_cgo;
  input input_mem_banks_bank_array_impl_data0_rsci_cgo_ir_unreg;
  input Datapath_for_1_ProductSum_cmp_cgo;
  input Datapath_for_1_ProductSum_cmp_cgo_ir_unreg;
  output Datapath_for_1_ProductSum_cmp_ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  assign weight_mem_banks_bank_array_impl_data0_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_array_impl_data0_rsci_cgo
      | weight_mem_banks_bank_array_impl_data0_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_array_impl_data1_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_array_impl_data1_rsci_cgo
      | weight_mem_banks_bank_array_impl_data1_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_array_impl_data2_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_array_impl_data2_rsci_cgo
      | weight_mem_banks_bank_array_impl_data2_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_array_impl_data3_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_array_impl_data3_rsci_cgo
      | weight_mem_banks_bank_array_impl_data3_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_array_impl_data4_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_array_impl_data4_rsci_cgo
      | weight_mem_banks_bank_array_impl_data4_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_array_impl_data5_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_array_impl_data5_rsci_cgo
      | weight_mem_banks_bank_array_impl_data5_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_array_impl_data6_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_array_impl_data6_rsci_cgo
      | weight_mem_banks_bank_array_impl_data6_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_array_impl_data7_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_array_impl_data7_rsci_cgo
      | weight_mem_banks_bank_array_impl_data7_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_array_impl_data8_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_array_impl_data8_rsci_cgo
      | weight_mem_banks_bank_array_impl_data8_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_array_impl_data9_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_array_impl_data9_rsci_cgo
      | weight_mem_banks_bank_array_impl_data9_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_array_impl_data10_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_array_impl_data10_rsci_cgo
      | weight_mem_banks_bank_array_impl_data10_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_array_impl_data11_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_array_impl_data11_rsci_cgo
      | weight_mem_banks_bank_array_impl_data11_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_array_impl_data12_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_array_impl_data12_rsci_cgo
      | weight_mem_banks_bank_array_impl_data12_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_array_impl_data13_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_array_impl_data13_rsci_cgo
      | weight_mem_banks_bank_array_impl_data13_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_array_impl_data14_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_array_impl_data14_rsci_cgo
      | weight_mem_banks_bank_array_impl_data14_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_array_impl_data15_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_array_impl_data15_rsci_cgo
      | weight_mem_banks_bank_array_impl_data15_rsci_cgo_ir_unreg);
  assign input_mem_banks_bank_array_impl_data0_rsci_clken_d = PECoreRun_wen & (input_mem_banks_bank_array_impl_data0_rsci_cgo
      | input_mem_banks_bank_array_impl_data0_rsci_cgo_ir_unreg);
  assign Datapath_for_1_ProductSum_cmp_ccs_ccore_en = PECoreRun_wen & (Datapath_for_1_ProductSum_cmp_cgo
      | Datapath_for_1_ProductSum_cmp_cgo_ir_unreg);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp
    (
  clk, rst, input_port_PopNB_mioi_idat_mxwt, input_port_PopNB_mioi_ivld_mxwt, input_port_PopNB_mioi_biwt,
      input_port_PopNB_mioi_bdwt, input_port_PopNB_mioi_idat, input_port_PopNB_mioi_ivld
);
  input clk;
  input rst;
  output [136:0] input_port_PopNB_mioi_idat_mxwt;
  output input_port_PopNB_mioi_ivld_mxwt;
  input input_port_PopNB_mioi_biwt;
  input input_port_PopNB_mioi_bdwt;
  input [137:0] input_port_PopNB_mioi_idat;
  input input_port_PopNB_mioi_ivld;


  // Interconnect Declarations
  reg input_port_PopNB_mioi_bcwt;
  reg [137:0] input_port_PopNB_mioi_idat_bfwt;
  reg input_port_PopNB_mioi_ivld_bfwt;
  wire [137:0] input_port_PopNB_mioi_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  assign input_port_PopNB_mioi_idat_mxwt_pconst = MUX_v_138_2_2(input_port_PopNB_mioi_idat,
      input_port_PopNB_mioi_idat_bfwt, input_port_PopNB_mioi_bcwt);
  assign input_port_PopNB_mioi_ivld_mxwt = MUX_s_1_2_2(input_port_PopNB_mioi_ivld,
      input_port_PopNB_mioi_ivld_bfwt, input_port_PopNB_mioi_bcwt);
  assign input_port_PopNB_mioi_idat_mxwt = {(input_port_PopNB_mioi_idat_mxwt_pconst[137:130])
      , (input_port_PopNB_mioi_idat_mxwt_pconst[128:0])};
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      input_port_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      input_port_PopNB_mioi_bcwt <= ~((~(input_port_PopNB_mioi_bcwt | input_port_PopNB_mioi_biwt))
          | input_port_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      input_port_PopNB_mioi_idat_bfwt <= 138'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      input_port_PopNB_mioi_ivld_bfwt <= 1'b0;
    end
    else if ( input_port_PopNB_mioi_biwt ) begin
      input_port_PopNB_mioi_idat_bfwt <= input_port_PopNB_mioi_idat;
      input_port_PopNB_mioi_ivld_bfwt <= input_port_PopNB_mioi_ivld;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [137:0] MUX_v_138_2_2;
    input [137:0] input_0;
    input [137:0] input_1;
    input  sel;
    reg [137:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_138_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl
    (
  PECoreRun_wen, PECoreRun_wten, input_port_PopNB_mioi_oswt, input_port_PopNB_mioi_biwt,
      input_port_PopNB_mioi_bdwt
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input input_port_PopNB_mioi_oswt;
  output input_port_PopNB_mioi_biwt;
  output input_port_PopNB_mioi_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign input_port_PopNB_mioi_bdwt = input_port_PopNB_mioi_oswt & PECoreRun_wen;
  assign input_port_PopNB_mioi_biwt = (~ PECoreRun_wten) & input_port_PopNB_mioi_oswt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi (
  clk, rst, start_val, start_rdy, start_msg, PECoreRun_wen, PECoreRun_wten, start_PopNB_mioi_oswt,
      start_PopNB_mioi_idat_mxwt, start_PopNB_mioi_ivld_mxwt
);
  input clk;
  input rst;
  input start_val;
  output start_rdy;
  input start_msg;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_idat_mxwt;
  output start_PopNB_mioi_ivld_mxwt;


  // Interconnect Declarations
  wire start_PopNB_mioi_biwt;
  wire start_PopNB_mioi_bdwt;
  wire start_PopNB_mioi_idat;
  wire start_PopNB_mioi_ivld;


  // Interconnect Declarations for Component Instantiations 
  PECore_ccs_conn_in_wait_v1 #(.width(32'sd1),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) start_PopNB_mioi (
      .vld(start_val),
      .rdy(start_rdy),
      .dat(start_msg),
      .idat(start_PopNB_mioi_idat),
      .irdy(start_PopNB_mioi_biwt),
      .ivld(start_PopNB_mioi_ivld),
      .clk(clk),
      .en(1'b0),
      .arst(rst),
      .srst(1'b1)
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .start_PopNB_mioi_oswt(start_PopNB_mioi_oswt),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt)
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .start_PopNB_mioi_idat_mxwt(start_PopNB_mioi_idat_mxwt),
      .start_PopNB_mioi_ivld_mxwt(start_PopNB_mioi_ivld_mxwt),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_idat(start_PopNB_mioi_idat),
      .start_PopNB_mioi_ivld(start_PopNB_mioi_ivld)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi (
  clk, rst, rva_out_val, rva_out_rdy, rva_out_msg, PECoreRun_wen, rva_out_Push_mioi_oswt,
      rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_idat
);
  input clk;
  input rst;
  output rva_out_val;
  input rva_out_rdy;
  output [127:0] rva_out_msg;
  input PECoreRun_wen;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input [127:0] rva_out_Push_mioi_idat;


  // Interconnect Declarations
  wire rva_out_Push_mioi_biwt;
  wire rva_out_Push_mioi_bdwt;
  wire rva_out_Push_mioi_bcwt;
  wire rva_out_Push_mioi_ivld_PECoreRun_sct;
  wire rva_out_Push_mioi_irdy;


  // Interconnect Declarations for Component Instantiations 
  PECore_ccs_conn_out_wait_v1 #(.width(32'sd128),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) rva_out_Push_mioi (
      .vld(rva_out_val),
      .rdy(rva_out_rdy),
      .dat(rva_out_msg),
      .idat(rva_out_Push_mioi_idat),
      .clk(clk),
      .en(1'b0),
      .arst(rst),
      .srst(1'b1),
      .ivld(rva_out_Push_mioi_ivld_PECoreRun_sct),
      .irdy(rva_out_Push_mioi_irdy)
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .rva_out_Push_mioi_oswt(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_bdwt(rva_out_Push_mioi_bdwt),
      .rva_out_Push_mioi_bcwt(rva_out_Push_mioi_bcwt),
      .rva_out_Push_mioi_ivld_PECoreRun_sct(rva_out_Push_mioi_ivld_PECoreRun_sct),
      .rva_out_Push_mioi_irdy(rva_out_Push_mioi_irdy)
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_Push_mioi_oswt(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_bdwt(rva_out_Push_mioi_bdwt),
      .rva_out_Push_mioi_bcwt(rva_out_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi (
  clk, rst, act_port_val, act_port_rdy, act_port_msg, PECoreRun_wen, act_port_Push_mioi_oswt,
      act_port_Push_mioi_wen_comp, act_port_Push_mioi_idat
);
  input clk;
  input rst;
  output act_port_val;
  input act_port_rdy;
  output [319:0] act_port_msg;
  input PECoreRun_wen;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_wen_comp;
  input [319:0] act_port_Push_mioi_idat;


  // Interconnect Declarations
  wire act_port_Push_mioi_biwt;
  wire act_port_Push_mioi_bdwt;
  wire act_port_Push_mioi_bcwt;
  wire act_port_Push_mioi_ivld_PECoreRun_sct;
  wire act_port_Push_mioi_irdy;


  // Interconnect Declarations for Component Instantiations 
  PECore_ccs_conn_out_wait_v1 #(.width(32'sd320),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) act_port_Push_mioi (
      .vld(act_port_val),
      .rdy(act_port_rdy),
      .dat(act_port_msg),
      .idat(act_port_Push_mioi_idat),
      .clk(clk),
      .en(1'b0),
      .arst(rst),
      .srst(1'b1),
      .ivld(act_port_Push_mioi_ivld_PECoreRun_sct),
      .irdy(act_port_Push_mioi_irdy)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .act_port_Push_mioi_oswt(act_port_Push_mioi_oswt),
      .act_port_Push_mioi_biwt(act_port_Push_mioi_biwt),
      .act_port_Push_mioi_bdwt(act_port_Push_mioi_bdwt),
      .act_port_Push_mioi_bcwt(act_port_Push_mioi_bcwt),
      .act_port_Push_mioi_ivld_PECoreRun_sct(act_port_Push_mioi_ivld_PECoreRun_sct),
      .act_port_Push_mioi_irdy(act_port_Push_mioi_irdy)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_port_Push_mioi_oswt(act_port_Push_mioi_oswt),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .act_port_Push_mioi_biwt(act_port_Push_mioi_biwt),
      .act_port_Push_mioi_bdwt(act_port_Push_mioi_bdwt),
      .act_port_Push_mioi_bcwt(act_port_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi (
  clk, rst, rva_in_val, rva_in_rdy, rva_in_msg, PECoreRun_wen, PECoreRun_wten, rva_in_PopNB_mioi_oswt,
      rva_in_PopNB_mioi_idat_mxwt, rva_in_PopNB_mioi_ivld_mxwt
);
  input clk;
  input rst;
  input rva_in_val;
  output rva_in_rdy;
  input [168:0] rva_in_msg;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output [168:0] rva_in_PopNB_mioi_idat_mxwt;
  output rva_in_PopNB_mioi_ivld_mxwt;


  // Interconnect Declarations
  wire rva_in_PopNB_mioi_biwt;
  wire rva_in_PopNB_mioi_bdwt;
  wire [168:0] rva_in_PopNB_mioi_idat;
  wire rva_in_PopNB_mioi_ivld;


  // Interconnect Declarations for Component Instantiations 
  PECore_ccs_conn_in_wait_v1 #(.width(32'sd169),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) rva_in_PopNB_mioi (
      .vld(rva_in_val),
      .rdy(rva_in_rdy),
      .dat(rva_in_msg),
      .idat(rva_in_PopNB_mioi_idat),
      .irdy(rva_in_PopNB_mioi_biwt),
      .ivld(rva_in_PopNB_mioi_ivld),
      .clk(clk),
      .en(1'b0),
      .arst(rst),
      .srst(1'b1)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .rva_in_PopNB_mioi_oswt(rva_in_PopNB_mioi_oswt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_PopNB_mioi_idat_mxwt(rva_in_PopNB_mioi_idat_mxwt),
      .rva_in_PopNB_mioi_ivld_mxwt(rva_in_PopNB_mioi_ivld_mxwt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_idat(rva_in_PopNB_mioi_idat),
      .rva_in_PopNB_mioi_ivld(rva_in_PopNB_mioi_ivld)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi (
  clk, rst, input_port_val, input_port_rdy, input_port_msg, PECoreRun_wen, PECoreRun_wten,
      input_port_PopNB_mioi_oswt, input_port_PopNB_mioi_idat_mxwt, input_port_PopNB_mioi_ivld_mxwt
);
  input clk;
  input rst;
  input input_port_val;
  output input_port_rdy;
  input [137:0] input_port_msg;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input input_port_PopNB_mioi_oswt;
  output [136:0] input_port_PopNB_mioi_idat_mxwt;
  output input_port_PopNB_mioi_ivld_mxwt;


  // Interconnect Declarations
  wire input_port_PopNB_mioi_biwt;
  wire input_port_PopNB_mioi_bdwt;
  wire [137:0] input_port_PopNB_mioi_idat;
  wire input_port_PopNB_mioi_ivld;
  wire [136:0] input_port_PopNB_mioi_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  PECore_ccs_conn_in_wait_v1 #(.width(32'sd138),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) input_port_PopNB_mioi (
      .vld(input_port_val),
      .rdy(input_port_rdy),
      .dat(input_port_msg),
      .idat(input_port_PopNB_mioi_idat),
      .irdy(input_port_PopNB_mioi_biwt),
      .ivld(input_port_PopNB_mioi_ivld),
      .clk(clk),
      .en(1'b0),
      .arst(rst),
      .srst(1'b1)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .input_port_PopNB_mioi_oswt(input_port_PopNB_mioi_oswt),
      .input_port_PopNB_mioi_biwt(input_port_PopNB_mioi_biwt),
      .input_port_PopNB_mioi_bdwt(input_port_PopNB_mioi_bdwt)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .input_port_PopNB_mioi_idat_mxwt(input_port_PopNB_mioi_idat_mxwt_pconst),
      .input_port_PopNB_mioi_ivld_mxwt(input_port_PopNB_mioi_ivld_mxwt),
      .input_port_PopNB_mioi_biwt(input_port_PopNB_mioi_biwt),
      .input_port_PopNB_mioi_bdwt(input_port_PopNB_mioi_bdwt),
      .input_port_PopNB_mioi_idat(input_port_PopNB_mioi_idat),
      .input_port_PopNB_mioi_ivld(input_port_PopNB_mioi_ivld)
    );
  assign input_port_PopNB_mioi_idat_mxwt = input_port_PopNB_mioi_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun (
  clk, rst, start_val, start_rdy, start_msg, input_port_val, input_port_rdy, input_port_msg,
      rva_in_val, rva_in_rdy, rva_in_msg, rva_out_val, rva_out_rdy, rva_out_msg,
      act_port_val, act_port_rdy, act_port_msg, SC_SRAM_CONFIG, weight_mem_banks_bank_array_impl_data0_rsci_clken_d,
      weight_mem_banks_bank_array_impl_data0_rsci_d_d, weight_mem_banks_bank_array_impl_data0_rsci_q_d,
      weight_mem_banks_bank_array_impl_data0_rsci_radr_d, weight_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data1_rsci_clken_d, weight_mem_banks_bank_array_impl_data1_rsci_d_d,
      weight_mem_banks_bank_array_impl_data1_rsci_q_d, weight_mem_banks_bank_array_impl_data1_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data1_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data2_rsci_clken_d, weight_mem_banks_bank_array_impl_data2_rsci_d_d,
      weight_mem_banks_bank_array_impl_data2_rsci_q_d, weight_mem_banks_bank_array_impl_data2_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data2_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data3_rsci_clken_d, weight_mem_banks_bank_array_impl_data3_rsci_d_d,
      weight_mem_banks_bank_array_impl_data3_rsci_q_d, weight_mem_banks_bank_array_impl_data3_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data3_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data4_rsci_clken_d, weight_mem_banks_bank_array_impl_data4_rsci_d_d,
      weight_mem_banks_bank_array_impl_data4_rsci_q_d, weight_mem_banks_bank_array_impl_data4_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data4_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data5_rsci_clken_d, weight_mem_banks_bank_array_impl_data5_rsci_d_d,
      weight_mem_banks_bank_array_impl_data5_rsci_q_d, weight_mem_banks_bank_array_impl_data5_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data5_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data6_rsci_clken_d, weight_mem_banks_bank_array_impl_data6_rsci_d_d,
      weight_mem_banks_bank_array_impl_data6_rsci_q_d, weight_mem_banks_bank_array_impl_data6_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data6_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data7_rsci_clken_d, weight_mem_banks_bank_array_impl_data7_rsci_d_d,
      weight_mem_banks_bank_array_impl_data7_rsci_q_d, weight_mem_banks_bank_array_impl_data7_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data7_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data8_rsci_clken_d, weight_mem_banks_bank_array_impl_data8_rsci_d_d,
      weight_mem_banks_bank_array_impl_data8_rsci_q_d, weight_mem_banks_bank_array_impl_data8_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data8_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data9_rsci_clken_d, weight_mem_banks_bank_array_impl_data9_rsci_d_d,
      weight_mem_banks_bank_array_impl_data9_rsci_q_d, weight_mem_banks_bank_array_impl_data9_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data9_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data10_rsci_clken_d, weight_mem_banks_bank_array_impl_data10_rsci_d_d,
      weight_mem_banks_bank_array_impl_data10_rsci_q_d, weight_mem_banks_bank_array_impl_data10_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data10_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data11_rsci_clken_d, weight_mem_banks_bank_array_impl_data11_rsci_d_d,
      weight_mem_banks_bank_array_impl_data11_rsci_q_d, weight_mem_banks_bank_array_impl_data11_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data11_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data12_rsci_clken_d, weight_mem_banks_bank_array_impl_data12_rsci_d_d,
      weight_mem_banks_bank_array_impl_data12_rsci_q_d, weight_mem_banks_bank_array_impl_data12_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data12_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data13_rsci_clken_d, weight_mem_banks_bank_array_impl_data13_rsci_d_d,
      weight_mem_banks_bank_array_impl_data13_rsci_q_d, weight_mem_banks_bank_array_impl_data13_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data13_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data14_rsci_clken_d, weight_mem_banks_bank_array_impl_data14_rsci_d_d,
      weight_mem_banks_bank_array_impl_data14_rsci_q_d, weight_mem_banks_bank_array_impl_data14_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data14_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data15_rsci_clken_d, weight_mem_banks_bank_array_impl_data15_rsci_d_d,
      weight_mem_banks_bank_array_impl_data15_rsci_q_d, weight_mem_banks_bank_array_impl_data15_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data15_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      input_mem_banks_bank_array_impl_data0_rsci_clken_d, input_mem_banks_bank_array_impl_data0_rsci_d_d,
      input_mem_banks_bank_array_impl_data0_rsci_q_d, input_mem_banks_bank_array_impl_data0_rsci_radr_d,
      input_mem_banks_bank_array_impl_data0_rsci_wadr_d, input_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_pff, weight_mem_banks_bank_array_impl_data0_rsci_we_d_pff,
      weight_mem_banks_bank_array_impl_data1_rsci_we_d_pff, weight_mem_banks_bank_array_impl_data2_rsci_we_d_pff,
      weight_mem_banks_bank_array_impl_data3_rsci_we_d_pff, weight_mem_banks_bank_array_impl_data4_rsci_we_d_pff,
      weight_mem_banks_bank_array_impl_data5_rsci_we_d_pff, weight_mem_banks_bank_array_impl_data6_rsci_we_d_pff,
      weight_mem_banks_bank_array_impl_data7_rsci_we_d_pff, weight_mem_banks_bank_array_impl_data8_rsci_we_d_pff,
      weight_mem_banks_bank_array_impl_data9_rsci_we_d_pff, weight_mem_banks_bank_array_impl_data10_rsci_we_d_pff,
      weight_mem_banks_bank_array_impl_data11_rsci_we_d_pff, weight_mem_banks_bank_array_impl_data12_rsci_we_d_pff,
      weight_mem_banks_bank_array_impl_data13_rsci_we_d_pff, weight_mem_banks_bank_array_impl_data14_rsci_we_d_pff,
      weight_mem_banks_bank_array_impl_data15_rsci_we_d_pff, input_mem_banks_bank_array_impl_data0_rsci_we_d_pff
);
  input clk;
  input rst;
  input start_val;
  output start_rdy;
  input start_msg;
  input input_port_val;
  output input_port_rdy;
  input [137:0] input_port_msg;
  input rva_in_val;
  output rva_in_rdy;
  input [168:0] rva_in_msg;
  output rva_out_val;
  input rva_out_rdy;
  output [127:0] rva_out_msg;
  output act_port_val;
  input act_port_rdy;
  output [319:0] act_port_msg;
  input [31:0] SC_SRAM_CONFIG;
  output weight_mem_banks_bank_array_impl_data0_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data0_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data0_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data0_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data1_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data1_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data1_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data1_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data1_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data2_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data2_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data2_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data2_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data2_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data3_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data3_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data3_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data3_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data3_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data4_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data4_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data4_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data4_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data4_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data5_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data5_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data5_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data5_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data5_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data6_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data6_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data6_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data6_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data6_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data7_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data7_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data7_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data7_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data7_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data8_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data8_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data8_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data8_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data8_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data9_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data9_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data9_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data9_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data9_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data10_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data10_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data10_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data10_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data10_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data11_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data11_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data11_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data11_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data11_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data12_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data12_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data12_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data12_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data12_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data13_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data13_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data13_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data13_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data13_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data14_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data14_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data14_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data14_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data14_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data15_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data15_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data15_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data15_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data15_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output input_mem_banks_bank_array_impl_data0_rsci_clken_d;
  output [127:0] input_mem_banks_bank_array_impl_data0_rsci_d_d;
  input [127:0] input_mem_banks_bank_array_impl_data0_rsci_q_d;
  output [7:0] input_mem_banks_bank_array_impl_data0_rsci_radr_d;
  output [7:0] input_mem_banks_bank_array_impl_data0_rsci_wadr_d;
  output input_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output [11:0] weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_pff;
  output weight_mem_banks_bank_array_impl_data0_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data1_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data2_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data3_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data4_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data5_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data6_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data7_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data8_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data9_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data10_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data11_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data12_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data13_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data14_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data15_rsci_we_d_pff;
  output input_mem_banks_bank_array_impl_data0_rsci_we_d_pff;


  // Interconnect Declarations
  wire PECoreRun_wen;
  wire PECoreRun_wten;
  wire [136:0] input_port_PopNB_mioi_idat_mxwt;
  wire input_port_PopNB_mioi_ivld_mxwt;
  wire [168:0] rva_in_PopNB_mioi_idat_mxwt;
  wire rva_in_PopNB_mioi_ivld_mxwt;
  wire act_port_Push_mioi_wen_comp;
  wire rva_out_Push_mioi_wen_comp;
  wire start_PopNB_mioi_idat_mxwt;
  wire start_PopNB_mioi_ivld_mxwt;
  wire [31:0] Datapath_for_1_ProductSum_cmp_out_rsc_z;
  wire Datapath_for_1_ProductSum_cmp_ccs_ccore_en;
  wire [31:0] Datapath_for_1_ProductSum_cmp_1_out_rsc_z;
  wire [31:0] Datapath_for_1_ProductSum_cmp_2_out_rsc_z;
  wire [31:0] Datapath_for_1_ProductSum_cmp_3_out_rsc_z;
  wire [12:0] PEManager_16U_GetWeightAddr_if_acc_4_cmp_z;
  reg [19:0] act_port_Push_mioi_idat_319_300;
  reg [19:0] act_port_Push_mioi_idat_299_280;
  reg [19:0] act_port_Push_mioi_idat_279_260;
  reg [19:0] act_port_Push_mioi_idat_259_240;
  reg [19:0] act_port_Push_mioi_idat_239_220;
  reg [19:0] act_port_Push_mioi_idat_219_200;
  reg [19:0] act_port_Push_mioi_idat_199_180;
  reg [19:0] act_port_Push_mioi_idat_179_160;
  reg [19:0] act_port_Push_mioi_idat_159_140;
  reg [19:0] act_port_Push_mioi_idat_139_120;
  reg [19:0] act_port_Push_mioi_idat_119_100;
  reg [19:0] act_port_Push_mioi_idat_99_80;
  reg [19:0] act_port_Push_mioi_idat_79_60;
  reg [19:0] act_port_Push_mioi_idat_59_40;
  reg [19:0] act_port_Push_mioi_idat_39_20;
  reg [19:0] act_port_Push_mioi_idat_19_0;
  reg [7:0] rva_out_Push_mioi_idat_127_120;
  reg [7:0] rva_out_Push_mioi_idat_119_112;
  reg [7:0] rva_out_Push_mioi_idat_111_104;
  reg [7:0] rva_out_Push_mioi_idat_103_96;
  reg [7:0] rva_out_Push_mioi_idat_95_88;
  reg [7:0] rva_out_Push_mioi_idat_87_80;
  reg [7:0] rva_out_Push_mioi_idat_79_72;
  reg [7:0] rva_out_Push_mioi_idat_71_64;
  reg [7:0] rva_out_Push_mioi_idat_63_56;
  reg [7:0] rva_out_Push_mioi_idat_55_48;
  reg [7:0] rva_out_Push_mioi_idat_47_40;
  reg [3:0] rva_out_Push_mioi_idat_39_36;
  reg [3:0] rva_out_Push_mioi_idat_35_32;
  reg [4:0] rva_out_Push_mioi_idat_31_27;
  reg [1:0] rva_out_Push_mioi_idat_26_25;
  reg rva_out_Push_mioi_idat_24;
  reg [4:0] rva_out_Push_mioi_idat_23_19;
  reg [1:0] rva_out_Push_mioi_idat_18_17;
  reg rva_out_Push_mioi_idat_16;
  reg [4:0] rva_out_Push_mioi_idat_15_11;
  reg [1:0] rva_out_Push_mioi_idat_10_9;
  reg rva_out_Push_mioi_idat_8;
  reg [6:0] rva_out_Push_mioi_idat_7_1;
  reg rva_out_Push_mioi_idat_0;
  wire [4:0] fsm_output;
  wire [8:0] operator_16_false_acc_tmp;
  wire [9:0] nl_operator_16_false_acc_tmp;
  wire [8:0] operator_8_false_acc_tmp;
  wire [9:0] nl_operator_8_false_acc_tmp;
  wire [4:0] operator_4_false_acc_tmp;
  wire [5:0] nl_operator_4_false_acc_tmp;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_239_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_238_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_237_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_236_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_235_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_234_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_232_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_231_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_230_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_229_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_228_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_227_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_226_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_225_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_224_tmp;
  wire [15:0] weight_mem_write_arbxbar_xbar_for_lshift_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_16_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_15_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_15_Arbiter_16U_Roundrobin_pick_priority_and_4_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_14_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_14_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_13_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_13_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_12_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_12_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_11_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_11_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_10_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_10_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_9_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_9_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_8_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_8_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_7_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_7_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_6_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_6_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_5_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_5_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_4_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_4_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_3_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_3_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_2_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_1_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_16_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_2_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_15_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_3_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_14_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_4_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_13_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_5_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_12_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_6_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_11_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_7_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_10_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_8_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_9_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_1_lshift_tmp;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_nor_7_tmp;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_nor_9_tmp;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_nor_11_tmp;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_nor_13_tmp;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_nor_15_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_233_tmp;
  wire or_tmp_18;
  wire or_tmp_20;
  wire or_dcpl;
  wire or_dcpl_34;
  wire and_dcpl_135;
  wire and_dcpl_210;
  wire and_dcpl_211;
  wire or_tmp_545;
  wire or_dcpl_247;
  wire and_dcpl_414;
  wire or_dcpl_251;
  wire or_tmp_1286;
  wire or_dcpl_285;
  wire or_dcpl_286;
  wire and_dcpl_437;
  wire and_dcpl_439;
  wire or_dcpl_295;
  wire and_dcpl_440;
  wire or_dcpl_300;
  wire or_dcpl_301;
  wire or_dcpl_302;
  wire or_dcpl_306;
  wire or_dcpl_310;
  wire or_dcpl_313;
  wire or_dcpl_327;
  wire or_dcpl_334;
  wire or_dcpl_362;
  wire or_dcpl_363;
  wire or_dcpl_364;
  wire or_dcpl_365;
  wire or_dcpl_369;
  wire and_dcpl_700;
  wire and_dcpl_702;
  wire or_dcpl_370;
  wire and_dcpl_704;
  wire and_dcpl_705;
  wire and_dcpl_706;
  wire and_dcpl_707;
  wire and_dcpl_708;
  wire and_dcpl_709;
  wire or_dcpl_374;
  wire or_dcpl_375;
  wire or_dcpl_378;
  wire and_dcpl_725;
  wire and_dcpl_726;
  wire and_dcpl_733;
  wire and_dcpl_748;
  wire and_dcpl_749;
  wire and_dcpl_756;
  wire and_dcpl_771;
  wire and_dcpl_772;
  wire and_dcpl_779;
  wire and_dcpl_794;
  wire and_dcpl_795;
  wire and_dcpl_802;
  wire and_dcpl_817;
  wire and_dcpl_818;
  wire and_dcpl_825;
  wire and_dcpl_840;
  wire and_dcpl_841;
  wire and_dcpl_848;
  wire and_dcpl_863;
  wire and_dcpl_864;
  wire and_dcpl_871;
  wire and_dcpl_886;
  wire and_dcpl_887;
  wire and_dcpl_894;
  wire and_dcpl_909;
  wire and_dcpl_910;
  wire and_dcpl_917;
  wire and_dcpl_932;
  wire and_dcpl_933;
  wire and_dcpl_939;
  wire and_dcpl_954;
  wire and_dcpl_955;
  wire and_dcpl_962;
  wire and_dcpl_977;
  wire and_dcpl_978;
  wire and_dcpl_985;
  wire and_dcpl_1000;
  wire and_dcpl_1001;
  wire and_dcpl_1008;
  wire and_dcpl_1023;
  wire and_dcpl_1024;
  wire and_dcpl_1029;
  wire and_dcpl_1043;
  wire and_dcpl_1044;
  wire and_dcpl_1051;
  wire and_dcpl_1066;
  wire and_dcpl_1067;
  wire and_dcpl_1074;
  wire or_tmp_1334;
  wire or_tmp_1655;
  wire or_tmp_2232;
  wire or_tmp_2557;
  wire PECore_RunMac_PECore_RunMac_and_2_cse;
  wire PECore_UpdateFSM_switch_lp_nor_6_cse;
  wire and_2164_cse;
  wire and_2907_cse;
  wire and_4616_cse;
  reg PECore_RunMac_nor_tmp;
  reg pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_pe_config_UpdateInputCounter_if_nor_svs;
  reg PECore_RunFSM_switch_lp_equal_tmp;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_1;
  reg PECore_RunFSM_switch_lp_equal_tmp_1;
  reg PECore_RunFSM_switch_lp_equal_tmp_2;
  reg state_2_0_sva_2;
  reg pe_config_is_valid_sva;
  reg is_start_sva;
  reg input_mem_banks_load_store_for_else_and_cse;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm;
  reg PECore_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva;
  reg PECore_CheckStart_start_reg_sva;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp;
  reg [168:0] rva_in_PopNB_mio_mrgout_dat_sva;
  reg PECore_DecodeAxiRead_switch_lp_nor_2_itm;
  reg state_2_0_sva_0;
  reg state_2_0_sva_1;
  wire input_mem_banks_load_store_for_else_and_cse_1;
  reg input_read_req_valid_lpi_1_dfm_5;
  reg input_write_req_valid_lpi_1_dfm_5;
  wire pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1;
  wire pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_nor_svs_1;
  wire pe_config_is_zero_first_sva_dfm_4_mx0;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
  wire PECore_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_mx1;
  wire weight_read_ack_15_lpi_1_dfm_15_mx0;
  wire weight_read_ack_14_lpi_1_dfm_15_mx0;
  wire weight_read_ack_13_lpi_1_dfm_15_mx0;
  wire weight_read_ack_12_lpi_1_dfm_15_mx0;
  wire weight_read_ack_11_lpi_1_dfm_15_mx0;
  wire weight_read_ack_10_lpi_1_dfm_15_mx0;
  wire weight_read_ack_8_lpi_1_dfm_15_mx0;
  wire weight_read_ack_7_lpi_1_dfm_15_mx0;
  wire weight_read_ack_6_lpi_1_dfm_15_mx0;
  wire weight_read_ack_5_lpi_1_dfm_15_mx0;
  wire weight_read_ack_4_lpi_1_dfm_15_mx0;
  wire weight_read_ack_3_lpi_1_dfm_15_mx0;
  wire weight_read_ack_2_lpi_1_dfm_15_mx0;
  wire weight_read_ack_1_lpi_1_dfm_15_mx0;
  wire weight_read_ack_0_lpi_1_dfm_15_mx0;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_15_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_2_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_15_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_15_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_15_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_15_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_15_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_15_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_15_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_15_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_15_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_15_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_15_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_2_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_2_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_2_1_sva_1;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_15_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_15_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_15_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_15_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_15_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_15_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_14_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_14_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_14_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_14_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_14_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_14_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_13_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_13_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_13_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_13_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_13_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_13_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_12_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_12_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_12_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_12_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_12_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_12_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_11_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_11_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_11_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_11_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_11_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_11_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_10_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_10_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_10_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_10_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_10_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_10_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_9_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_9_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_9_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_9_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_9_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_9_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_8_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_8_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_8_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_8_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_8_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_8_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_7_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_7_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_7_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_7_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_7_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_7_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_6_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_6_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_6_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_6_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_6_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_6_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_5_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_5_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_5_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_5_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_5_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_5_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_4_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_4_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_4_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_4_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_4_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_4_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_3_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_3_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_3_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_2_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_2_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_2_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_1_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_1_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_1_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_0_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_7_sva;
  wire [168:0] rva_in_PopNB_mio_mrgout_dat_sva_1;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_nor_tmp_1;
  wire PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_5;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_31;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_4;
  wire PECore_DecodeAxiRead_switch_lp_nor_tmp_mx0w0;
  wire PECore_RunFSM_switch_lp_equal_tmp_3;
  reg pe_config_is_bias_sva;
  wire PECore_RunFSM_switch_lp_nor_3_cse_1;
  wire PECore_RunFSM_switch_lp_equal_tmp_5;
  wire PECore_RunFSM_switch_lp_equal_tmp_4;
  wire PECore_RunBias_if_for_11_operator_32_true_slc_operator_32_true_acc_13_svs_mx0;
  reg while_and_46_tmp_1;
  wire PECore_RunBias_if_for_10_operator_32_true_slc_operator_32_true_acc_13_svs_mx0;
  wire PECore_RunBias_if_for_7_operator_32_true_slc_operator_32_true_acc_13_svs_mx0;
  wire PECore_RunBias_if_for_6_operator_32_true_slc_operator_32_true_acc_13_svs_mx0;
  wire PECore_RunBias_if_for_2_operator_32_true_slc_operator_32_true_acc_13_svs_mx2;
  wire PECore_RunBias_if_for_12_operator_32_true_slc_operator_32_true_acc_13_svs_mx2;
  wire PECore_RunBias_if_for_1_operator_32_true_slc_operator_32_true_acc_13_svs_mx2;
  wire PECore_RunBias_if_for_16_operator_32_true_slc_operator_32_true_acc_13_svs_mx1;
  wire while_and_48_tmp_1;
  wire PECore_RunBias_if_for_15_operator_32_true_slc_operator_32_true_acc_13_svs_mx1;
  wire PECore_RunBias_if_for_14_operator_32_true_slc_operator_32_true_acc_13_svs_mx1;
  wire PECore_RunBias_if_for_13_operator_32_true_slc_operator_32_true_acc_13_svs_mx1;
  wire weight_read_ack_9_lpi_1_dfm_15_mx0;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  reg while_stage_0_2;
  reg while_asn_41_itm_1;
  reg adpfloat_tmp_is_zero_land_11_lpi_1_dfm;
  reg adpfloat_tmp_is_zero_land_11_lpi_1_dfm_st;
  reg adpfloat_tmp_is_zero_land_10_lpi_1_dfm;
  reg adpfloat_tmp_is_zero_land_10_lpi_1_dfm_st;
  reg PECore_UpdateFSM_case_4_is_output_end_pe_config_UpdateManagerCounter_nand_itm;
  reg PECore_UpdateFSM_switch_lp_unequal_tmp;
  reg [127:0] input_mem_banks_read_read_data_lpi_1;
  reg adpfloat_tmp_is_zero_land_7_lpi_1_dfm;
  reg adpfloat_tmp_is_zero_land_7_lpi_1_dfm_st;
  reg adpfloat_tmp_is_zero_land_6_lpi_1_dfm;
  reg adpfloat_tmp_is_zero_land_6_lpi_1_dfm_st;
  reg while_and_29_itm_1;
  reg while_and_30_itm_1;
  reg PECore_RunBias_if_for_14_operator_32_true_slc_operator_32_true_acc_13_svs;
  reg PECore_RunBias_if_for_15_operator_32_true_slc_operator_32_true_acc_13_svs;
  reg PECore_RunBias_if_for_13_operator_32_true_slc_operator_32_true_acc_13_svs;
  reg PECore_RunBias_if_for_16_operator_32_true_slc_operator_32_true_acc_13_svs;
  reg PECore_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva;
  reg w_axi_rsp_lpi_1_dfm_1;
  reg pe_config_is_zero_first_sva;
  reg pe_manager_zero_active_1_sva;
  reg pe_manager_zero_active_0_sva;
  reg pe_config_is_cluster_sva;
  reg [3:0] pe_config_manager_counter_sva;
  reg [15:0] weight_mem_write_arbxbar_xbar_for_empty_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_16_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_15_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_14_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_13_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_12_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_11_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_10_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_9_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_8_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_7_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_6_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_5_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_4_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_3_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_2_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_1_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg PECore_DecodeAxiRead_case_4_switch_lp_and_2_itm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_15_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_14_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_13_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_9_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_11_lpi_1_dfm;
  wire [31:0] PECore_RunBias_if_accum_vector_out_data_11_lpi_1_dfm_mx2;
  wire [31:0] PECore_RunBias_if_accum_vector_out_data_10_lpi_1_dfm_mx2;
  wire [31:0] PECore_RunBias_if_accum_vector_out_data_7_lpi_1_dfm_mx2;
  wire [31:0] PECore_RunBias_if_accum_vector_out_data_6_lpi_1_dfm_mx2;
  wire pe_config_manager_counter_sva_dfm_4_mx0_0;
  reg PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva;
  wire while_and_71_m1c;
  wire while_and_73_m1c;
  wire while_and_65_m1c;
  wire while_and_79_m1c;
  wire while_and_63_m1c;
  wire while_and_61_m1c;
  wire while_and_59_m1c;
  wire while_and_57_m1c;
  wire while_and_87_m1c;
  wire while_and_85_m1c;
  wire while_and_83_m1c;
  wire while_and_81_m1c;
  reg [19:0] reg_PECore_RunBias_if_accum_vector_out_data_11_lpi_1_dfm_ftd_12;
  reg [19:0] reg_PECore_RunBias_if_accum_vector_out_data_10_lpi_1_dfm_ftd_12;
  reg [19:0] reg_PECore_RunBias_if_accum_vector_out_data_7_lpi_1_dfm_ftd_12;
  reg [19:0] reg_PECore_RunBias_if_accum_vector_out_data_6_lpi_1_dfm_ftd_12;
  wire while_and_67_m1c;
  wire while_and_69_m1c;
  wire while_and_75_m1c;
  wire while_and_77_m1c;
  wire weight_mem_banks_write_if_for_if_mux_cse;
  wire weight_mem_banks_write_if_for_if_mux_1_cse;
  wire weight_mem_banks_read_for_mux_cse;
  wire weight_mem_banks_read_for_mux_1_cse;
  wire weight_mem_banks_write_if_for_if_mux_4_cse;
  wire weight_mem_banks_write_if_for_if_mux_5_cse;
  wire weight_mem_banks_read_for_mux_4_cse;
  wire weight_mem_banks_read_for_mux_5_cse;
  wire weight_mem_banks_write_if_for_if_mux_8_cse;
  wire weight_mem_banks_write_if_for_if_mux_9_cse;
  wire weight_mem_banks_read_for_mux_8_cse;
  wire weight_mem_banks_read_for_mux_9_cse;
  wire weight_mem_banks_write_if_for_if_mux_12_cse;
  wire weight_mem_banks_write_if_for_if_mux_13_cse;
  wire weight_mem_banks_read_for_mux_12_cse;
  wire weight_mem_banks_read_for_mux_13_cse;
  wire weight_mem_banks_write_if_for_if_mux_16_cse;
  wire weight_mem_banks_write_if_for_if_mux_17_cse;
  wire weight_mem_banks_read_for_mux_16_cse;
  wire weight_mem_banks_read_for_mux_17_cse;
  wire weight_mem_banks_write_if_for_if_mux_20_cse;
  wire weight_mem_banks_write_if_for_if_mux_21_cse;
  wire weight_mem_banks_read_for_mux_20_cse;
  wire weight_mem_banks_read_for_mux_21_cse;
  wire weight_mem_banks_write_if_for_if_mux_24_cse;
  wire weight_mem_banks_write_if_for_if_mux_25_cse;
  wire weight_mem_banks_read_for_mux_24_cse;
  wire weight_mem_banks_read_for_mux_25_cse;
  wire weight_mem_banks_write_if_for_if_mux_28_cse;
  wire weight_mem_banks_write_if_for_if_mux_29_cse;
  wire weight_mem_banks_read_for_mux_28_cse;
  wire weight_mem_banks_read_for_mux_29_cse;
  wire weight_mem_banks_write_if_for_if_mux_32_cse;
  wire weight_mem_banks_write_if_for_if_mux_33_cse;
  wire weight_mem_banks_read_for_mux_32_cse;
  wire weight_mem_banks_read_for_mux_33_cse;
  wire weight_mem_banks_write_if_for_if_mux_36_cse;
  wire weight_mem_banks_write_if_for_if_mux_37_cse;
  wire weight_mem_banks_read_for_mux_36_cse;
  wire weight_mem_banks_read_for_mux_37_cse;
  wire weight_mem_banks_write_if_for_if_mux_40_cse;
  wire weight_mem_banks_write_if_for_if_mux_41_cse;
  wire weight_mem_banks_read_for_mux_40_cse;
  wire weight_mem_banks_read_for_mux_41_cse;
  wire weight_mem_banks_write_if_for_if_mux_44_cse;
  wire weight_mem_banks_write_if_for_if_mux_45_cse;
  wire weight_mem_banks_read_for_mux_44_cse;
  wire weight_mem_banks_read_for_mux_45_cse;
  wire weight_mem_banks_write_if_for_if_mux_48_cse;
  wire weight_mem_banks_write_if_for_if_mux_49_cse;
  wire weight_mem_banks_read_for_mux_48_cse;
  wire weight_mem_banks_read_for_mux_49_cse;
  wire weight_mem_banks_write_if_for_if_mux_52_cse;
  wire weight_mem_banks_write_if_for_if_mux_53_cse;
  wire weight_mem_banks_read_for_mux_52_cse;
  wire weight_mem_banks_read_for_mux_53_cse;
  wire weight_mem_banks_write_if_for_if_mux_56_cse;
  wire weight_mem_banks_write_if_for_if_mux_57_cse;
  wire weight_mem_banks_read_for_mux_56_cse;
  wire weight_mem_banks_read_for_mux_57_cse;
  wire weight_mem_banks_write_if_for_if_mux_60_cse;
  wire weight_mem_banks_write_if_for_if_mux_61_cse;
  wire weight_mem_banks_read_for_mux_60_cse;
  wire weight_mem_banks_read_for_mux_61_cse;
  wire input_mem_banks_write_if_for_if_mux_1_cse;
  wire input_mem_banks_write_if_for_if_mux_2_cse;
  wire input_mem_banks_read_for_mux_cse;
  wire input_mem_banks_read_for_mux_1_cse;
  reg reg_input_port_PopNB_mioi_oswt_cse;
  reg reg_rva_in_PopNB_mioi_oswt_cse;
  wire PECore_RunMac_if_and_208_cse;
  wire PECore_RunMac_if_and_209_cse;
  wire PECore_RunMac_if_and_176_cse;
  wire PECore_RunMac_if_and_177_cse;
  wire PECore_RunMac_if_and_144_cse;
  wire PECore_RunMac_if_and_145_cse;
  wire PECore_RunMac_if_and_112_cse;
  wire PECore_RunMac_if_and_113_cse;
  wire PECore_PushAxiRsp_if_and_cse;
  wire PECore_PushAxiRsp_if_and_10_cse;
  wire PECore_PushOutput_if_and_cse;
  reg reg_Datapath_for_1_ProductSum_cmp_cgo_ir_3_cse;
  reg reg_input_mem_banks_bank_array_impl_data0_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data15_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data14_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data13_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data12_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data11_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data10_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data9_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data8_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data7_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data6_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data5_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data4_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data3_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data2_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data1_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data0_rsci_cgo_ir_cse;
  reg reg_start_PopNB_mioi_iswt0_cse;
  reg reg_rva_out_Push_mioi_iswt0_cse;
  reg reg_act_port_Push_mioi_iswt0_cse;
  wire pe_manager_adplfloat_bias_weight_and_cse;
  wire pe_manager_adplfloat_bias_weight_and_1_cse;
  wire pe_manager_cluster_lut_data_and_cse;
  wire pe_manager_cluster_lut_data_and_1_cse;
  wire pe_config_num_output_and_cse;
  wire and_5345_cse;
  wire PECore_RunMac_if_and_12_cse;
  wire PECore_RunMac_if_and_13_cse;
  wire PECore_RunMac_if_and_10_cse;
  wire PECore_RunMac_if_and_11_cse;
  wire or_1405_cse;
  wire or_1409_cse;
  wire or_1413_cse;
  wire or_1417_cse;
  wire or_1421_cse;
  wire or_1425_cse;
  wire or_1429_cse;
  wire or_1433_cse;
  wire or_1437_cse;
  wire or_1441_cse;
  wire or_1445_cse;
  wire or_1449_cse;
  wire or_1453_cse;
  wire or_1457_cse;
  wire or_1461_cse;
  wire or_1465_cse;
  wire or_1183_cse;
  wire [127:0] input_mem_banks_write_if_for_if_mux_cse;
  wire or_500_cse;
  wire and_cse;
  wire and_3039_cse;
  wire and_3035_cse;
  wire and_3031_cse;
  wire and_3027_cse;
  wire and_3023_cse;
  wire and_3019_cse;
  wire and_3015_cse;
  wire and_3011_cse;
  wire and_3007_cse;
  wire and_3003_cse;
  wire and_2999_cse;
  wire and_2995_cse;
  wire and_2991_cse;
  wire and_2987_cse;
  wire and_2983_cse;
  wire and_2979_cse;
  wire nor_499_cse;
  wire and_5335_cse;
  wire or_55_cse;
  wire nand_199_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_450_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_452_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_453_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_454_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_455_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_456_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_457_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_420_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_422_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_423_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_424_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_425_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_426_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_427_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_390_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_392_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_393_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_394_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_395_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_396_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_397_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_360_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_362_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_363_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_364_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_365_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_366_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_367_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_330_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_332_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_333_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_334_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_335_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_336_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_337_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_300_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_302_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_303_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_304_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_305_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_306_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_307_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_270_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_272_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_273_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_274_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_275_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_276_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_277_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_240_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_242_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_243_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_244_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_245_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_246_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_247_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_210_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_212_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_213_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_214_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_215_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_216_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_217_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_180_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_182_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_183_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_184_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_185_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_186_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_187_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_150_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_152_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_153_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_154_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_155_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_156_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_157_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_120_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_122_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_123_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_124_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_125_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_126_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_127_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_90_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_92_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_93_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_94_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_95_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_96_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_97_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_60_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_62_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_63_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_64_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_65_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_66_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_67_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_30_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_32_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_33_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_34_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_35_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_36_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_37_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_2_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_3_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_4_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_5_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_6_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_7_cse;
  wire PECore_PushAxiRsp_if_and_45_cse;
  wire pe_config_is_valid_and_cse;
  wire or_1584_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_1_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_2_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_3_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_4_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_5_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_6_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_7_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_8_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_9_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_10_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_11_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_12_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_13_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_14_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_15_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_16_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire and_2973_cse;
  wire rva_out_reg_data_and_2_cse;
  wire [7:0] weight_write_data_data_mux1h_14_rmff;
  wire [7:0] weight_write_data_data_mux1h_13_rmff;
  wire [7:0] weight_write_data_data_mux1h_12_rmff;
  wire [7:0] weight_write_data_data_mux1h_11_rmff;
  wire [7:0] weight_write_data_data_mux1h_10_rmff;
  wire [7:0] weight_write_data_data_mux1h_9_rmff;
  wire [7:0] weight_write_data_data_mux1h_8_rmff;
  wire [7:0] weight_write_data_data_mux1h_7_rmff;
  wire [7:0] weight_write_data_data_mux1h_6_rmff;
  wire [7:0] weight_write_data_data_mux1h_5_rmff;
  wire [7:0] weight_write_data_data_mux1h_4_rmff;
  wire [7:0] weight_write_data_data_mux1h_3_rmff;
  wire [7:0] weight_write_data_data_mux1h_2_rmff;
  wire [7:0] weight_write_data_data_mux1h_1_rmff;
  wire [7:0] weight_write_data_data_mux1h_rmff;
  wire [127:0] input_mem_banks_read_read_data_mux_rmff;
  wire or_2419_rmff;
  wire or_2438_rmff;
  wire or_2437_rmff;
  wire or_2436_rmff;
  wire or_2435_rmff;
  wire or_2434_rmff;
  wire or_2433_rmff;
  wire or_2432_rmff;
  wire or_2431_rmff;
  wire or_2430_rmff;
  wire or_2429_rmff;
  wire or_2428_rmff;
  wire or_2427_rmff;
  wire or_2426_rmff;
  wire or_2425_rmff;
  wire or_2424_rmff;
  wire or_2423_rmff;
  wire or_2422_rmff;
  wire or_2421_rmff;
  reg [7:0] pe_config_output_counter_sva;
  reg [7:0] pe_manager_num_input_0_sva;
  reg [7:0] pe_manager_num_input_1_sva;
  reg [7:0] pe_config_input_counter_sva;
  reg [7:0] PECore_RunMac_if_mux_175_itm;
  reg [7:0] pe_manager_cluster_lut_data_0_0_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_1_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_2_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_3_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_4_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_5_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_6_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_7_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_8_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_9_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_10_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_11_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_12_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_13_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_14_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_15_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_0_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_1_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_2_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_3_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_4_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_5_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_6_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_7_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_8_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_9_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_10_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_11_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_12_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_13_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_14_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_15_sva_dfm_4;
  wire [7:0] weight_port_read_out_data_7_15_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_15_15_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_15_itm;
  reg [7:0] PECore_RunMac_if_mux_174_itm;
  reg [7:0] weight_port_read_out_data_15_14_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_173_itm;
  wire [7:0] weight_port_read_out_data_7_14_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_15_13_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_13_itm;
  reg [7:0] PECore_RunMac_if_mux_172_itm;
  reg [7:0] weight_port_read_out_data_15_12_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_13_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] rva_out_reg_data_79_72_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_171_itm;
  wire [7:0] weight_port_read_out_data_7_13_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_15_11_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_12_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_170_itm;
  reg [7:0] weight_port_read_out_data_15_10_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_11_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_169_itm;
  wire [7:0] weight_port_read_out_data_7_12_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_15_9_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_10_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_9_itm;
  reg [7:0] PECore_RunMac_if_mux_168_itm;
  reg [7:0] weight_port_read_out_data_15_8_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_9_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_8_itm;
  reg [7:0] PECore_RunMac_if_mux_167_itm;
  wire [7:0] weight_port_read_out_data_7_11_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_15_7_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_8_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_7_itm;
  reg [7:0] PECore_RunMac_if_mux_166_itm;
  reg [7:0] weight_port_read_out_data_15_6_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_7_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_6_itm;
  reg [7:0] PECore_RunMac_if_mux_165_itm;
  wire [7:0] weight_port_read_out_data_7_10_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_15_5_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_6_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_5_itm;
  reg [7:0] PECore_RunMac_if_mux_164_itm;
  reg [7:0] weight_port_read_out_data_15_4_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_5_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_4_itm;
  reg [7:0] PECore_RunMac_if_mux_163_itm;
  wire [7:0] weight_port_read_out_data_7_9_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_15_3_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_4_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_3_itm;
  reg [7:0] PECore_RunMac_if_mux_162_itm;
  reg [7:0] weight_port_read_out_data_15_2_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_3_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_2_itm;
  reg [7:0] PECore_RunMac_if_mux_161_itm;
  wire [7:0] weight_port_read_out_data_7_8_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_15_1_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_2_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_160_itm;
  reg [7:0] weight_port_read_out_data_15_0_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_1_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_itm;
  reg [7:0] PECore_RunMac_if_mux_95_itm;
  wire [7:0] weight_port_read_out_data_6_15_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_13_15_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_191_itm;
  reg [7:0] PECore_RunMac_if_mux_79_itm;
  reg [7:0] PECore_RunMac_if_mux_94_itm;
  reg [7:0] weight_port_read_out_data_13_14_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_190_itm;
  reg [7:0] PECore_RunMac_if_mux_78_itm;
  reg [7:0] PECore_RunMac_if_mux_93_itm;
  wire [7:0] weight_port_read_out_data_6_14_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_13_13_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_15;
  reg [7:0] PECore_RunMac_if_mux_189_itm;
  reg [7:0] PECore_RunMac_if_mux_77_itm;
  reg [7:0] PECore_RunMac_if_mux_92_itm;
  reg [7:0] weight_port_read_out_data_13_12_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_17;
  reg [7:0] PECore_RunMac_if_mux_188_itm;
  reg [7:0] PECore_RunMac_if_mux_76_itm;
  reg [7:0] PECore_RunMac_if_mux_91_itm;
  wire [7:0] weight_port_read_out_data_6_13_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_13_11_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_19;
  reg [7:0] PECore_RunMac_if_mux_187_itm;
  reg [7:0] PECore_RunMac_if_mux_75_itm;
  reg [7:0] PECore_RunMac_if_mux_90_itm;
  reg [7:0] weight_port_read_out_data_13_10_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_21;
  reg [7:0] PECore_RunMac_if_mux_186_itm;
  reg [7:0] PECore_RunMac_if_mux_74_itm;
  reg [7:0] PECore_RunMac_if_mux_89_itm;
  wire [7:0] weight_port_read_out_data_6_12_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_13_9_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_23;
  reg [7:0] PECore_RunMac_if_mux_185_itm;
  reg [7:0] PECore_RunMac_if_mux_73_itm;
  reg [7:0] PECore_RunMac_if_mux_88_itm;
  reg [7:0] weight_port_read_out_data_13_8_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_25;
  reg [7:0] PECore_RunMac_if_mux_184_itm;
  reg [7:0] PECore_RunMac_if_mux_72_itm;
  reg [7:0] PECore_RunMac_if_mux_87_itm;
  wire [7:0] weight_port_read_out_data_6_11_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_13_7_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_27;
  reg [7:0] PECore_RunMac_if_mux_183_itm;
  reg [7:0] PECore_RunMac_if_mux_71_itm;
  reg [7:0] PECore_RunMac_if_mux_86_itm;
  reg [7:0] weight_port_read_out_data_13_6_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_29;
  reg [7:0] PECore_RunMac_if_mux_182_itm;
  reg [7:0] PECore_RunMac_if_mux_70_itm;
  reg [7:0] PECore_RunMac_if_mux_85_itm;
  wire [7:0] weight_port_read_out_data_6_10_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_13_5_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_31;
  reg [7:0] PECore_RunMac_if_mux_181_itm;
  reg [7:0] PECore_RunMac_if_mux_69_itm;
  reg [7:0] PECore_RunMac_if_mux_84_itm;
  reg [7:0] weight_port_read_out_data_13_4_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_33;
  reg [7:0] PECore_RunMac_if_mux_180_itm;
  reg [7:0] PECore_RunMac_if_mux_68_itm;
  reg [7:0] PECore_RunMac_if_mux_83_itm;
  wire [7:0] weight_port_read_out_data_6_9_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_13_3_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_35;
  reg [7:0] PECore_RunMac_if_mux_179_itm;
  reg [7:0] PECore_RunMac_if_mux_67_itm;
  reg [7:0] PECore_RunMac_if_mux_82_itm;
  reg [7:0] weight_port_read_out_data_13_2_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_37;
  reg [7:0] PECore_RunMac_if_mux_178_itm;
  reg [7:0] PECore_RunMac_if_mux_66_itm;
  reg [7:0] PECore_RunMac_if_mux_81_itm;
  wire [7:0] weight_port_read_out_data_6_8_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_13_1_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_39;
  reg [7:0] PECore_RunMac_if_mux_177_itm;
  reg [7:0] PECore_RunMac_if_mux_65_itm;
  reg [7:0] PECore_RunMac_if_mux_80_itm;
  reg [7:0] weight_port_read_out_data_13_0_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_41;
  reg [7:0] PECore_RunMac_if_mux_176_itm;
  reg [7:0] PECore_RunMac_if_mux_64_itm;
  reg [7:0] PECore_RunMac_if_mux_111_itm;
  wire [7:0] weight_port_read_out_data_7_7_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_14_15_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_63_itm;
  reg [7:0] PECore_RunMac_if_mux_110_itm;
  reg [7:0] weight_port_read_out_data_14_14_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_62_itm;
  reg [7:0] PECore_RunMac_if_mux_109_itm;
  wire [7:0] weight_port_read_out_data_7_6_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_14_13_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_61_itm;
  reg [7:0] PECore_RunMac_if_mux_108_itm;
  reg [7:0] weight_port_read_out_data_14_12_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_13_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_60_itm;
  reg [7:0] PECore_RunMac_if_mux_107_itm;
  wire [7:0] weight_port_read_out_data_7_5_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_14_11_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_12_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_59_itm;
  reg [7:0] PECore_RunMac_if_mux_106_itm;
  reg [7:0] weight_port_read_out_data_14_10_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_11_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_58_itm;
  reg [7:0] PECore_RunMac_if_mux_105_itm;
  wire [7:0] weight_port_read_out_data_7_4_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_14_9_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_10_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_57_itm;
  reg [7:0] weight_port_read_out_data_14_8_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_9_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_136_itm;
  reg [7:0] PECore_RunMac_if_mux_56_itm;
  wire [7:0] weight_port_read_out_data_7_3_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_14_7_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_8_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_135_itm;
  reg [7:0] PECore_RunMac_if_mux_55_itm;
  reg [7:0] weight_port_read_out_data_14_6_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_7_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_134_itm;
  reg [7:0] PECore_RunMac_if_mux_54_itm;
  wire [7:0] weight_port_read_out_data_7_2_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_14_5_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_6_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_133_itm;
  reg [7:0] PECore_RunMac_if_mux_53_itm;
  reg [7:0] weight_port_read_out_data_14_4_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_5_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_132_itm;
  reg [7:0] PECore_RunMac_if_mux_52_itm;
  reg [7:0] PECore_RunMac_if_mux_99_itm;
  wire [7:0] weight_port_read_out_data_7_1_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_14_3_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_4_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_131_itm;
  reg [7:0] PECore_RunMac_if_mux_51_itm;
  reg [7:0] PECore_RunMac_if_mux_98_itm;
  reg [7:0] weight_port_read_out_data_14_2_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_3_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_130_itm;
  reg [7:0] PECore_RunMac_if_mux_50_itm;
  reg [7:0] PECore_RunMac_if_mux_97_itm;
  wire [7:0] weight_port_read_out_data_7_0_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_14_1_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_2_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_49_itm;
  reg [7:0] PECore_RunMac_if_mux_96_itm;
  reg [7:0] weight_port_read_out_data_14_0_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_1_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_48_itm;
  reg [7:0] PECore_RunMac_if_mux_159_itm;
  wire [7:0] weight_port_read_out_data_6_7_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_12_15_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1;
  reg [7:0] PECore_RunMac_if_mux_47_itm;
  reg [7:0] PECore_RunMac_if_mux_158_itm;
  reg [7:0] weight_port_read_out_data_12_14_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1;
  reg [7:0] PECore_RunMac_if_mux_46_itm;
  reg [7:0] PECore_RunMac_if_mux_157_itm;
  wire [7:0] weight_port_read_out_data_6_6_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_12_13_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1;
  reg [7:0] PECore_RunMac_if_mux_45_itm;
  reg [7:0] PECore_RunMac_if_mux_156_itm;
  reg [7:0] weight_port_read_out_data_12_12_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1;
  reg [7:0] PECore_RunMac_if_mux_44_itm;
  reg [7:0] PECore_RunMac_if_mux_155_itm;
  wire [7:0] weight_port_read_out_data_6_5_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_12_11_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1;
  reg [7:0] PECore_RunMac_if_mux_43_itm;
  reg [7:0] PECore_RunMac_if_mux_154_itm;
  reg [7:0] weight_port_read_out_data_12_10_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1;
  reg [7:0] PECore_RunMac_if_mux_42_itm;
  reg [7:0] PECore_RunMac_if_mux_153_itm;
  wire [7:0] weight_port_read_out_data_6_4_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_12_9_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1;
  reg [7:0] rva_out_reg_data_95_88_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_41_itm;
  reg [7:0] PECore_RunMac_if_mux_152_itm;
  reg [7:0] weight_port_read_out_data_12_8_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1;
  reg [7:0] rva_out_reg_data_87_80_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_40_itm;
  reg [7:0] PECore_RunMac_if_mux_151_itm;
  wire [7:0] weight_port_read_out_data_6_3_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_12_7_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1;
  reg [7:0] rva_out_reg_data_71_64_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_39_itm;
  reg [7:0] PECore_RunMac_if_mux_150_itm;
  reg [7:0] weight_port_read_out_data_12_6_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1;
  reg [7:0] rva_out_reg_data_63_56_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_38_itm;
  reg [7:0] PECore_RunMac_if_mux_149_itm;
  wire [7:0] weight_port_read_out_data_6_2_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_12_5_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_37_itm;
  reg [7:0] PECore_RunMac_if_mux_148_itm;
  reg [7:0] weight_port_read_out_data_12_4_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1;
  reg [7:0] rva_out_reg_data_47_40_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_36_itm;
  reg [7:0] PECore_RunMac_if_mux_147_itm;
  wire [7:0] weight_port_read_out_data_6_1_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_12_3_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1;
  reg [7:0] rva_out_reg_data_127_120_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_35_itm;
  reg [7:0] PECore_RunMac_if_mux_146_itm;
  reg [7:0] weight_port_read_out_data_12_2_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1;
  reg [7:0] rva_out_reg_data_119_112_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_34_itm;
  reg [7:0] PECore_RunMac_if_mux_145_itm;
  wire [7:0] weight_port_read_out_data_6_0_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_12_1_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1;
  reg [7:0] rva_out_reg_data_111_104_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_33_itm;
  reg [7:0] PECore_RunMac_if_mux_144_itm;
  reg [7:0] weight_port_read_out_data_12_0_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1;
  reg [7:0] rva_out_reg_data_103_96_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_32_itm;
  wire while_and_127_cse_1;
  wire [11:0] weight_read_addrs_0_15_4_lpi_1_dfm_5_mx0;
  wire [15:0] weight_read_addrs_1_lpi_1_dfm_2;
  wire [14:0] weight_read_addrs_2_15_1_lpi_1_dfm_2;
  wire [15:0] weight_read_addrs_3_lpi_1_dfm_2;
  wire [13:0] weight_read_addrs_4_15_2_lpi_1_dfm_2;
  wire [15:0] weight_read_addrs_5_lpi_1_dfm_2;
  wire [14:0] weight_read_addrs_6_15_1_lpi_1_dfm_2;
  wire [15:0] weight_read_addrs_7_lpi_1_dfm_2;
  wire [12:0] weight_read_addrs_8_15_3_lpi_1_dfm_3;
  wire [15:0] weight_read_addrs_9_lpi_1_dfm_3;
  wire [14:0] weight_read_addrs_10_15_1_lpi_1_dfm_3;
  wire [15:0] weight_read_addrs_11_lpi_1_dfm_3;
  wire [13:0] weight_read_addrs_12_15_2_lpi_1_dfm_3;
  wire [15:0] weight_read_addrs_13_lpi_1_dfm_3;
  wire [14:0] weight_read_addrs_14_15_1_lpi_1_dfm_3;
  wire [15:0] weight_read_addrs_15_lpi_1_dfm_3;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_3_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_3_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_3_0_sva_1;
  wire [15:0] weight_write_addrs_lpi_1_dfm_6;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_4_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_4_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_4_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_5_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_5_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_5_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_6_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_6_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_6_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_7_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_7_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_7_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_8_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_8_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_8_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_9_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_9_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_9_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_10_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_10_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_10_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_11_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_11_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_11_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_12_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_12_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_12_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_13_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_13_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_13_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_14_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_14_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_14_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_15_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_15_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_15_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_16_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_16_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_16_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_17_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_17_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_17_0_sva_1;
  reg [15:0] pe_manager_base_input_0_sva;
  reg [15:0] pe_manager_base_input_1_sva;
  reg [15:0] pe_manager_base_bias_0_sva;
  reg [15:0] pe_manager_base_bias_1_sva;
  wire or_dcpl_717;
  wire or_dcpl_718;
  wire or_dcpl_724;
  reg [31:0] PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_11_sva;
  reg [31:0] PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_1_sva;
  reg [31:0] PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_5_sva;
  reg [31:0] PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_4_sva;
  wire PECore_DecodeAxiRead_switch_lp_nor_10_cse_1;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_5;
  reg [7:0] weight_port_read_out_data_0_0_sva_dfm;
  reg [31:0] accum_vector_data_4_sva;
  reg [31:0] accum_vector_data_3_sva;
  reg [31:0] accum_vector_data_2_sva;
  reg [19:0] act_port_reg_data_10_sva;
  reg [19:0] act_port_reg_data_9_sva;
  reg [19:0] act_port_reg_data_6_sva;
  reg [19:0] act_port_reg_data_5_sva;
  reg [31:0] accum_vector_data_9_sva;
  reg [31:0] accum_vector_data_6_sva;
  reg [31:0] accum_vector_data_5_sva;
  reg [31:0] PECore_RunBias_if_accum_vector_out_data_14_lpi_1_dfm;
  reg [31:0] PECore_RunBias_if_accum_vector_out_data_15_lpi_1_dfm;
  wire and_tmp;
  wire PECore_PushAxiRsp_if_asn_70;
  wire and_5501_cse;
  wire and_5502_cse;
  wire or_1593_cse;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_or_6_cse_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_6_sva_1;
  wire [7:0] while_while_and_18_itm;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_15;
  wire [4:0] z_out_4;
  wire [5:0] nl_z_out_4;
  wire [7:0] z_out_5;
  wire [8:0] nl_z_out_5;
  wire [19:0] z_out_17;
  wire [20:0] nl_z_out_17;
  wire [19:0] z_out_18;
  wire [20:0] nl_z_out_18;
  wire [19:0] z_out_19;
  wire [20:0] nl_z_out_19;
  wire [19:0] z_out_20;
  wire [20:0] nl_z_out_20;
  wire [31:0] z_out_25;
  wire [32:0] nl_z_out_25;
  wire [31:0] z_out_26;
  wire [32:0] nl_z_out_26;
  wire [31:0] z_out_27;
  wire [32:0] nl_z_out_27;
  wire [31:0] z_out_28;
  wire [32:0] nl_z_out_28;
  wire [31:0] z_out_29;
  wire [32:0] nl_z_out_29;
  wire [31:0] z_out_30;
  wire [32:0] nl_z_out_30;
  wire [31:0] z_out_31;
  wire [32:0] nl_z_out_31;
  wire [31:0] z_out_32;
  wire [32:0] nl_z_out_32;
  wire [31:0] z_out_37;
  wire [31:0] z_out_38;
  wire [31:0] z_out_39;
  wire [31:0] z_out_40;
  wire or_tmp_3038;
  wire [7:0] z_out_41;
  wire [19:0] z_out_43;
  wire [19:0] z_out_44;
  wire [19:0] z_out_45;
  wire [19:0] z_out_46;
  wire [19:0] z_out_47;
  wire [19:0] z_out_48;
  wire [19:0] z_out_49;
  wire [3:0] z_out_50;
  wire [4:0] nl_z_out_50;
  reg weight_mem_read_arbxbar_arbiters_next_7_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_1_sva;
  reg [2:0] pe_manager_adplfloat_bias_weight_0_sva;
  reg [2:0] pe_manager_adplfloat_bias_weight_1_sva;
  reg [2:0] pe_manager_adplfloat_bias_bias_0_sva;
  reg [2:0] pe_manager_adplfloat_bias_bias_1_sva;
  reg [2:0] pe_manager_adplfloat_bias_input_0_sva;
  reg [2:0] pe_manager_adplfloat_bias_input_1_sva;
  reg [15:0] pe_manager_base_weight_0_sva;
  reg [15:0] pe_manager_base_weight_1_sva;
  reg [3:0] pe_config_num_manager_sva;
  reg [7:0] pe_config_num_output_sva;
  reg [31:0] accum_vector_data_7_sva;
  reg [31:0] accum_vector_data_8_sva;
  reg [31:0] accum_vector_data_12_sva;
  reg [31:0] accum_vector_data_13_sva;
  reg [31:0] accum_vector_data_14_sva;
  reg [31:0] accum_vector_data_15_sva;
  reg [19:0] act_port_reg_data_7_sva;
  reg [19:0] act_port_reg_data_8_sva;
  reg [19:0] act_port_reg_data_4_sva;
  reg [19:0] act_port_reg_data_11_sva;
  reg [19:0] act_port_reg_data_3_sva;
  reg [19:0] act_port_reg_data_12_sva;
  reg [19:0] act_port_reg_data_2_sva;
  reg [19:0] act_port_reg_data_13_sva;
  reg [19:0] act_port_reg_data_1_sva;
  reg [19:0] act_port_reg_data_14_sva;
  reg [19:0] act_port_reg_data_0_sva;
  reg [19:0] act_port_reg_data_15_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm;
  reg [7:0] weight_port_read_out_data_0_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_15_sva_dfm;
  reg PECore_RunBias_if_for_1_operator_32_true_slc_operator_32_true_acc_13_svs;
  reg PECore_RunBias_if_for_2_operator_32_true_slc_operator_32_true_acc_13_svs;
  reg PECore_RunBias_if_for_12_operator_32_true_slc_operator_32_true_acc_13_svs;
  reg [31:0] PECore_RunBias_if_accum_vector_out_data_13_lpi_1_dfm;
  reg [31:0] PECore_RunBias_if_accum_vector_out_data_lpi_1_dfm;
  reg PECore_DecodeAxiRead_case_4_switch_lp_and_itm;
  reg PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm;
  reg PECore_DecodeAxiRead_case_4_switch_lp_and_5_itm;
  reg [7:0] PECore_RunMac_if_mux_31_itm;
  reg [7:0] PECore_RunMac_if_mux_30_itm;
  reg [7:0] PECore_RunMac_if_mux_29_itm;
  reg [7:0] PECore_RunMac_if_mux_28_itm;
  reg [7:0] PECore_RunMac_if_mux_27_itm;
  reg [7:0] PECore_RunMac_if_mux_26_itm;
  reg [7:0] PECore_RunMac_if_mux_25_itm;
  reg [7:0] PECore_RunMac_if_mux_24_itm;
  reg [7:0] PECore_RunMac_if_mux_23_itm;
  reg [7:0] PECore_RunMac_if_mux_22_itm;
  reg [7:0] PECore_RunMac_if_mux_21_itm;
  reg [7:0] PECore_RunMac_if_mux_20_itm;
  reg [7:0] PECore_RunMac_if_mux_19_itm;
  reg [7:0] PECore_RunMac_if_mux_18_itm;
  reg [7:0] PECore_RunMac_if_mux_17_itm;
  reg [7:0] PECore_RunMac_if_mux_16_itm;
  reg PECore_RunBias_if_for_6_operator_4_false_slc_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_0_itm;
  reg PECore_RunBias_if_for_7_operator_4_false_slc_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_0_itm;
  reg PECore_RunBias_if_for_10_operator_4_false_slc_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_0_itm;
  reg PECore_RunBias_if_for_11_operator_4_false_slc_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_0_itm;
  reg [19:0] act_port_reg_data_asn_itm;
  reg [19:0] act_port_reg_data_asn_1_itm;
  reg [19:0] act_port_reg_data_asn_2_itm;
  reg [19:0] act_port_reg_data_asn_3_itm;
  reg pe_manager_cluster_lut_data_1_0_sva_0;
  reg pe_manager_cluster_lut_data_1_1_sva_0;
  reg pe_manager_cluster_lut_data_1_2_sva_0;
  reg pe_manager_cluster_lut_data_1_3_sva_0;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  wire [7:0] weight_port_read_out_data_5_8_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_9_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_10_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_11_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_12_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_13_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_14_sva_dfm_mx1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  wire [7:0] weight_port_read_out_data_5_15_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_0_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_1_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_2_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_3_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_4_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_5_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_6_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_7_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_8_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_9_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_10_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_11_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_12_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_13_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_14_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_15_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_8_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_9_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_10_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_11_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_12_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_13_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_14_sva_dfm_mx1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  wire [7:0] weight_port_read_out_data_3_15_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_0_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_1_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_2_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_3_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_4_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_5_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_6_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_7_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_0_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_1_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_2_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_3_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_4_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_5_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_6_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_7_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_8_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_9_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_10_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_11_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_12_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_13_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_14_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_15_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_8_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_9_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_10_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_11_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_12_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_13_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_14_sva_dfm_mx1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  wire [7:0] weight_port_read_out_data_1_15_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_0_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_1_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_2_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_3_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_4_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_5_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_6_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_7_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_8_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_9_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_10_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_11_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_12_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_13_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_14_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_15_sva_dfm_mx1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_1_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  wire [7:0] weight_port_read_out_data_0_0_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_1_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_2_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_3_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_4_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_5_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_6_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_7_sva_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm_mx1;
  wire adpfloat_tmp_is_zero_land_11_lpi_1_dfm_mx1w0;
  wire adpfloat_tmp_is_zero_land_10_lpi_1_dfm_mx1w0;
  wire adpfloat_tmp_is_zero_land_7_lpi_1_dfm_mx1w0;
  wire adpfloat_tmp_is_zero_land_6_lpi_1_dfm_mx1w0;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  wire [7:0] weight_port_read_out_data_5_0_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_1_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_2_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_3_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_4_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_5_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_6_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_7_sva_dfm_mx1;
  wire while_and_32_cse_1;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm_1;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm_1;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm_1;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm_1;
  wire input_read_req_valid_lpi_1_dfm_6;
  wire PECore_DecodeAxiRead_switch_lp_nor_2_itm_mx0w0;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_13_cse_1;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_12_cse_1;
  wire PECore_DecodeAxiRead_switch_lp_nor_14_cse_1;
  wire [12:0] PEManager_16U_GetWeightAddr_if_acc_2_psp_sva_1;
  wire [13:0] nl_PEManager_16U_GetWeightAddr_if_acc_2_psp_sva_1;
  wire [15:0] PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx1;
  wire [11:0] PEManager_16U_GetWeightAddr_1_else_acc_2_psp_sva_1;
  wire [12:0] nl_PEManager_16U_GetWeightAddr_1_else_acc_2_psp_sva_1;
  wire [2:0] weight_read_addrs_8_2_0_lpi_1_dfm_1;
  wire [3:0] while_asn_294_mx0w0;
  wire [3:0] pe_config_manager_counter_sva_dfm_4_mx1;
  wire [7:0] pe_config_input_counter_sva_dfm_4_mx0;
  wire [7:0] pe_config_output_counter_sva_dfm_4_mx0;
  wire [1:0] weight_read_addrs_4_1_0_lpi_1_dfm_1;
  wire weight_read_addrs_0_2_0_lpi_1_dfm_4_2_mx0;
  wire weight_read_addrs_0_2_0_lpi_1_dfm_4_1_mx0;
  wire weight_read_addrs_0_2_0_lpi_1_dfm_4_0_mx0;
  wire weight_read_addrs_0_3_lpi_1_dfm_6;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_14_sva_1;
  wire weight_read_addrs_0_3_lpi_1_dfm_5_mx0;
  wire weight_mem_run_1_if_for_land_1_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_2_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_3_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_4_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_5_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_6_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_7_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_8_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_9_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_10_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_11_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_12_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_13_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_14_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_15_lpi_1_dfm_1;
  wire weight_read_req_valid_0_lpi_1_dfm_4_mx0;
  wire Arbiter_16U_Roundrobin_pick_return_0_1_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_2_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_3_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_4_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_5_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_6_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_7_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_8_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_9_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_10_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_11_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_12_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_13_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_14_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_15_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_lpi_1_dfm_2;
  wire input_write_req_valid_lpi_1_dfm_6;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_1_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_1_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_1_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_1_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_1_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_1_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_1_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_1_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_2_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_2_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_2_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_2_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_2_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_2_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_2_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_2_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_3_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_3_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_3_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_3_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_3_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_3_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_3_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_3_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_4_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_4_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_4_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_4_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_4_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_4_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_4_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_4_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_5_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_5_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_5_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_5_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_5_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_5_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_5_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_5_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_6_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_6_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_6_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_6_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_6_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_6_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_6_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_7_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_7_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_7_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_7_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_7_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_7_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_7_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_7_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_8_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_8_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_8_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_8_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_8_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_8_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_8_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_8_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_8_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_8_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_8_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_9_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_9_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_9_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_9_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_9_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_9_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_9_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_9_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_9_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_9_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_9_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_10_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_10_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_10_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_10_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_10_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_10_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_10_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_10_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_10_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_10_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_10_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_11_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_11_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_11_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_11_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_11_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_11_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_11_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_11_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_11_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_11_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_11_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_12_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_12_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_12_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_12_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_12_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_12_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_12_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_12_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_12_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_12_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_12_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_13_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_13_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_13_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_13_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_13_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_13_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_13_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_13_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_13_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_13_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_13_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_14_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_14_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_14_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_14_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_14_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_14_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_14_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_14_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_14_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_14_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_14_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_15_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_15_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_15_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_15_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_15_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_15_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_15_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_15_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_15_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_15_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_15_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_sva_1;
  wire [3:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_lpi_1_dfm_1;
  wire [3:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_14_lpi_1_dfm_1;
  wire [1:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_13_3_2_lpi_1_dfm_1;
  wire [1:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_13_1_0_lpi_1_dfm_1;
  wire [3:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_12_lpi_1_dfm_1;
  wire [2:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_3_1_lpi_1_dfm_1;
  wire [2:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_2_0_lpi_1_dfm_1;
  wire [3:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_8_lpi_1_dfm_1;
  wire [2:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_3_1_lpi_1_dfm_1;
  wire [3:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_6_lpi_1_dfm_1;
  wire [1:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_5_3_2_lpi_1_dfm_1;
  wire [1:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_5_1_0_lpi_1_dfm_1;
  wire [3:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_4_lpi_1_dfm_1;
  wire [2:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_3_1_lpi_1_dfm_1;
  wire [3:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_2_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_14_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_14_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_14_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_14_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_14_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_14_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_14_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_14_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_14_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_14_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_14_sva_1;
  wire pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_pe_config_UpdateInputCounter_if_nor_svs_1;
  wire PECore_UpdateFSM_switch_lp_unequal_tmp_1;
  wire weight_read_req_valid_8_lpi_1_dfm_1;
  wire weight_read_addrs_10_0_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire [3:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_10_lpi_1_dfm_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_241;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_243;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_245;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_247;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_249;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_251;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_253;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_255;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_257;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_259;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_261;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_263;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_265;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_267;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_269;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_271;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_1_sva_mx0w2;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_1_sva_mx0w2;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_12_sva_mx0w1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_12_sva_mx0w1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_2_sva_mx0w1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_2_sva_mx0w1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_3_sva_mx0w1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_3_sva_mx0w1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_4_sva_mx0w1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_4_sva_mx0w1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_5_sva_mx0w1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_5_sva_mx0w1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_8_sva_mx0w1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_8_sva_mx0w1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_9_sva_mx0w1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_9_sva_mx0w1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_12_mx1w2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_11_mx1w2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_13_mx1w2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_0_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_1_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_2_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_3_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_4_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_5_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_6_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_7_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_8_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_9_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_10_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_11_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_12_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_13_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_14_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_15_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_15_lpi_1_dfm_3;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1;
  wire [3:0] operator_4_false_acc_psp_1_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_1_sva_1;
  wire [3:0] operator_4_false_acc_psp_2_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_2_sva_1;
  wire [3:0] operator_4_false_acc_psp_3_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_3_sva_1;
  wire [3:0] operator_4_false_acc_psp_4_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_4_sva_1;
  wire [3:0] operator_4_false_acc_psp_5_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_5_sva_1;
  wire [3:0] operator_4_false_acc_psp_8_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_8_sva_1;
  wire [3:0] operator_4_false_acc_psp_9_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_9_sva_1;
  wire [3:0] operator_4_false_acc_psp_12_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_12_sva_1;
  wire [3:0] operator_4_false_acc_psp_13_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_13_sva_1;
  wire [3:0] operator_4_false_acc_psp_14_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_14_sva_1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_14_sva_1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_14_sva_1;
  wire [3:0] operator_4_false_acc_psp_15_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_15_sva_1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_15_sva_1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_15_sva_1;
  wire [3:0] operator_4_false_acc_psp_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_sva_1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_sva_1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_sva_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_6_sva_1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_6_sva_1;
  wire [3:0] operator_4_false_acc_psp_6_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_6_sva_1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_7_sva_1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_7_sva_1;
  wire [3:0] operator_4_false_acc_psp_7_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_7_sva_1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_10_sva_1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_10_sva_1;
  wire [3:0] operator_4_false_acc_psp_10_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_10_sva_1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_11_sva_1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_11_sva_1;
  wire [3:0] operator_4_false_acc_psp_11_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_11_sva_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44;
  wire [2:0] PECore_RunBias_if_for_if_bias_tmp2_mux_17;
  wire PECore_PushAxiRsp_if_asn_66;
  wire PECore_PushAxiRsp_if_asn_68;
  wire [3:0] PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx0_3_0;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1_3;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1_2;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1_1;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1_0;
  wire [2:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_15_lpi_1_dfm_1_3_1;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_15_lpi_1_dfm_1_0;
  reg [7:0] reg_Datapath_for_conc_4_ftd;
  reg [7:0] reg_Datapath_for_conc_4_ftd_1;
  reg [7:0] reg_Datapath_for_conc_4_ftd_2;
  reg [7:0] reg_Datapath_for_conc_4_ftd_3;
  reg [7:0] reg_Datapath_for_conc_4_ftd_4;
  reg [7:0] reg_Datapath_for_conc_4_ftd_5;
  reg [7:0] reg_Datapath_for_conc_4_ftd_6;
  reg [7:0] reg_Datapath_for_conc_4_ftd_7;
  reg [7:0] reg_Datapath_for_conc_4_ftd_8;
  reg [7:0] reg_Datapath_for_conc_4_ftd_9;
  reg [7:0] reg_Datapath_for_conc_4_ftd_10;
  reg [7:0] reg_Datapath_for_conc_4_ftd_11;
  reg [7:0] reg_Datapath_for_conc_4_ftd_12;
  reg [7:0] reg_Datapath_for_conc_4_ftd_13;
  reg [7:0] reg_Datapath_for_conc_4_ftd_14;
  reg [7:0] reg_Datapath_for_conc_4_ftd_15;
  reg reg_PECore_RunMac_if_mux_143_ftd;
  reg [6:0] reg_PECore_RunMac_if_mux_143_ftd_1;
  reg [3:0] reg_PECore_RunMac_if_mux_142_ftd;
  reg [3:0] reg_PECore_RunMac_if_mux_142_ftd_1;
  reg [2:0] reg_PECore_RunMac_if_mux_141_ftd;
  reg [4:0] reg_PECore_RunMac_if_mux_141_ftd_1;
  reg [5:0] reg_PECore_RunMac_if_mux_140_ftd;
  reg [1:0] reg_PECore_RunMac_if_mux_140_ftd_1;
  reg [2:0] reg_PECore_RunMac_if_mux_14_ftd;
  reg [4:0] reg_PECore_RunMac_if_mux_14_ftd_1;
  reg [5:0] reg_PECore_RunMac_if_mux_139_ftd;
  reg [1:0] reg_PECore_RunMac_if_mux_139_ftd_1;
  reg [2:0] reg_PECore_RunMac_if_mux_138_ftd;
  reg [4:0] reg_PECore_RunMac_if_mux_138_ftd_1;
  reg [5:0] reg_PECore_RunMac_if_mux_137_ftd;
  reg [1:0] reg_PECore_RunMac_if_mux_137_ftd_1;
  reg [3:0] reg_PECore_RunMac_if_mux_129_ftd;
  reg [3:0] reg_PECore_RunMac_if_mux_129_ftd_1;
  reg [3:0] reg_PECore_RunMac_if_mux_128_ftd;
  reg [3:0] reg_PECore_RunMac_if_mux_128_ftd_1;
  reg [3:0] reg_PECore_RunMac_if_mux_127_ftd;
  reg [3:0] reg_PECore_RunMac_if_mux_127_ftd_1;
  reg [3:0] reg_PECore_RunMac_if_mux_126_ftd;
  reg [3:0] reg_PECore_RunMac_if_mux_126_ftd_1;
  reg [3:0] reg_PECore_RunMac_if_mux_125_ftd;
  reg [3:0] reg_PECore_RunMac_if_mux_125_ftd_1;
  reg [3:0] reg_PECore_RunMac_if_mux_124_ftd;
  reg [3:0] reg_PECore_RunMac_if_mux_124_ftd_1;
  reg [3:0] reg_PECore_RunMac_if_mux_123_ftd;
  reg [3:0] reg_PECore_RunMac_if_mux_123_ftd_1;
  reg [3:0] reg_PECore_RunMac_if_mux_11_ftd;
  reg [3:0] reg_PECore_RunMac_if_mux_11_ftd_1;
  reg [3:0] reg_PECore_RunMac_if_mux_122_ftd;
  reg [3:0] reg_PECore_RunMac_if_mux_122_ftd_1;
  wire PECore_RunBias_if_for_or_m1c_5;
  wire and_4031_m1c;
  wire PECore_RunMac_if_or_5_m1c;
  wire PECore_DecodeAxiRead_switch_lp_and_3_rgt;
  wire operator_32_true_and_6_rgt;
  wire PECore_RunBias_if_for_and_50_rgt;
  wire operator_32_true_and_2_rgt;
  wire PECore_RunMac_if_nand_56_rgt;
  wire PECore_RunMac_if_and_674_rgt;
  wire PECore_RunMac_if_and_675_rgt;
  wire PECore_RunMac_if_and_676_rgt;
  wire PECore_RunMac_if_and_627_rgt;
  wire PECore_RunMac_if_and_628_rgt;
  wire PECore_RunMac_if_and_580_rgt;
  wire PECore_RunMac_if_and_569_rgt;
  wire PECore_RunMac_if_and_570_rgt;
  wire PECore_RunMac_if_and_571_rgt;
  wire PECore_RunBias_if_for_and_45_rgt;
  wire PECore_RunBias_if_for_and_34_rgt;
  wire rva_out_reg_data_and_87_rgt;
  wire rva_out_reg_data_and_88_rgt;
  wire PECore_RunMac_if_and_346_rgt;
  reg reg_PECore_RunMac_asn_15_itm_1_ftd;
  reg reg_PECore_RunMac_asn_15_itm_1_ftd_1;
  reg reg_PECore_RunMac_asn_15_itm_1_ftd_2;
  wire PECore_RunMac_if_and_721_ssc;
  reg [2:0] reg_PECore_RunMac_if_mux_100_ftd;
  reg [4:0] reg_PECore_RunMac_if_mux_100_ftd_1;
  reg [2:0] reg_PECore_RunMac_if_mux_101_ftd;
  reg [4:0] reg_PECore_RunMac_if_mux_101_ftd_1;
  wire PECore_RunMac_if_and_723_ssc;
  reg [2:0] reg_PECore_RunMac_if_mux_102_ftd;
  reg [4:0] reg_PECore_RunMac_if_mux_102_ftd_1;
  reg [2:0] reg_PECore_RunMac_if_mux_103_ftd;
  reg [4:0] reg_PECore_RunMac_if_mux_103_ftd_1;
  reg [2:0] reg_PECore_RunMac_if_mux_104_ftd;
  reg [4:0] reg_PECore_RunMac_if_mux_104_ftd_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_1_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_2_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_3_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_4_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_5_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_6_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_7_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_8_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_9_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_10_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_11_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_12_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_13_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_14_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_0;
  wire weight_mem_read_arbxbar_xbar_for_3_1_operator_31_false_operator_31_false_operator_31_false_or_seb;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_1_lpi_1_dfm_3_0;
  wire weight_mem_read_arbxbar_xbar_for_3_2_operator_31_false_operator_31_false_operator_31_false_or_seb;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_2_lpi_1_dfm_3_0;
  wire weight_mem_read_arbxbar_xbar_for_3_3_operator_31_false_operator_31_false_operator_31_false_or_seb;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_3_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_4_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_5_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_6_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_7_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_8_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_9_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_10_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_11_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_12_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_13_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_14_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_15_lpi_1_dfm_3_0;
  wire is_start_and_cse;
  wire [31:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_15_cse;
  wire [31:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_14_cse;
  wire [19:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_25_cse;
  wire [19:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_26_cse;
  wire [19:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_21_cse;
  wire [19:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_22_cse;
  wire pe_config_manager_counter_and_cse;
  wire [31:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_2_cse;
  wire [31:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_3_cse;
  wire [31:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_4_cse;
  wire [31:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_12_cse;
  wire [31:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_1_cse;
  wire [31:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_13_cse;
  wire PECore_RunMac_if_and_572_cse;
  wire PECore_RunMac_if_and_cse;
  wire [31:0] PECore_RunBias_if_accum_vector_out_data_mux_5_cse;
  wire [31:0] PECore_RunBias_if_accum_vector_out_data_mux_9_cse;
  wire [31:0] PECore_RunBias_if_accum_vector_out_data_mux_11_cse;
  wire [31:0] PECore_RunBias_if_accum_vector_out_data_mux_7_cse;
  wire PECore_RunMac_if_and_434_cse;
  wire PECore_RunMac_if_and_433_cse;
  wire and_5541_cse;
  wire or_796_cse;
  wire or_3399_cse;
  wire PECore_RunMac_if_and_470_cse;
  wire PECore_RunMac_if_and_444_cse;
  wire PECore_RunMac_if_and_445_cse;
  wire PECore_RunMac_if_and_398_cse;
  wire PECore_RunMac_if_and_399_cse;
  wire PECore_RunMac_if_and_390_cse;
  wire PECore_RunMac_if_and_391_cse;
  wire while_and_74_cse;
  wire while_and_66_cse;
  reg [2:0] reg_PECore_RunMac_if_mux_10_ftd;
  reg [4:0] reg_PECore_RunMac_if_mux_10_ftd_1;
  reg [2:0] reg_PECore_RunMac_if_mux_1_ftd;
  reg [4:0] reg_PECore_RunMac_if_mux_1_ftd_1;
  wire PECore_RunMac_if_or_140_m1c;
  wire PECore_RunMac_if_or_143_m1c;
  wire PECore_RunMac_if_or_145_m1c;
  wire PECore_RunBias_if_accum_vector_out_data_and_15_rgt;
  wire PECore_RunMac_if_and_817_rgt;
  wire PECore_RunMac_if_and_472_rgt;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_2;
  wire accum_vector_data_and_6_cse;
  wire act_port_reg_data_and_8_cse;
  wire weight_port_read_out_data_and_cse;
  wire weight_port_read_out_data_and_16_cse;
  wire weight_port_read_out_data_and_32_cse;
  wire weight_port_read_out_data_and_48_cse;
  wire weight_port_read_out_data_and_64_cse;
  wire weight_port_read_out_data_and_80_cse;
  wire weight_port_read_out_data_and_96_cse;
  wire weight_port_read_out_data_and_112_cse;
  wire weight_port_read_out_data_and_128_cse;
  wire weight_port_read_out_data_and_136_cse;
  wire weight_port_read_out_data_and_152_cse;
  wire weight_port_read_out_data_and_168_cse;
  wire weight_port_read_out_data_and_184_cse;
  wire weight_port_read_out_data_and_200_cse;
  wire accum_vector_data_and_9_cse;
  wire PECore_DecodeAxi_if_and_3_cse;
  wire or_1534_cse;
  wire PECore_CheckStart_start_reg_and_cse;
  wire operator_4_false_and_cse;
  wire adpfloat_tmp_is_zero_aelse_and_cse;
  wire operator_32_true_and_12_cse;
  wire weight_port_read_out_data_and_216_cse;
  wire weight_port_read_out_data_and_232_cse;
  wire adpfloat_tmp_is_zero_aelse_and_4_cse;
  wire accum_vector_data_and_15_cse;
  wire adpfloat_tmp_is_zero_aelse_and_6_cse;
  wire PECore_RunMac_if_and_685_cse;
  wire PECore_RunMac_if_and_701_cse;
  wire PECore_RunMac_if_and_717_cse;
  wire PECore_RunMac_if_and_726_cse;
  wire while_and_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_2_cse;
  wire PECore_RunBias_if_for_and_47_cse;
  wire PECore_RunBias_if_for_and_48_cse;
  wire and_2966_cse;
  wire act_port_reg_data_and_24_cse;
  wire rva_out_reg_data_and_91_cse;
  wire pe_config_UpdateInputCounter_if_and_cse;
  wire PECore_RunBias_if_for_and_42_cse;
  wire or_1521_cse;
  wire PECore_RunBias_if_for_and_cse;
  wire PECore_RunMac_if_and_359_cse;
  wire PECore_RunMac_if_and_360_cse;
  wire PECore_RunMac_if_and_361_cse;
  wire PECore_RunMac_if_and_834_rgt;
  wire PECore_RunMac_if_and_820_rgt;
  wire PECore_RunMac_if_and_430_cse;
  wire PECore_RunMac_if_and_431_cse;
  wire PECore_RunBias_if_accum_vector_out_data_and_17_cse;
  wire PECore_RunMac_if_and_859_cse;
  wire PECore_RunMac_if_and_867_cse;
  wire PECore_RunMac_if_and_872_cse;
  wire pe_config_UpdateManagerCounter_if_unequal_tmp;
  wire and_5872_cse;
  wire and_5844_cse;
  wire and_5871_cse;
  reg reg_PECore_RunMac_if_mux_123_1_enexo;
  reg reg_PECore_RunMac_if_mux_142_1_enexo;
  reg reg_rva_out_reg_data_47_40_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_63_56_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_71_64_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_79_72_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_87_80_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_95_88_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_103_96_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_111_104_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_119_112_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_127_120_sva_dfm_4_enexo;
  reg reg_act_port_reg_data_0_enexo;
  reg reg_act_port_reg_data_1_enexo;
  reg reg_act_port_reg_data_2_enexo;
  reg reg_act_port_reg_data_3_enexo;
  reg reg_act_port_reg_data_4_enexo;
  reg reg_act_port_reg_data_5_enexo;
  reg reg_act_port_reg_data_6_enexo;
  reg reg_act_port_reg_data_9_enexo;
  reg reg_act_port_reg_data_10_enexo;
  reg reg_act_port_reg_data_asn_3_enexo;
  reg reg_act_port_reg_data_asn_2_enexo;
  reg reg_act_port_reg_data_asn_1_enexo;
  reg reg_act_port_reg_data_asn_enexo;
  reg reg_act_port_reg_data_14_enexo;
  reg reg_act_port_reg_data_13_enexo;
  reg reg_act_port_reg_data_12_enexo;
  reg reg_act_port_reg_data_15_enexo;
  reg reg_PECore_RunMac_if_mux_31_enexo;
  wire PECore_PushAxiRsp_if_and_47_enex5;
  wire PECore_PushAxiRsp_if_and_48_enex5;
  wire PECore_PushAxiRsp_if_and_49_enex5;
  wire PECore_PushAxiRsp_if_and_50_enex5;
  wire PECore_PushAxiRsp_if_and_51_enex5;
  wire PECore_PushAxiRsp_if_and_52_enex5;
  wire PECore_PushAxiRsp_if_and_53_enex5;
  wire PECore_PushAxiRsp_if_and_54_enex5;
  wire PECore_PushAxiRsp_if_and_55_enex5;
  wire PECore_PushAxiRsp_if_and_56_enex5;
  wire PECore_PushAxiRsp_if_and_57_enex5;
  wire PECore_PushAxiRsp_if_and_58_enex5;
  wire PECore_PushAxiRsp_if_and_59_enex5;
  wire PECore_PushOutput_if_and_16_enex5;
  wire PECore_PushOutput_if_and_17_enex5;
  wire PECore_PushOutput_if_and_18_enex5;
  wire PECore_PushOutput_if_and_19_enex5;
  wire PECore_PushOutput_if_and_20_enex5;
  wire PECore_PushOutput_if_and_21_enex5;
  wire PECore_PushOutput_if_and_22_enex5;
  wire PECore_PushOutput_if_and_25_enex5;
  wire PECore_PushOutput_if_and_26_enex5;
  wire PECore_PushOutput_if_and_28_enex5;
  wire PECore_PushOutput_if_and_29_enex5;
  wire PECore_PushOutput_if_and_30_enex5;
  wire PECore_PushOutput_if_and_31_enex5;
  wire act_port_reg_data_and_enex5;
  wire act_port_reg_data_and_28_enex5;
  wire act_port_reg_data_and_29_enex5;
  wire act_port_reg_data_and_30_enex5;
  wire Datapath_for_and_enex5;
  wire PECore_RunMac_if_and_854_tmp;
  wire PECore_RunMac_if_and_865_tmp;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_15_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse;
  wire PECore_RunMac_if_and_860_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_1_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_2_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_3_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_4_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_5_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_6_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_7_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_8_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_9_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_10_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_11_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_12_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_13_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_14_itm;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_1;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_2;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_3;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_4;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_5;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_6;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_7;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_8;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_9;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_10;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_11;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_12;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_13;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_14;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_14;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_13;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_12;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_11;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_10;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_9;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_8;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_7;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_6;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_5;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_4;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_3;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_2;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_1;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_2;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_14;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_13;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_12;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_11;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_10;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_9;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_8;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_7;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_6;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_5;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_4;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_3;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_2;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_1;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_0;
  wire [11:0] operator_16_false_1_mux_10_cse;
  wire operator_16_false_1_mux_14_cse;
  wire z_out_10_13;
  wire z_out_11_13;
  wire z_out_12_13;
  wire z_out_13_13;
  wire z_out_21_32;
  wire z_out_22_32;
  wire z_out_23_32;
  wire z_out_24_32;
  wire [15:0] operator_16_false_1_mux_16_cse;
  wire while_mux_440_cse;
  wire adpfloat_tmp_to_fixed_20U_14U_mux1h_28_tmp;
  wire or_3880_tmp;
  wire while_while_mux_15_m1c;
  wire while_mux1h_62_m1c;
  wire while_while_mux_13_m1c;
  wire while_mux1h_57_m1c;
  wire while_while_mux_11_m1c;
  wire while_mux1h_52_m1c;
  wire while_while_mux_9_m1c;
  wire while_mux1h_47_m1c;
  wire PEManager_16U_GetInputAddr_1_PEManager_16U_GetInputAddr_1_mux_5_tmp;
  wire adpfloat_tmp_to_fixed_20U_14U_mux1h_29_tmp;
  wire adpfloat_tmp_to_fixed_20U_14U_mux1h_30_tmp;
  wire adpfloat_tmp_to_fixed_20U_14U_mux1h_32_tmp;
  wire while_while_nor_cse;
  wire while_and_268_cse;

  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_10;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_10;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_11;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_12;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_12;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_13;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_28;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_28;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_28;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_28;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_14;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_14;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_29;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_29;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_29;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_29;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_30;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_30;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_30;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_30;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_15;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_31;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_31;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_31;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_31;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_32;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_32;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_32;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_32;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_16;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_16;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_33;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_33;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_33;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_33;
  wire PECore_PushAxiRsp_if_else_mux_14_nl;
  wire PECore_DecodeAxi_mux_139_nl;
  wire PECore_DecodeAxi_if_mux_74_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_19_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_11_nl;
  wire[6:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_18_nl;
  wire PECore_PushAxiRsp_if_else_mux_15_nl;
  wire PECore_DecodeAxi_mux_141_nl;
  wire PECore_DecodeAxi_if_mux_126_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_17_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_8_nl;
  wire[1:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl;
  wire[4:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_15_nl;
  wire PECore_PushAxiRsp_if_else_mux_16_nl;
  wire PECore_DecodeAxi_mux_143_nl;
  wire PECore_DecodeAxi_if_mux_127_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_13_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_5_nl;
  wire[1:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_12_nl;
  wire[4:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_10_nl;
  wire PECore_PushAxiRsp_if_else_mux_17_nl;
  wire PECore_DecodeAxi_mux_145_nl;
  wire PECore_DecodeAxi_if_mux_128_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_12_nl;
  wire[1:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_9_nl;
  wire[4:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl;
  wire input_mem_banks_read_read_data_and_nl;
  wire mux_594_nl;
  wire or_1536_nl;
  wire mux_593_nl;
  wire mux_592_nl;
  wire mux_591_nl;
  wire nor_244_nl;
  wire or_1531_nl;
  wire or_1530_nl;
  wire mux_596_nl;
  wire mux_595_nl;
  wire nor_242_nl;
  wire nor_243_nl;
  wire mux_600_nl;
  wire mux_599_nl;
  wire mux_598_nl;
  wire nor_241_nl;
  wire mux_597_nl;
  wire PECore_UpdateFSM_switch_lp_mux_6_nl;
  wire PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_7_nl;
  wire and_3383_nl;
  wire PECore_UpdateFSM_switch_lp_mux1h_42_nl;
  wire PECore_UpdateFSM_switch_lp_not_47_nl;
  wire PECore_UpdateFSM_switch_lp_not_48_nl;
  wire PECore_UpdateFSM_switch_lp_not_49_nl;
  wire while_and_221_nl;
  wire while_and_225_nl;
  wire while_and_226_nl;
  wire while_and_227_nl;
  wire[19:0] mux1h_12_nl;
  wire while_or_11_nl;
  wire while_and_288_nl;
  wire while_and_289_nl;
  wire while_mux1h_46_nl;
  wire while_and_222_nl;
  wire while_and_223_nl;
  wire while_and_224_nl;
  wire while_and_290_nl;
  wire while_mux1h_48_nl;
  wire PECore_RunBias_if_for_and_55_nl;
  wire PECore_RunBias_if_for_and_56_nl;
  wire PECore_RunBias_if_for_and_57_nl;
  wire while_mux1h_49_nl;
  wire while_and_228_nl;
  wire while_and_229_nl;
  wire while_and_230_nl;
  wire PECore_UpdateFSM_switch_lp_not_65_nl;
  wire while_and_231_nl;
  wire while_and_235_nl;
  wire while_and_236_nl;
  wire while_and_237_nl;
  wire[19:0] mux1h_13_nl;
  wire while_or_10_nl;
  wire while_and_283_nl;
  wire while_and_284_nl;
  wire while_mux1h_51_nl;
  wire while_and_232_nl;
  wire while_and_233_nl;
  wire while_and_234_nl;
  wire while_and_285_nl;
  wire while_mux1h_53_nl;
  wire PECore_RunBias_if_for_and_58_nl;
  wire PECore_RunBias_if_for_and_59_nl;
  wire PECore_RunBias_if_for_and_60_nl;
  wire while_mux1h_54_nl;
  wire while_and_238_nl;
  wire while_and_239_nl;
  wire while_and_240_nl;
  wire PECore_UpdateFSM_switch_lp_not_66_nl;
  wire while_and_241_nl;
  wire while_and_245_nl;
  wire while_and_246_nl;
  wire while_and_247_nl;
  wire[19:0] mux1h_14_nl;
  wire while_or_9_nl;
  wire while_and_278_nl;
  wire while_and_279_nl;
  wire while_mux1h_56_nl;
  wire while_and_242_nl;
  wire while_and_243_nl;
  wire while_and_244_nl;
  wire while_and_280_nl;
  wire while_mux1h_58_nl;
  wire PECore_RunBias_if_for_and_61_nl;
  wire PECore_RunBias_if_for_and_62_nl;
  wire PECore_RunBias_if_for_and_63_nl;
  wire while_mux1h_59_nl;
  wire while_and_248_nl;
  wire PECore_UpdateFSM_switch_lp_not_67_nl;
  wire while_and_249_nl;
  wire while_and_253_nl;
  wire while_and_254_nl;
  wire while_and_255_nl;
  wire[19:0] mux1h_15_nl;
  wire while_or_nl;
  wire while_and_273_nl;
  wire while_and_274_nl;
  wire while_mux1h_61_nl;
  wire while_and_250_nl;
  wire while_and_251_nl;
  wire while_and_252_nl;
  wire while_and_275_nl;
  wire while_mux1h_63_nl;
  wire PECore_RunBias_if_for_and_64_nl;
  wire PECore_RunBias_if_for_and_65_nl;
  wire PECore_RunBias_if_for_and_66_nl;
  wire while_mux1h_64_nl;
  wire while_and_256_nl;
  wire PECore_UpdateFSM_switch_lp_not_38_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_if_1_crossbar_spec_PE_Weight_WordType_16U_16U_for_if_1_crossbar_spec_PE_Weight_WordType_16U_16U_for_if_1_nor_5_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_252_nl;
  wire[3:0] pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_and_1_nl;
  wire pe_config_UpdateManagerCounter_if_not_7_nl;
  wire and_3501_nl;
  wire[31:0] while_mux1h_67_nl;
  wire while_and_269_nl;
  wire while_and_270_nl;
  wire PECore_UpdateFSM_switch_lp_not_55_nl;
  wire[31:0] while_mux_nl;
  wire PECore_UpdateFSM_switch_lp_not_56_nl;
  wire[31:0] while_mux1h_65_nl;
  wire PECore_UpdateFSM_switch_lp_not_57_nl;
  wire[31:0] while_mux_449_nl;
  wire PECore_UpdateFSM_switch_lp_not_58_nl;
  wire[19:0] while_while_mux1h_12_nl;
  wire while_and_202_nl;
  wire while_and_203_nl;
  wire while_and_204_nl;
  wire PECore_RunBias_if_for_and_25_nl;
  wire while_and_82_nl;
  wire PECore_UpdateFSM_switch_lp_not_36_nl;
  wire[19:0] while_while_mux1h_13_nl;
  wire while_and_199_nl;
  wire while_and_200_nl;
  wire while_and_201_nl;
  wire PECore_RunBias_if_for_and_27_nl;
  wire while_and_84_nl;
  wire PECore_UpdateFSM_switch_lp_not_64_nl;
  wire[19:0] while_while_mux1h_14_nl;
  wire while_and_196_nl;
  wire while_and_197_nl;
  wire while_and_198_nl;
  wire PECore_RunBias_if_for_and_29_nl;
  wire while_and_86_nl;
  wire PECore_UpdateFSM_switch_lp_not_63_nl;
  wire[19:0] while_while_mux1h_15_nl;
  wire while_and_193_nl;
  wire while_and_194_nl;
  wire while_and_195_nl;
  wire PECore_RunBias_if_for_and_31_nl;
  wire while_and_88_nl;
  wire PECore_UpdateFSM_switch_lp_not_62_nl;
  wire PECore_UpdateFSM_switch_lp_mux_7_nl;
  wire pe_config_UpdateManagerCounter_mux_1_nl;
  wire pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl;
  wire and_3991_nl;
  wire[7:0] pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl;
  wire pe_config_UpdateInputCounter_if_not_2_nl;
  wire PECore_UpdateFSM_switch_lp_and_nl;
  wire[7:0] pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl;
  wire pe_config_UpdateManagerCounter_if_not_9_nl;
  wire and_4037_nl;
  wire PECore_UpdateFSM_switch_lp_not_50_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_94_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_92_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_90_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_88_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_86_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_84_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_82_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_80_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_81_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_83_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_85_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_87_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_89_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_91_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_93_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_95_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_78_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_76_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_74_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_72_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_70_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_68_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_66_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_64_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_65_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_67_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_69_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_71_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_73_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_75_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_77_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_79_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_62_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_60_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_58_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_56_nl;
  wire[2:0] PEManager_16U_ClusterLookup_for_mux_54_nl;
  wire[4:0] PECore_RunBias_if_for_10_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_10_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_10_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_10_operator_33_true_acc_nl;
  wire[4:0] PEManager_16U_ClusterLookup_for_mux_139_nl;
  wire[2:0] PEManager_16U_ClusterLookup_for_mux_52_nl;
  wire[4:0] PECore_RunBias_if_for_11_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_11_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_11_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_11_operator_33_true_acc_nl;
  wire[4:0] PEManager_16U_ClusterLookup_for_mux_140_nl;
  wire[2:0] PEManager_16U_ClusterLookup_for_mux_50_nl;
  wire[4:0] PEManager_16U_ClusterLookup_for_mux_141_nl;
  wire[4:0] PECore_RunBias_if_for_5_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_5_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_5_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_5_operator_33_true_acc_nl;
  wire PECore_RunMac_if_and_829_nl;
  wire[2:0] PEManager_16U_ClusterLookup_for_mux_48_nl;
  wire[4:0] PECore_RunBias_if_for_6_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_6_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_6_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_6_operator_33_true_acc_nl;
  wire[4:0] PEManager_16U_ClusterLookup_for_mux_142_nl;
  wire[2:0] PEManager_16U_ClusterLookup_for_mux_49_nl;
  wire[4:0] PECore_RunBias_if_for_7_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_7_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_7_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_7_operator_33_true_acc_nl;
  wire[4:0] PEManager_16U_ClusterLookup_for_mux_143_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_51_nl;
  wire[4:0] PECore_RunBias_if_for_8_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_8_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_8_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_8_operator_33_true_acc_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_53_nl;
  wire[4:0] PECore_RunBias_if_for_9_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_9_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_9_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_9_operator_33_true_acc_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_55_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_57_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_59_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_61_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_63_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_46_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_44_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_42_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_40_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_38_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_36_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_34_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_32_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_33_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_35_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_37_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_39_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_41_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_43_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_45_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_47_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_2_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux1h_6_nl;
  wire PECore_RunBias_if_for_and_49_nl;
  wire PECore_RunBias_if_for_and_40_nl;
  wire PECore_RunBias_if_for_and_36_nl;
  wire PECore_DecodeAxi_mux_133_nl;
  wire PECore_DecodeAxi_if_mux_67_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_or_1_nl;
  wire adpfloat_tmp_is_zero_if_adpfloat_tmp_is_zero_if_nor_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_29_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_7_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_62_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_28_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_8_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_60_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_27_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_9_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_58_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_26_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_10_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_56_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_25_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_19_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_49_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_18_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_51_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_20_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_48_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_21_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_4_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_22_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_52_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_20_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_23_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_50_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_and_3_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_9_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_11_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_54_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux1h_13_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux1h_11_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux1h_16_nl;
  wire PECore_DecodeAxi_mux_138_nl;
  wire PECore_DecodeAxi_if_mux_125_nl;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_or_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_258_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_257_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_256_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_255_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_254_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_251_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_250_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_249_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_248_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_247_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_246_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_245_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_244_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_253_nl;
  wire PECore_RunMac_nor_nl;
  wire PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl;
  wire PECore_UpdateFSM_case_1_if_mux_nl;
  wire pe_manager_zero_active_mux_nl;
  wire PECore_DecodeAxi_mux_127_nl;
  wire PECore_DecodeAxi_if_mux_57_nl;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_34_nl;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_32_nl;
  wire pe_manager_zero_active_mux_1_nl;
  wire PECore_DecodeAxi_mux_125_nl;
  wire PECore_DecodeAxi_if_mux_55_nl;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_35_nl;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_33_nl;
  wire[2:0] PEManager_16U_ClusterLookup_for_mux_15_nl;
  wire[4:0] PEManager_16U_ClusterLookup_for_mux_145_nl;
  wire[4:0] PECore_RunBias_if_for_3_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_3_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_3_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_3_operator_33_true_acc_nl;
  wire[2:0] PEManager_16U_ClusterLookup_for_mux_6_nl;
  wire[4:0] PEManager_16U_ClusterLookup_for_mux_144_nl;
  wire[4:0] PECore_RunBias_if_for_4_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_4_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_4_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_4_operator_33_true_acc_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_3_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_74_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_72_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_70_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_68_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_66_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_64_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_65_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_30_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_94_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_31_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_92_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_32_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_90_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_33_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_88_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_34_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_86_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_35_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_84_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_36_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_82_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_37_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_80_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_38_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_81_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_39_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_83_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_40_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_85_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_41_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_87_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_42_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_89_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_43_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_91_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_44_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_93_nl;
  wire[7:0] data_in_tmp_operator_for_mux_34_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_95_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_46_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_44_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_42_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_40_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_38_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_36_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_34_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_32_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_33_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_35_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_37_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_39_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_41_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_43_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_45_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_47_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_30_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_28_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_26_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_24_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_22_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_20_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_18_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_16_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_17_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_19_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_21_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_23_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_25_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_27_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_29_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_31_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_30_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_28_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_26_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_24_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_22_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_20_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_18_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_16_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_17_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_19_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_21_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_23_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_25_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_27_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_29_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_31_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_1_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_2_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_3_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_4_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_5_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_6_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_7_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_8_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_9_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_10_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_11_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_12_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_13_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_14_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_15_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_14_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_13_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_12_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_11_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_10_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_9_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_8_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_7_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_1_nl;
  wire mux_22_nl;
  wire nand_198_nl;
  wire nor_475_nl;
  wire pe_config_is_cluster_not_39_nl;
  wire[11:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_40_nl;
  wire[11:0] PECore_RunFSM_switch_lp_mux_28_nl;
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_43_nl;
  wire PECore_RunFSM_switch_lp_mux_29_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3212_nl;
  wire weight_mem_run_1_if_for_if_and_702_nl;
  wire PECore_DecodeAxi_mux_134_nl;
  wire PECore_DecodeAxi_if_mux_122_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_mux_5_nl;
  wire PECore_DecodeAxi_mux_135_nl;
  wire PECore_DecodeAxi_if_mux_123_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_or_nl;
  wire PECore_RunFSM_case_0_if_mux_1_nl;
  wire or_1624_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_465_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_466_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_468_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_469_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_470_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_471_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_472_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_473_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_474_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_475_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_476_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_477_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_478_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_479_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_1_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_2995_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_2994_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_2992_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_2988_nl;
  wire[15:0] operator_16_false_1_acc_12_nl;
  wire[16:0] nl_operator_16_false_1_acc_12_nl;
  wire[14:0] operator_16_false_1_acc_nl;
  wire[15:0] nl_operator_16_false_1_acc_nl;
  wire[15:0] operator_16_false_1_acc_11_nl;
  wire[16:0] nl_operator_16_false_1_acc_11_nl;
  wire[13:0] operator_16_false_1_acc_8_nl;
  wire[14:0] nl_operator_16_false_1_acc_8_nl;
  wire[13:0] operator_16_false_1_mux_20_nl;
  wire[15:0] operator_16_false_1_acc_10_nl;
  wire[16:0] nl_operator_16_false_1_acc_10_nl;
  wire[14:0] operator_16_false_1_acc_7_nl;
  wire[15:0] nl_operator_16_false_1_acc_7_nl;
  wire[15:0] operator_16_false_1_acc_9_nl;
  wire[16:0] nl_operator_16_false_1_acc_9_nl;
  wire[12:0] operator_16_false_1_acc_3_nl;
  wire[13:0] nl_operator_16_false_1_acc_3_nl;
  wire[15:0] PECore_RunFSM_case_2_else_for_10_operator_16_false_1_acc_nl;
  wire[16:0] nl_PECore_RunFSM_case_2_else_for_10_operator_16_false_1_acc_nl;
  wire[14:0] operator_16_false_1_acc_4_nl;
  wire[15:0] nl_operator_16_false_1_acc_4_nl;
  wire[15:0] PECore_RunFSM_case_2_else_for_12_operator_16_false_1_acc_nl;
  wire[16:0] nl_PECore_RunFSM_case_2_else_for_12_operator_16_false_1_acc_nl;
  wire[13:0] operator_16_false_1_acc_5_nl;
  wire[14:0] nl_operator_16_false_1_acc_5_nl;
  wire[15:0] PECore_RunFSM_case_2_else_for_14_operator_16_false_1_acc_nl;
  wire[16:0] nl_PECore_RunFSM_case_2_else_for_14_operator_16_false_1_acc_nl;
  wire[14:0] operator_16_false_1_acc_6_nl;
  wire[15:0] nl_operator_16_false_1_acc_6_nl;
  wire[15:0] PECore_RunFSM_case_2_else_for_16_operator_16_false_1_acc_nl;
  wire[16:0] nl_PECore_RunFSM_case_2_else_for_16_operator_16_false_1_acc_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_1_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_435_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_436_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_438_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_439_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_440_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_441_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_442_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_443_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_444_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_445_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_446_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_447_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_448_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_449_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_2_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3009_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3008_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3006_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3002_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_2_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_405_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_406_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_408_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_409_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_410_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_411_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_412_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_413_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_414_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_415_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_416_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_417_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_418_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_419_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_3_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3023_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3022_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3020_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3016_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_3_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_375_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_376_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_378_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_379_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_380_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_381_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_382_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_383_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_384_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_385_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_386_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_387_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_388_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_389_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_4_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3037_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3036_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3034_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3030_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_4_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_345_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_346_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_348_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_349_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_350_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_351_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_352_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_353_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_354_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_355_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_356_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_357_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_358_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_359_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_5_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3051_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3050_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3048_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3044_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_5_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_315_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_316_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_318_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_319_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_320_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_321_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_322_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_323_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_324_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_325_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_326_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_327_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_328_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_329_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_6_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3065_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3064_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3062_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3058_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_6_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_285_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_286_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_288_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_289_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_290_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_291_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_292_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_293_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_294_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_295_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_296_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_297_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_298_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_299_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_7_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3079_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3078_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3076_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3072_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_7_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_255_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_256_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_258_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_259_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_260_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_261_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_262_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_263_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_264_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_265_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_266_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_267_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_268_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_269_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_8_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3093_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3092_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3090_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3086_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_8_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_225_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_226_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_228_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_229_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_230_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_231_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_232_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_233_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_234_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_235_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_236_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_237_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_238_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_239_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_9_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3107_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3106_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3104_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3100_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_9_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_195_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_196_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_198_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_199_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_200_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_201_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_202_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_203_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_204_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_205_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_206_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_207_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_208_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_209_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_10_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3121_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3120_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3118_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3114_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_10_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_165_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_166_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_168_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_169_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_170_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_171_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_172_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_173_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_174_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_175_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_176_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_177_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_178_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_179_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_11_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3135_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3134_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3132_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3128_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_11_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_135_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_136_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_138_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_139_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_140_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_141_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_142_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_143_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_144_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_145_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_146_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_147_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_148_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_149_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_12_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3149_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3148_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3146_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3142_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_12_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_105_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_106_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_108_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_109_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_110_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_111_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_112_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_113_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_114_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_115_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_116_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_117_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_118_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_119_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_13_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3163_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3162_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3160_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3156_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_13_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_75_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_76_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_78_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_79_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_80_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_81_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_82_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_83_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_84_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_85_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_86_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_87_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_88_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_89_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_14_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3177_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3176_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3174_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3170_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_14_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_45_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_46_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_48_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_49_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_50_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_51_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_52_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_53_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_54_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_55_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_56_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_57_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_58_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_59_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_15_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3191_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3190_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3188_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3184_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_15_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_15_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_16_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_18_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_19_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_20_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_21_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_22_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_23_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_24_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_25_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_26_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_27_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_28_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_29_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_16_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3216_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3218_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3219_nl;
  wire weight_mem_run_1_if_for_if_and_697_nl;
  wire weight_mem_run_1_if_for_if_and_693_nl;
  wire weight_mem_run_1_if_for_if_and_689_nl;
  wire weight_mem_run_1_if_for_if_and_690_nl;
  wire weight_mem_run_1_if_for_if_and_694_nl;
  wire weight_mem_run_1_if_for_if_and_698_nl;
  wire weight_mem_run_1_if_for_if_and_703_nl;
  wire weight_mem_run_1_if_for_if_and_701_nl;
  wire weight_mem_run_1_if_for_if_and_699_nl;
  wire weight_mem_run_1_if_for_if_and_695_nl;
  wire weight_mem_run_1_if_for_if_and_688_nl;
  wire weight_mem_run_1_if_for_if_and_692_nl;
  wire weight_mem_run_1_if_for_if_and_696_nl;
  wire weight_mem_run_1_if_for_if_and_700_nl;
  wire PECore_DecodeAxi_mux_149_nl;
  wire PECore_DecodeAxi_if_mux_135_nl;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_56_nl;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_54_nl;
  wire[7:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_mux1h_nl;
  wire PECore_UpdateFSM_switch_lp_or_nl;
  wire PECore_UpdateFSM_switch_lp_and_2_nl;
  wire PECore_UpdateFSM_switch_lp_and_3_nl;
  wire[7:0] PECore_DecodeAxi_if_mux_68_nl;
  wire[3:0] PECore_DecodeAxi_if_mux_69_nl;
  wire weight_mem_run_1_if_for_if_and_691_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_260_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_262_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_264_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_266_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_268_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_270_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_272_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_274_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_276_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_278_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_280_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_282_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_284_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_286_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_256_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_258_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_332_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_347_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_362_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_377_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_392_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_407_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_422_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_437_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_452_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_467_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_482_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_497_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_512_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_527_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_302_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_317_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_331_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_346_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_361_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_376_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_391_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_406_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_421_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_436_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_451_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_466_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_481_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_496_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_511_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_526_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_301_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_316_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_330_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_345_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_360_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_375_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_390_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_405_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_420_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_435_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_450_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_465_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_480_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_495_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_510_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_525_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_300_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_315_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_329_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_344_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_359_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_374_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_389_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_404_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_419_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_434_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_449_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_464_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_479_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_494_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_509_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_524_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_299_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_314_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_328_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_343_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_358_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_373_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_388_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_403_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_418_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_433_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_448_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_463_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_478_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_493_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_508_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_523_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_298_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_313_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_327_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_342_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_357_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_372_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_387_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_402_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_417_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_432_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_447_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_462_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_477_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_492_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_507_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_522_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_297_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_312_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_326_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_341_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_356_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_371_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_386_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_401_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_416_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_431_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_446_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_461_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_476_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_491_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_506_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_521_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_296_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_311_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_325_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_340_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_355_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_370_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_385_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_400_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_415_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_430_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_445_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_460_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_475_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_490_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_505_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_520_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_295_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_310_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_324_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_339_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_354_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_369_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_384_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_399_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_414_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_429_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_444_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_459_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_474_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_489_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_504_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_519_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_294_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_309_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_323_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_338_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_353_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_368_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_383_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_398_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_413_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_428_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_443_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_458_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_473_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_488_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_503_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_518_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_293_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_308_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_322_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_337_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_352_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_367_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_382_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_397_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_412_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_427_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_442_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_457_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_472_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_487_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_502_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_517_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_292_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_307_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_321_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_336_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_351_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_366_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_381_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_396_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_411_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_426_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_441_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_456_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_471_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_486_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_501_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_516_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_291_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_306_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_320_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_335_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_350_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_365_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_380_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_395_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_410_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_425_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_440_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_455_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_470_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_485_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_500_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_515_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_290_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_305_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_319_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_334_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_349_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_364_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_379_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_394_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_409_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_424_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_439_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_454_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_469_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_484_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_499_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_514_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_289_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_304_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_318_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_333_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_348_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_363_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_378_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_393_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_408_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_423_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_438_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_453_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_468_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_483_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_498_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_513_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_288_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_303_nl;
  wire[7:0] while_mux_111_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_36_nl;
  wire[7:0] while_mux_110_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_35_nl;
  wire[7:0] while_mux_109_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_34_nl;
  wire[7:0] while_mux_108_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_33_nl;
  wire[7:0] while_mux_107_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_32_nl;
  wire[7:0] while_mux_106_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_31_nl;
  wire[7:0] while_mux_105_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_30_nl;
  wire[7:0] while_mux_104_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_29_nl;
  wire[7:0] while_mux_103_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_28_nl;
  wire[7:0] while_mux_102_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_27_nl;
  wire[7:0] while_mux_101_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_26_nl;
  wire[7:0] while_mux_100_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_25_nl;
  wire[7:0] while_mux_99_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_24_nl;
  wire[7:0] while_mux_98_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_23_nl;
  wire[7:0] while_mux_97_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_22_nl;
  wire[7:0] while_mux_96_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_21_nl;
  wire[7:0] mux1h_7_nl;
  wire[7:0] PEManager_16U_GetInputAddr_1_acc_nl;
  wire[8:0] nl_PEManager_16U_GetInputAddr_1_acc_nl;
  wire[7:0] PEManager_16U_GetBiasAddr_acc_nl;
  wire[8:0] nl_PEManager_16U_GetBiasAddr_acc_nl;
  wire PECore_DecodeAxi_if_and_nl;
  wire PECore_DecodeAxi_if_and_1_nl;
  wire not_3760_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_35_nl;
  wire[7:0] PEManager_16U_GetInputAddr_acc_nl;
  wire[8:0] nl_PEManager_16U_GetInputAddr_acc_nl;
  wire or_1589_nl;
  wire mux_601_nl;
  wire and_1488_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_53_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_133_nl;
  wire[3:0] PEManager_16U_ClusterLookup_for_mux_5_nl;
  wire[3:0] PEManager_16U_ClusterLookup_for_mux_138_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_55_nl;
  wire[3:0] PECore_DecodeAxiRead_case_4_switch_lp_and_1_nl;
  wire[3:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_5_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_132_nl;
  wire and_5134_nl;
  wire and_5136_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_and_1_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_and_2_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_57_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_131_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_59_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_130_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_61_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_129_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_63_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_128_nl;
  wire[3:0] PEManager_16U_ClusterLookup_for_mux_78_nl;
  wire[3:0] PEManager_16U_ClusterLookup_for_mux_137_nl;
  wire[3:0] PEManager_16U_ClusterLookup_for_mux_76_nl;
  wire[3:0] PEManager_16U_ClusterLookup_for_mux_136_nl;
  wire[5:0] PEManager_16U_ClusterLookup_for_mux_67_nl;
  wire[1:0] PECore_DecodeAxiRead_case_4_switch_lp_and_9_nl;
  wire[1:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_10_nl;
  wire[1:0] PEManager_16U_ClusterLookup_for_mux_135_nl;
  wire[2:0] PEManager_16U_ClusterLookup_for_mux_69_nl;
  wire[4:0] PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_12_nl;
  wire[4:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_2_nl;
  wire[4:0] PECore_RunBias_if_for_12_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_12_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_12_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_12_operator_33_true_acc_nl;
  wire[4:0] PEManager_16U_ClusterLookup_for_mux_134_nl;
  wire[5:0] PEManager_16U_ClusterLookup_for_mux_71_nl;
  wire[1:0] PECore_DecodeAxiRead_case_4_switch_lp_and_7_nl;
  wire[1:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_4_nl;
  wire[1:0] PEManager_16U_ClusterLookup_for_mux_133_nl;
  wire[2:0] PEManager_16U_ClusterLookup_for_mux_2_nl;
  wire[4:0] PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_10_nl;
  wire[4:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_nl;
  wire[4:0] PEManager_16U_ClusterLookup_for_mux_132_nl;
  wire[5:0] PEManager_16U_ClusterLookup_for_mux_73_nl;
  wire[1:0] PECore_DecodeAxiRead_case_4_switch_lp_and_6_nl;
  wire[1:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_1_nl;
  wire[1:0] PEManager_16U_ClusterLookup_for_mux_131_nl;
  wire[2:0] PEManager_16U_ClusterLookup_for_mux_75_nl;
  wire[4:0] PEManager_16U_ClusterLookup_for_mux_130_nl;
  wire[4:0] PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_11_nl;
  wire[4:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_1_nl;
  wire[4:0] PECore_RunBias_if_for_2_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_2_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_2_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_2_operator_33_true_acc_nl;
  wire PECore_RunMac_if_and_803_nl;
  wire[3:0] PEManager_16U_ClusterLookup_for_mux_77_nl;
  wire[3:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl;
  wire[3:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_24_nl;
  wire[3:0] PEManager_16U_ClusterLookup_for_mux_129_nl;
  wire rva_out_reg_data_and_1_nl;
  wire PECore_RunMac_if_and_801_nl;
  wire PEManager_16U_ClusterLookup_for_mux_79_nl;
  wire[6:0] PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_13_nl;
  wire[6:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl;
  wire[6:0] PEManager_16U_ClusterLookup_for_mux_128_nl;
  wire[3:0] operator_4_false_mux_2_nl;
  wire[2:0] PECore_RunBias_if_for_1_operator_33_true_acc_1_nl;
  wire[3:0] nl_PECore_RunBias_if_for_1_operator_33_true_acc_1_nl;
  wire[7:0] operator_8_false_mux_2_nl;
  wire and_5952_nl;
  wire[13:0] operator_32_true_acc_nl;
  wire[14:0] nl_operator_32_true_acc_nl;
  wire[12:0] operator_32_true_mux1h_40_nl;
  wire[13:0] operator_32_true_acc_1_nl;
  wire[14:0] nl_operator_32_true_acc_1_nl;
  wire[12:0] operator_32_true_mux1h_41_nl;
  wire[13:0] operator_32_true_acc_2_nl;
  wire[14:0] nl_operator_32_true_acc_2_nl;
  wire[12:0] operator_32_true_mux1h_42_nl;
  wire[13:0] operator_32_true_acc_3_nl;
  wire[14:0] nl_operator_32_true_acc_3_nl;
  wire[12:0] operator_32_true_mux1h_43_nl;
  wire[19:0] adpfloat_tmp_to_fixed_20U_14U_if_1_adpfloat_tmp_to_fixed_20U_14U_if_1_mux_2_nl;
  wire[19:0] adpfloat_tmp_to_fixed_20U_14U_if_1_mux1h_8_nl;
  wire[19:0] adpfloat_tmp_to_fixed_20U_14U_if_1_adpfloat_tmp_to_fixed_20U_14U_if_1_mux_3_nl;
  wire[19:0] adpfloat_tmp_to_fixed_20U_14U_if_1_mux1h_9_nl;
  wire[32:0] operator_32_true_acc_nl_1;
  wire[33:0] nl_operator_32_true_acc_nl_1;
  wire[31:0] operator_32_true_mux1h_8_nl;
  wire[32:0] operator_32_true_acc_1_nl_1;
  wire[33:0] nl_operator_32_true_acc_1_nl_1;
  wire[31:0] operator_32_true_mux1h_9_nl;
  wire[32:0] operator_32_true_acc_2_nl_1;
  wire[33:0] nl_operator_32_true_acc_2_nl_1;
  wire[31:0] operator_32_true_mux1h_10_nl;
  wire[32:0] operator_32_true_acc_3_nl_1;
  wire[33:0] nl_operator_32_true_acc_3_nl_1;
  wire[31:0] operator_32_true_mux1h_11_nl;
  wire[31:0] PECore_RunMac_if_for_mux1h_4_nl;
  wire[31:0] PECore_RunMac_if_for_mux1h_5_nl;
  wire[31:0] PECore_RunMac_if_for_mux1h_6_nl;
  wire[31:0] PECore_RunMac_if_for_mux1h_7_nl;
  wire[19:0] and_5953_nl;
  wire[19:0] mux1h_16_nl;
  wire[19:0] PECore_RunBias_if_for_if_or_8_nl;
  wire[19:0] PECore_RunBias_if_for_if_mux1h_4_nl;
  wire PECore_RunBias_if_for_if_and_8_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_8_nl;
  wire PECore_RunBias_if_for_if_or_9_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_12_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_13_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_14_nl;
  wire nor_599_nl;
  wire[19:0] and_5961_nl;
  wire[19:0] mux_645_nl;
  wire[19:0] PECore_RunBias_if_for_if_or_10_nl;
  wire[19:0] PECore_RunBias_if_for_if_mux1h_5_nl;
  wire PECore_RunBias_if_for_if_and_9_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_9_nl;
  wire PECore_RunBias_if_for_if_and_10_nl;
  wire or_3882_nl;
  wire nor_603_nl;
  wire[19:0] and_5968_nl;
  wire[19:0] mux_646_nl;
  wire[19:0] PECore_RunBias_if_for_if_or_11_nl;
  wire[19:0] PECore_RunBias_if_for_if_mux1h_6_nl;
  wire PECore_RunBias_if_for_if_and_11_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_10_nl;
  wire PECore_RunBias_if_for_if_and_12_nl;
  wire or_3883_nl;
  wire nor_607_nl;
  wire[19:0] and_5975_nl;
  wire[19:0] mux_647_nl;
  wire[19:0] PECore_RunBias_if_for_if_or_12_nl;
  wire[19:0] PECore_RunBias_if_for_if_mux1h_7_nl;
  wire PECore_RunBias_if_for_if_and_13_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_11_nl;
  wire PECore_RunBias_if_for_if_and_14_nl;
  wire or_3884_nl;
  wire nor_611_nl;
  wire[2:0] operator_3_false_mux_2_nl;
  wire[2:0] PECore_RunBias_if_right_shift_mux_2_nl;
  wire[2:0] operator_3_false_mux_3_nl;
  wire[2:0] PECore_RunBias_if_right_shift_mux_3_nl;
  wire and_5982_nl;
  wire PEManager_16U_GetInputAddr_1_PEManager_16U_GetInputAddr_1_nor_nl;
  wire PEManager_16U_GetInputAddr_1_and_1_nl;
  wire PEManager_16U_GetInputAddr_1_and_2_nl;
  wire PEManager_16U_GetInputAddr_1_and_3_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_adpfloat_tmp_to_fixed_20U_14U_nor_8_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_16_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_17_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_18_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_adpfloat_tmp_to_fixed_20U_14U_nor_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_20_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_21_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_22_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_23_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_24_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_25_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_26_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_27_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[7:0] PECore_RunMac_if_mux1h_63_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_127_nl;
  wire[7:0] PECore_RunMac_if_mux1h_62_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_126_nl;
  wire[7:0] PECore_RunMac_if_mux1h_61_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_124_nl;
  wire[7:0] PECore_RunMac_if_mux1h_60_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_122_nl;
  wire[7:0] PECore_RunMac_if_mux1h_59_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_120_nl;
  wire[7:0] PECore_RunMac_if_mux1h_58_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_118_nl;
  wire[7:0] PECore_RunMac_if_mux1h_57_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_116_nl;
  wire[7:0] PECore_RunMac_if_mux1h_56_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_114_nl;
  wire[7:0] PECore_RunMac_if_mux1h_55_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_112_nl;
  wire[7:0] PECore_RunMac_if_mux1h_54_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_113_nl;
  wire[7:0] PECore_RunMac_if_mux1h_53_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_115_nl;
  wire[7:0] PECore_RunMac_if_mux1h_52_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_117_nl;
  wire[7:0] PECore_RunMac_if_mux1h_51_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_119_nl;
  wire[7:0] PECore_RunMac_if_mux1h_50_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_121_nl;
  wire[7:0] PECore_RunMac_if_mux1h_49_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_123_nl;
  wire[7:0] PECore_RunMac_if_mux1h_48_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_125_nl;
  wire [127:0] nl_Datapath_for_1_ProductSum_cmp_in_1_data_rsc_dat;
  assign PEManager_16U_ClusterLookup_1_for_mux_127_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_15_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_63_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_175_itm,
      PEManager_16U_ClusterLookup_1_for_mux_127_nl, weight_port_read_out_data_15_15_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      PECore_RunMac_if_mux_15_itm, reg_Datapath_for_conc_4_ftd, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_112_cse , PECore_RunMac_if_and_113_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_126_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_15_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_62_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_174_itm,
      PEManager_16U_ClusterLookup_1_for_mux_126_nl, weight_port_read_out_data_15_14_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      ({reg_PECore_RunMac_if_mux_14_ftd , reg_PECore_RunMac_if_mux_14_ftd_1}), reg_Datapath_for_conc_4_ftd_1,
      {or_tmp_1334 , PECore_RunMac_if_and_434_cse , PECore_RunMac_if_and_112_cse
      , PECore_RunMac_if_and_113_cse , (fsm_output[3]) , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_124_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_14_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_61_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_173_itm,
      PEManager_16U_ClusterLookup_1_for_mux_124_nl, weight_port_read_out_data_15_13_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      PECore_RunMac_if_mux_13_itm, reg_Datapath_for_conc_4_ftd_2, {or_tmp_1334 ,
      PECore_RunMac_if_and_434_cse , PECore_RunMac_if_and_112_cse , PECore_RunMac_if_and_113_cse
      , (fsm_output[3]) , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_122_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_14_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_60_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_172_itm,
      PEManager_16U_ClusterLookup_1_for_mux_122_nl, weight_port_read_out_data_15_12_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_13_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      rva_out_reg_data_79_72_sva_dfm_4, reg_Datapath_for_conc_4_ftd_3, {or_tmp_1334
      , PECore_RunMac_if_and_434_cse , PECore_RunMac_if_and_112_cse , PECore_RunMac_if_and_113_cse
      , (fsm_output[3]) , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_120_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_13_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_59_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_171_itm,
      PEManager_16U_ClusterLookup_1_for_mux_120_nl, weight_port_read_out_data_15_11_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_12_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      ({reg_PECore_RunMac_if_mux_11_ftd , reg_PECore_RunMac_if_mux_11_ftd_1}), reg_Datapath_for_conc_4_ftd_4,
      {or_tmp_1334 , PECore_RunMac_if_and_434_cse , PECore_RunMac_if_and_112_cse
      , PECore_RunMac_if_and_113_cse , (fsm_output[3]) , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_118_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_13_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_58_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_170_itm,
      PEManager_16U_ClusterLookup_1_for_mux_118_nl, weight_port_read_out_data_15_10_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_11_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      ({reg_PECore_RunMac_if_mux_10_ftd , reg_PECore_RunMac_if_mux_10_ftd_1}), reg_Datapath_for_conc_4_ftd_5,
      {or_tmp_1334 , PECore_RunMac_if_and_434_cse , PECore_RunMac_if_and_112_cse
      , PECore_RunMac_if_and_113_cse , (fsm_output[3]) , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_116_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_12_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_57_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_169_itm,
      PEManager_16U_ClusterLookup_1_for_mux_116_nl, weight_port_read_out_data_15_9_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_10_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      PECore_RunMac_if_mux_9_itm, reg_Datapath_for_conc_4_ftd_6, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_112_cse , PECore_RunMac_if_and_113_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_114_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_12_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_56_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_168_itm,
      PEManager_16U_ClusterLookup_1_for_mux_114_nl, weight_port_read_out_data_15_8_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_9_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      PECore_RunMac_if_mux_8_itm, reg_Datapath_for_conc_4_ftd_7, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_112_cse , PECore_RunMac_if_and_113_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_112_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_11_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_55_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_167_itm,
      PEManager_16U_ClusterLookup_1_for_mux_112_nl, weight_port_read_out_data_15_7_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_8_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      PECore_RunMac_if_mux_7_itm, reg_Datapath_for_conc_4_ftd_8, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_112_cse , PECore_RunMac_if_and_113_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_113_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_11_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_54_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_166_itm,
      PEManager_16U_ClusterLookup_1_for_mux_113_nl, weight_port_read_out_data_15_6_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_7_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      PECore_RunMac_if_mux_6_itm, reg_Datapath_for_conc_4_ftd_9, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_112_cse , PECore_RunMac_if_and_113_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_115_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_10_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_53_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_165_itm,
      PEManager_16U_ClusterLookup_1_for_mux_115_nl, weight_port_read_out_data_15_5_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_6_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      PECore_RunMac_if_mux_5_itm, reg_Datapath_for_conc_4_ftd_10, {or_tmp_1334 ,
      PECore_RunMac_if_and_434_cse , PECore_RunMac_if_and_112_cse , PECore_RunMac_if_and_113_cse
      , (fsm_output[3]) , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_117_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_10_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_52_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_164_itm,
      PEManager_16U_ClusterLookup_1_for_mux_117_nl, weight_port_read_out_data_15_4_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_5_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      PECore_RunMac_if_mux_4_itm, reg_Datapath_for_conc_4_ftd_11, {or_tmp_1334 ,
      PECore_RunMac_if_and_434_cse , PECore_RunMac_if_and_112_cse , PECore_RunMac_if_and_113_cse
      , (fsm_output[3]) , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_119_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_9_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_51_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_163_itm,
      PEManager_16U_ClusterLookup_1_for_mux_119_nl, weight_port_read_out_data_15_3_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_4_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      PECore_RunMac_if_mux_3_itm, reg_Datapath_for_conc_4_ftd_12, {or_tmp_1334 ,
      PECore_RunMac_if_and_434_cse , PECore_RunMac_if_and_112_cse , PECore_RunMac_if_and_113_cse
      , (fsm_output[3]) , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_121_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_9_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_50_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_162_itm,
      PEManager_16U_ClusterLookup_1_for_mux_121_nl, weight_port_read_out_data_15_2_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_3_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      PECore_RunMac_if_mux_2_itm, reg_Datapath_for_conc_4_ftd_13, {or_tmp_1334 ,
      PECore_RunMac_if_and_434_cse , PECore_RunMac_if_and_112_cse , PECore_RunMac_if_and_113_cse
      , (fsm_output[3]) , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_123_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_8_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_49_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_161_itm,
      PEManager_16U_ClusterLookup_1_for_mux_123_nl, weight_port_read_out_data_15_1_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_2_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      ({reg_PECore_RunMac_if_mux_1_ftd , reg_PECore_RunMac_if_mux_1_ftd_1}), reg_Datapath_for_conc_4_ftd_14,
      {or_tmp_1334 , PECore_RunMac_if_and_434_cse , PECore_RunMac_if_and_112_cse
      , PECore_RunMac_if_and_113_cse , (fsm_output[3]) , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_125_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_8_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_48_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_160_itm,
      PEManager_16U_ClusterLookup_1_for_mux_125_nl, weight_port_read_out_data_15_0_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_1_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      PECore_RunMac_if_mux_itm, reg_Datapath_for_conc_4_ftd_15, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_112_cse , PECore_RunMac_if_and_113_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign nl_Datapath_for_1_ProductSum_cmp_in_1_data_rsc_dat = {PECore_RunMac_if_mux1h_63_nl
      , PECore_RunMac_if_mux1h_62_nl , PECore_RunMac_if_mux1h_61_nl , PECore_RunMac_if_mux1h_60_nl
      , PECore_RunMac_if_mux1h_59_nl , PECore_RunMac_if_mux1h_58_nl , PECore_RunMac_if_mux1h_57_nl
      , PECore_RunMac_if_mux1h_56_nl , PECore_RunMac_if_mux1h_55_nl , PECore_RunMac_if_mux1h_54_nl
      , PECore_RunMac_if_mux1h_53_nl , PECore_RunMac_if_mux1h_52_nl , PECore_RunMac_if_mux1h_51_nl
      , PECore_RunMac_if_mux1h_50_nl , PECore_RunMac_if_mux1h_49_nl , PECore_RunMac_if_mux1h_48_nl};
  wire[7:0] PECore_RunMac_if_mux1h_47_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_111_nl;
  wire[7:0] PECore_RunMac_if_mux1h_46_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_109_nl;
  wire[7:0] PECore_RunMac_if_mux1h_45_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_107_nl;
  wire[7:0] PECore_RunMac_if_mux1h_44_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_105_nl;
  wire[7:0] PECore_RunMac_if_mux1h_43_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_103_nl;
  wire[7:0] PECore_RunMac_if_mux1h_42_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_101_nl;
  wire[7:0] PECore_RunMac_if_mux1h_41_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_99_nl;
  wire[7:0] PECore_RunMac_if_mux1h_40_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_97_nl;
  wire[7:0] PECore_RunMac_if_mux1h_39_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_96_nl;
  wire[7:0] PECore_RunMac_if_mux1h_38_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_98_nl;
  wire[7:0] PECore_RunMac_if_mux1h_37_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_100_nl;
  wire[7:0] PECore_RunMac_if_mux1h_36_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_102_nl;
  wire[7:0] PECore_RunMac_if_mux1h_35_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_104_nl;
  wire[7:0] PECore_RunMac_if_mux1h_34_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_106_nl;
  wire[7:0] PECore_RunMac_if_mux1h_33_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_108_nl;
  wire[7:0] PECore_RunMac_if_mux1h_32_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_110_nl;
  wire [127:0] nl_Datapath_for_1_ProductSum_cmp_1_in_1_data_rsc_dat;
  assign PEManager_16U_ClusterLookup_1_for_mux_111_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_15_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_47_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_95_itm,
      PEManager_16U_ClusterLookup_1_for_mux_111_nl, weight_port_read_out_data_13_15_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      PECore_RunMac_if_mux_191_itm, PECore_RunMac_if_mux_79_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_144_cse , PECore_RunMac_if_and_145_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_109_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_15_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_46_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_94_itm,
      PEManager_16U_ClusterLookup_1_for_mux_109_nl, weight_port_read_out_data_13_14_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      PECore_RunMac_if_mux_190_itm, PECore_RunMac_if_mux_78_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_144_cse , PECore_RunMac_if_and_145_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_107_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_14_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_45_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_93_itm,
      PEManager_16U_ClusterLookup_1_for_mux_107_nl, weight_port_read_out_data_13_13_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_15,
      PECore_RunMac_if_mux_189_itm, PECore_RunMac_if_mux_77_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_144_cse , PECore_RunMac_if_and_145_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_105_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_14_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_44_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_92_itm,
      PEManager_16U_ClusterLookup_1_for_mux_105_nl, weight_port_read_out_data_13_12_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_17,
      PECore_RunMac_if_mux_188_itm, PECore_RunMac_if_mux_76_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_144_cse , PECore_RunMac_if_and_145_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_103_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_13_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_43_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_91_itm,
      PEManager_16U_ClusterLookup_1_for_mux_103_nl, weight_port_read_out_data_13_11_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_19,
      PECore_RunMac_if_mux_187_itm, PECore_RunMac_if_mux_75_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_144_cse , PECore_RunMac_if_and_145_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_101_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_13_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_42_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_90_itm,
      PEManager_16U_ClusterLookup_1_for_mux_101_nl, weight_port_read_out_data_13_10_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_21,
      PECore_RunMac_if_mux_186_itm, PECore_RunMac_if_mux_74_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_144_cse , PECore_RunMac_if_and_145_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_99_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_12_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_41_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_89_itm,
      PEManager_16U_ClusterLookup_1_for_mux_99_nl, weight_port_read_out_data_13_9_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_23,
      PECore_RunMac_if_mux_185_itm, PECore_RunMac_if_mux_73_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_144_cse , PECore_RunMac_if_and_145_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_97_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_12_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_40_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_88_itm,
      PEManager_16U_ClusterLookup_1_for_mux_97_nl, weight_port_read_out_data_13_8_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_25,
      PECore_RunMac_if_mux_184_itm, PECore_RunMac_if_mux_72_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_144_cse , PECore_RunMac_if_and_145_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_96_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_11_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_39_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_87_itm,
      PEManager_16U_ClusterLookup_1_for_mux_96_nl, weight_port_read_out_data_13_7_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_27,
      PECore_RunMac_if_mux_183_itm, PECore_RunMac_if_mux_71_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_144_cse , PECore_RunMac_if_and_145_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_98_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_11_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_38_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_86_itm,
      PEManager_16U_ClusterLookup_1_for_mux_98_nl, weight_port_read_out_data_13_6_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_29,
      PECore_RunMac_if_mux_182_itm, PECore_RunMac_if_mux_70_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_144_cse , PECore_RunMac_if_and_145_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_100_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_10_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_37_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_85_itm,
      PEManager_16U_ClusterLookup_1_for_mux_100_nl, weight_port_read_out_data_13_5_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_31,
      PECore_RunMac_if_mux_181_itm, PECore_RunMac_if_mux_69_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_144_cse , PECore_RunMac_if_and_145_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_102_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_10_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_36_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_84_itm,
      PEManager_16U_ClusterLookup_1_for_mux_102_nl, weight_port_read_out_data_13_4_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_33,
      PECore_RunMac_if_mux_180_itm, PECore_RunMac_if_mux_68_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_144_cse , PECore_RunMac_if_and_145_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_104_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_9_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_35_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_83_itm,
      PEManager_16U_ClusterLookup_1_for_mux_104_nl, weight_port_read_out_data_13_3_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_35,
      PECore_RunMac_if_mux_179_itm, PECore_RunMac_if_mux_67_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_144_cse , PECore_RunMac_if_and_145_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_106_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_9_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_34_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_82_itm,
      PEManager_16U_ClusterLookup_1_for_mux_106_nl, weight_port_read_out_data_13_2_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_37,
      PECore_RunMac_if_mux_178_itm, PECore_RunMac_if_mux_66_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_144_cse , PECore_RunMac_if_and_145_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_108_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_8_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_33_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_81_itm,
      PEManager_16U_ClusterLookup_1_for_mux_108_nl, weight_port_read_out_data_13_1_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_39,
      PECore_RunMac_if_mux_177_itm, PECore_RunMac_if_mux_65_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_144_cse , PECore_RunMac_if_and_145_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_110_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_8_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_32_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_80_itm,
      PEManager_16U_ClusterLookup_1_for_mux_110_nl, weight_port_read_out_data_13_0_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_41,
      PECore_RunMac_if_mux_176_itm, PECore_RunMac_if_mux_64_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_144_cse , PECore_RunMac_if_and_145_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign nl_Datapath_for_1_ProductSum_cmp_1_in_1_data_rsc_dat = {PECore_RunMac_if_mux1h_47_nl
      , PECore_RunMac_if_mux1h_46_nl , PECore_RunMac_if_mux1h_45_nl , PECore_RunMac_if_mux1h_44_nl
      , PECore_RunMac_if_mux1h_43_nl , PECore_RunMac_if_mux1h_42_nl , PECore_RunMac_if_mux1h_41_nl
      , PECore_RunMac_if_mux1h_40_nl , PECore_RunMac_if_mux1h_39_nl , PECore_RunMac_if_mux1h_38_nl
      , PECore_RunMac_if_mux1h_37_nl , PECore_RunMac_if_mux1h_36_nl , PECore_RunMac_if_mux1h_35_nl
      , PECore_RunMac_if_mux1h_34_nl , PECore_RunMac_if_mux1h_33_nl , PECore_RunMac_if_mux1h_32_nl};
  wire[7:0] PECore_RunMac_if_mux1h_31_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_127_nl;
  wire[7:0] PECore_RunMac_if_mux1h_30_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_125_nl;
  wire[7:0] PECore_RunMac_if_mux1h_29_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_123_nl;
  wire[7:0] PECore_RunMac_if_mux1h_28_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_121_nl;
  wire[7:0] PECore_RunMac_if_mux1h_27_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_119_nl;
  wire[7:0] PECore_RunMac_if_mux1h_26_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_117_nl;
  wire[7:0] PECore_RunMac_if_mux1h_25_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_115_nl;
  wire[7:0] PECore_RunMac_if_mux1h_24_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_113_nl;
  wire[7:0] PECore_RunMac_if_mux1h_23_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_112_nl;
  wire[7:0] PECore_RunMac_if_mux1h_22_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_114_nl;
  wire[7:0] PECore_RunMac_if_mux1h_21_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_116_nl;
  wire[7:0] PECore_RunMac_if_mux1h_20_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_118_nl;
  wire[7:0] PECore_RunMac_if_mux1h_19_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_120_nl;
  wire[7:0] PECore_RunMac_if_mux1h_18_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_122_nl;
  wire[7:0] PECore_RunMac_if_mux1h_17_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_124_nl;
  wire[7:0] PECore_RunMac_if_mux1h_16_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_126_nl;
  wire [127:0] nl_Datapath_for_1_ProductSum_cmp_2_in_1_data_rsc_dat;
  assign PEManager_16U_ClusterLookup_for_mux_127_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_7_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_31_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_111_itm,
      PEManager_16U_ClusterLookup_for_mux_127_nl, weight_port_read_out_data_14_15_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      ({reg_PECore_RunMac_if_mux_143_ftd , reg_PECore_RunMac_if_mux_143_ftd_1}),
      PECore_RunMac_if_mux_63_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse ,
      PECore_RunMac_if_and_176_cse , PECore_RunMac_if_and_177_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_125_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_7_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_30_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_110_itm,
      PEManager_16U_ClusterLookup_for_mux_125_nl, weight_port_read_out_data_14_14_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      ({reg_PECore_RunMac_if_mux_142_ftd , reg_PECore_RunMac_if_mux_142_ftd_1}),
      PECore_RunMac_if_mux_62_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse ,
      PECore_RunMac_if_and_176_cse , PECore_RunMac_if_and_177_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_123_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_6_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_29_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_109_itm,
      PEManager_16U_ClusterLookup_for_mux_123_nl, weight_port_read_out_data_14_13_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      ({reg_PECore_RunMac_if_mux_141_ftd , reg_PECore_RunMac_if_mux_141_ftd_1}),
      PECore_RunMac_if_mux_61_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse ,
      PECore_RunMac_if_and_176_cse , PECore_RunMac_if_and_177_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_121_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_6_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_28_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_108_itm,
      PEManager_16U_ClusterLookup_for_mux_121_nl, weight_port_read_out_data_14_12_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_13_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      ({reg_PECore_RunMac_if_mux_140_ftd , reg_PECore_RunMac_if_mux_140_ftd_1}),
      PECore_RunMac_if_mux_60_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse ,
      PECore_RunMac_if_and_176_cse , PECore_RunMac_if_and_177_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_119_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_5_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_27_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_107_itm,
      PEManager_16U_ClusterLookup_for_mux_119_nl, weight_port_read_out_data_14_11_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_12_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      ({reg_PECore_RunMac_if_mux_139_ftd , reg_PECore_RunMac_if_mux_139_ftd_1}),
      PECore_RunMac_if_mux_59_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse ,
      PECore_RunMac_if_and_176_cse , PECore_RunMac_if_and_177_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_117_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_5_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_26_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_106_itm,
      PEManager_16U_ClusterLookup_for_mux_117_nl, weight_port_read_out_data_14_10_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_11_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      ({reg_PECore_RunMac_if_mux_138_ftd , reg_PECore_RunMac_if_mux_138_ftd_1}),
      PECore_RunMac_if_mux_58_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse ,
      PECore_RunMac_if_and_176_cse , PECore_RunMac_if_and_177_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_115_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_4_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_25_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_105_itm,
      PEManager_16U_ClusterLookup_for_mux_115_nl, weight_port_read_out_data_14_9_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_10_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      ({reg_PECore_RunMac_if_mux_137_ftd , reg_PECore_RunMac_if_mux_137_ftd_1}),
      PECore_RunMac_if_mux_57_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse ,
      PECore_RunMac_if_and_176_cse , PECore_RunMac_if_and_177_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_113_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_4_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_24_nl = MUX1HOT_v_8_6_2(({reg_PECore_RunMac_if_mux_104_ftd
      , reg_PECore_RunMac_if_mux_104_ftd_1}), PEManager_16U_ClusterLookup_for_mux_113_nl,
      weight_port_read_out_data_14_8_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_9_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      PECore_RunMac_if_mux_136_itm, PECore_RunMac_if_mux_56_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_176_cse , PECore_RunMac_if_and_177_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_112_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_3_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_23_nl = MUX1HOT_v_8_6_2(({reg_PECore_RunMac_if_mux_103_ftd
      , reg_PECore_RunMac_if_mux_103_ftd_1}), PEManager_16U_ClusterLookup_for_mux_112_nl,
      weight_port_read_out_data_14_7_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_8_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      PECore_RunMac_if_mux_135_itm, PECore_RunMac_if_mux_55_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_176_cse , PECore_RunMac_if_and_177_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_114_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_3_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_22_nl = MUX1HOT_v_8_6_2(({reg_PECore_RunMac_if_mux_102_ftd
      , reg_PECore_RunMac_if_mux_102_ftd_1}), PEManager_16U_ClusterLookup_for_mux_114_nl,
      weight_port_read_out_data_14_6_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_7_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      PECore_RunMac_if_mux_134_itm, PECore_RunMac_if_mux_54_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_176_cse , PECore_RunMac_if_and_177_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_116_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_2_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_21_nl = MUX1HOT_v_8_6_2(({reg_PECore_RunMac_if_mux_101_ftd
      , reg_PECore_RunMac_if_mux_101_ftd_1}), PEManager_16U_ClusterLookup_for_mux_116_nl,
      weight_port_read_out_data_14_5_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_6_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      PECore_RunMac_if_mux_133_itm, PECore_RunMac_if_mux_53_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_176_cse , PECore_RunMac_if_and_177_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_118_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_2_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_20_nl = MUX1HOT_v_8_6_2(({reg_PECore_RunMac_if_mux_100_ftd
      , reg_PECore_RunMac_if_mux_100_ftd_1}), PEManager_16U_ClusterLookup_for_mux_118_nl,
      weight_port_read_out_data_14_4_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_5_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      PECore_RunMac_if_mux_132_itm, PECore_RunMac_if_mux_52_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_176_cse , PECore_RunMac_if_and_177_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_120_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_1_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_19_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_99_itm,
      PEManager_16U_ClusterLookup_for_mux_120_nl, weight_port_read_out_data_14_3_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_4_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      PECore_RunMac_if_mux_131_itm, PECore_RunMac_if_mux_51_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_176_cse , PECore_RunMac_if_and_177_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_122_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_1_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_18_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_98_itm,
      PEManager_16U_ClusterLookup_for_mux_122_nl, weight_port_read_out_data_14_2_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_3_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      PECore_RunMac_if_mux_130_itm, PECore_RunMac_if_mux_50_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse
      , PECore_RunMac_if_and_176_cse , PECore_RunMac_if_and_177_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_124_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_0_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_17_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_97_itm,
      PEManager_16U_ClusterLookup_for_mux_124_nl, weight_port_read_out_data_14_1_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_2_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      ({reg_PECore_RunMac_if_mux_129_ftd , reg_PECore_RunMac_if_mux_129_ftd_1}),
      PECore_RunMac_if_mux_49_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse ,
      PECore_RunMac_if_and_176_cse , PECore_RunMac_if_and_177_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_126_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_7_0_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_16_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_96_itm,
      PEManager_16U_ClusterLookup_for_mux_126_nl, weight_port_read_out_data_14_0_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_1_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      ({reg_PECore_RunMac_if_mux_128_ftd , reg_PECore_RunMac_if_mux_128_ftd_1}),
      PECore_RunMac_if_mux_48_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse ,
      PECore_RunMac_if_and_176_cse , PECore_RunMac_if_and_177_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign nl_Datapath_for_1_ProductSum_cmp_2_in_1_data_rsc_dat = {PECore_RunMac_if_mux1h_31_nl
      , PECore_RunMac_if_mux1h_30_nl , PECore_RunMac_if_mux1h_29_nl , PECore_RunMac_if_mux1h_28_nl
      , PECore_RunMac_if_mux1h_27_nl , PECore_RunMac_if_mux1h_26_nl , PECore_RunMac_if_mux1h_25_nl
      , PECore_RunMac_if_mux1h_24_nl , PECore_RunMac_if_mux1h_23_nl , PECore_RunMac_if_mux1h_22_nl
      , PECore_RunMac_if_mux1h_21_nl , PECore_RunMac_if_mux1h_20_nl , PECore_RunMac_if_mux1h_19_nl
      , PECore_RunMac_if_mux1h_18_nl , PECore_RunMac_if_mux1h_17_nl , PECore_RunMac_if_mux1h_16_nl};
  wire[7:0] PECore_RunMac_if_mux1h_15_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_111_nl;
  wire[7:0] PECore_RunMac_if_mux1h_14_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_109_nl;
  wire[7:0] PECore_RunMac_if_mux1h_13_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_107_nl;
  wire[7:0] PECore_RunMac_if_mux1h_12_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_105_nl;
  wire[7:0] PECore_RunMac_if_mux1h_11_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_103_nl;
  wire[7:0] PECore_RunMac_if_mux1h_10_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_101_nl;
  wire[7:0] PECore_RunMac_if_mux1h_9_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_99_nl;
  wire[7:0] PECore_RunMac_if_mux1h_8_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_97_nl;
  wire[7:0] PECore_RunMac_if_mux1h_7_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_96_nl;
  wire[7:0] PECore_RunMac_if_mux1h_6_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_98_nl;
  wire[7:0] PECore_RunMac_if_mux1h_5_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_100_nl;
  wire[7:0] PECore_RunMac_if_mux1h_4_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_102_nl;
  wire[7:0] PECore_RunMac_if_mux1h_3_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_104_nl;
  wire[7:0] PECore_RunMac_if_mux1h_2_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_106_nl;
  wire[7:0] PECore_RunMac_if_mux1h_1_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_108_nl;
  wire[7:0] PECore_RunMac_if_mux1h_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_110_nl;
  wire [127:0] nl_Datapath_for_1_ProductSum_cmp_3_in_1_data_rsc_dat;
  assign PEManager_16U_ClusterLookup_for_mux_111_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_7_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_15_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_159_itm,
      PEManager_16U_ClusterLookup_for_mux_111_nl, weight_port_read_out_data_12_15_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1,
      ({reg_PECore_RunMac_if_mux_127_ftd , reg_PECore_RunMac_if_mux_127_ftd_1}),
      PECore_RunMac_if_mux_47_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse ,
      PECore_RunMac_if_and_208_cse , PECore_RunMac_if_and_209_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_109_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_7_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_14_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_158_itm,
      PEManager_16U_ClusterLookup_for_mux_109_nl, weight_port_read_out_data_12_14_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1,
      ({reg_PECore_RunMac_if_mux_126_ftd , reg_PECore_RunMac_if_mux_126_ftd_1}),
      PECore_RunMac_if_mux_46_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse ,
      PECore_RunMac_if_and_208_cse , PECore_RunMac_if_and_209_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_107_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_6_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_13_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_157_itm,
      PEManager_16U_ClusterLookup_for_mux_107_nl, weight_port_read_out_data_12_13_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1,
      ({reg_PECore_RunMac_if_mux_125_ftd , reg_PECore_RunMac_if_mux_125_ftd_1}),
      PECore_RunMac_if_mux_45_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse ,
      PECore_RunMac_if_and_208_cse , PECore_RunMac_if_and_209_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_105_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_6_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_12_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_156_itm,
      PEManager_16U_ClusterLookup_for_mux_105_nl, weight_port_read_out_data_12_12_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1,
      ({reg_PECore_RunMac_if_mux_124_ftd , reg_PECore_RunMac_if_mux_124_ftd_1}),
      PECore_RunMac_if_mux_44_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse ,
      PECore_RunMac_if_and_208_cse , PECore_RunMac_if_and_209_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_103_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_5_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_11_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_155_itm,
      PEManager_16U_ClusterLookup_for_mux_103_nl, weight_port_read_out_data_12_11_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1,
      ({reg_PECore_RunMac_if_mux_123_ftd , reg_PECore_RunMac_if_mux_123_ftd_1}),
      PECore_RunMac_if_mux_43_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse ,
      PECore_RunMac_if_and_208_cse , PECore_RunMac_if_and_209_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_101_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_5_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_10_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_154_itm,
      PEManager_16U_ClusterLookup_for_mux_101_nl, weight_port_read_out_data_12_10_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1,
      ({reg_PECore_RunMac_if_mux_122_ftd , reg_PECore_RunMac_if_mux_122_ftd_1}),
      PECore_RunMac_if_mux_42_itm, {or_tmp_1334 , PECore_RunMac_if_and_434_cse ,
      PECore_RunMac_if_and_208_cse , PECore_RunMac_if_and_209_cse , (fsm_output[3])
      , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_99_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_4_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_9_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_153_itm,
      PEManager_16U_ClusterLookup_for_mux_99_nl, weight_port_read_out_data_12_9_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1,
      rva_out_reg_data_95_88_sva_dfm_4, PECore_RunMac_if_mux_41_itm, {or_tmp_1334
      , PECore_RunMac_if_and_434_cse , PECore_RunMac_if_and_208_cse , PECore_RunMac_if_and_209_cse
      , (fsm_output[3]) , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_97_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_4_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_8_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_152_itm,
      PEManager_16U_ClusterLookup_for_mux_97_nl, weight_port_read_out_data_12_8_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1,
      rva_out_reg_data_87_80_sva_dfm_4, PECore_RunMac_if_mux_40_itm, {or_tmp_1334
      , PECore_RunMac_if_and_434_cse , PECore_RunMac_if_and_208_cse , PECore_RunMac_if_and_209_cse
      , (fsm_output[3]) , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_96_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_3_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_7_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_151_itm,
      PEManager_16U_ClusterLookup_for_mux_96_nl, weight_port_read_out_data_12_7_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1,
      rva_out_reg_data_71_64_sva_dfm_4, PECore_RunMac_if_mux_39_itm, {or_tmp_1334
      , PECore_RunMac_if_and_434_cse , PECore_RunMac_if_and_208_cse , PECore_RunMac_if_and_209_cse
      , (fsm_output[3]) , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_98_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_3_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_6_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_150_itm,
      PEManager_16U_ClusterLookup_for_mux_98_nl, weight_port_read_out_data_12_6_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1,
      rva_out_reg_data_63_56_sva_dfm_4, PECore_RunMac_if_mux_38_itm, {or_tmp_1334
      , PECore_RunMac_if_and_434_cse , PECore_RunMac_if_and_208_cse , PECore_RunMac_if_and_209_cse
      , (fsm_output[3]) , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_100_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_2_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_5_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_149_itm,
      PEManager_16U_ClusterLookup_for_mux_100_nl, weight_port_read_out_data_12_5_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1,
      rva_out_reg_data_55_48_sva_dfm_4, PECore_RunMac_if_mux_37_itm, {or_tmp_1334
      , PECore_RunMac_if_and_434_cse , PECore_RunMac_if_and_208_cse , PECore_RunMac_if_and_209_cse
      , (fsm_output[3]) , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_102_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_2_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_4_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_148_itm,
      PEManager_16U_ClusterLookup_for_mux_102_nl, weight_port_read_out_data_12_4_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1,
      rva_out_reg_data_47_40_sva_dfm_4, PECore_RunMac_if_mux_36_itm, {or_tmp_1334
      , PECore_RunMac_if_and_434_cse , PECore_RunMac_if_and_208_cse , PECore_RunMac_if_and_209_cse
      , (fsm_output[3]) , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_104_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_1_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_3_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_147_itm,
      PEManager_16U_ClusterLookup_for_mux_104_nl, weight_port_read_out_data_12_3_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1,
      rva_out_reg_data_127_120_sva_dfm_4, PECore_RunMac_if_mux_35_itm, {or_tmp_1334
      , PECore_RunMac_if_and_434_cse , PECore_RunMac_if_and_208_cse , PECore_RunMac_if_and_209_cse
      , (fsm_output[3]) , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_106_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_1_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_2_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_146_itm,
      PEManager_16U_ClusterLookup_for_mux_106_nl, weight_port_read_out_data_12_2_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1,
      rva_out_reg_data_119_112_sva_dfm_4, PECore_RunMac_if_mux_34_itm, {or_tmp_1334
      , PECore_RunMac_if_and_434_cse , PECore_RunMac_if_and_208_cse , PECore_RunMac_if_and_209_cse
      , (fsm_output[3]) , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_108_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_0_sva_dfm_mx1[7:4])});
  assign PECore_RunMac_if_mux1h_1_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_145_itm,
      PEManager_16U_ClusterLookup_for_mux_108_nl, weight_port_read_out_data_12_1_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1,
      rva_out_reg_data_111_104_sva_dfm_4, PECore_RunMac_if_mux_33_itm, {or_tmp_1334
      , PECore_RunMac_if_and_434_cse , PECore_RunMac_if_and_208_cse , PECore_RunMac_if_and_209_cse
      , (fsm_output[3]) , (fsm_output[4])});
  assign PEManager_16U_ClusterLookup_for_mux_110_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_6_0_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_if_mux1h_nl = MUX1HOT_v_8_6_2(PECore_RunMac_if_mux_144_itm,
      PEManager_16U_ClusterLookup_for_mux_110_nl, weight_port_read_out_data_12_0_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1,
      rva_out_reg_data_103_96_sva_dfm_4, PECore_RunMac_if_mux_32_itm, {or_tmp_1334
      , PECore_RunMac_if_and_434_cse , PECore_RunMac_if_and_208_cse , PECore_RunMac_if_and_209_cse
      , (fsm_output[3]) , (fsm_output[4])});
  assign nl_Datapath_for_1_ProductSum_cmp_3_in_1_data_rsc_dat = {PECore_RunMac_if_mux1h_15_nl
      , PECore_RunMac_if_mux1h_14_nl , PECore_RunMac_if_mux1h_13_nl , PECore_RunMac_if_mux1h_12_nl
      , PECore_RunMac_if_mux1h_11_nl , PECore_RunMac_if_mux1h_10_nl , PECore_RunMac_if_mux1h_9_nl
      , PECore_RunMac_if_mux1h_8_nl , PECore_RunMac_if_mux1h_7_nl , PECore_RunMac_if_mux1h_6_nl
      , PECore_RunMac_if_mux1h_5_nl , PECore_RunMac_if_mux1h_4_nl , PECore_RunMac_if_mux1h_3_nl
      , PECore_RunMac_if_mux1h_2_nl , PECore_RunMac_if_mux1h_1_nl , PECore_RunMac_if_mux1h_nl};
  wire [7:0] nl_PEManager_16U_GetWeightAddr_if_acc_4_cmp_a;
  assign nl_PEManager_16U_GetWeightAddr_if_acc_4_cmp_a = pe_config_output_counter_sva;
  wire [7:0] nl_PEManager_16U_GetWeightAddr_if_acc_4_cmp_b;
  assign nl_PEManager_16U_GetWeightAddr_if_acc_4_cmp_b = MUX_v_8_2_2(pe_manager_num_input_0_sva,
      pe_manager_num_input_1_sva, pe_config_manager_counter_sva[0]);
  wire [7:0] nl_PEManager_16U_GetWeightAddr_if_acc_4_cmp_c;
  assign nl_PEManager_16U_GetWeightAddr_if_acc_4_cmp_c = pe_config_input_counter_sva;
  wire  nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a;
  assign nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a = PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0
      & (rva_in_PopNB_mio_mrgout_dat_sva_1[168]) & PECore_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_mx1
      & (~ is_start_sva);
  wire [3:0] nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s;
  assign nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s = weight_write_addrs_lpi_1_dfm_6[3:0];
  wire [3:0] nl_weight_mem_read_arbxbar_xbar_for_15_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_for_15_lshift_rg_s = {(weight_read_addrs_14_15_1_lpi_1_dfm_3[2:0])
      , weight_read_addrs_10_0_lpi_1_dfm_2};
  wire [3:0] nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s = {weight_read_addrs_0_3_lpi_1_dfm_5_mx0
      , weight_read_addrs_0_2_0_lpi_1_dfm_4_2_mx0 , weight_read_addrs_0_2_0_lpi_1_dfm_4_1_mx0
      , weight_read_addrs_0_2_0_lpi_1_dfm_4_0_mx0};
  wire [3:0] nl_weight_mem_read_arbxbar_xbar_for_11_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_for_11_lshift_rg_s = {(weight_read_addrs_10_15_1_lpi_1_dfm_3[2:0])
      , weight_read_addrs_10_0_lpi_1_dfm_2};
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_50_nl;
  wire [3:0] nl_weight_mem_read_arbxbar_xbar_for_13_lshift_rg_s;
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_50_nl
      = (weight_read_addrs_8_2_0_lpi_1_dfm_1[1]) & PECore_RunFSM_switch_lp_equal_tmp_5;
  assign nl_weight_mem_read_arbxbar_xbar_for_13_lshift_rg_s = {(weight_read_addrs_12_15_2_lpi_1_dfm_3[1:0])
      , PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_50_nl
      , weight_read_addrs_10_0_lpi_1_dfm_2};
  wire [3:0] nl_weight_mem_read_arbxbar_xbar_for_16_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_for_16_lshift_rg_s = weight_read_addrs_15_lpi_1_dfm_3[3:0];
  wire [3:0] nl_weight_mem_read_arbxbar_xbar_for_12_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_for_12_lshift_rg_s = weight_read_addrs_11_lpi_1_dfm_3[3:0];
  wire [3:0] nl_weight_mem_read_arbxbar_xbar_for_14_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_for_14_lshift_rg_s = weight_read_addrs_13_lpi_1_dfm_3[3:0];
  wire [3:0] nl_weight_mem_read_arbxbar_xbar_for_7_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_for_7_lshift_rg_s = {(weight_read_addrs_6_15_1_lpi_1_dfm_2[2:0])
      , (weight_read_addrs_4_1_0_lpi_1_dfm_1[0])};
  wire[2:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_46_nl;
  wire [3:0] nl_weight_mem_read_arbxbar_xbar_for_9_lshift_rg_s;
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_46_nl
      = MUX_v_3_2_2(3'b000, weight_read_addrs_8_2_0_lpi_1_dfm_1, PECore_RunFSM_switch_lp_equal_tmp_5);
  assign nl_weight_mem_read_arbxbar_xbar_for_9_lshift_rg_s = {(weight_read_addrs_8_15_3_lpi_1_dfm_3[0])
      , PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_46_nl};
  wire [3:0] nl_weight_mem_read_arbxbar_xbar_for_3_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_for_3_lshift_rg_s = {(weight_read_addrs_2_15_1_lpi_1_dfm_2[2:0])
      , (weight_read_addrs_4_1_0_lpi_1_dfm_1[0])};
  wire [3:0] nl_weight_mem_read_arbxbar_xbar_for_5_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_for_5_lshift_rg_s = {(weight_read_addrs_4_15_2_lpi_1_dfm_2[1:0])
      , weight_read_addrs_4_1_0_lpi_1_dfm_1};
  wire [3:0] nl_weight_mem_read_arbxbar_xbar_for_8_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_for_8_lshift_rg_s = weight_read_addrs_7_lpi_1_dfm_2[3:0];
  wire [3:0] nl_weight_mem_read_arbxbar_xbar_for_4_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_for_4_lshift_rg_s = weight_read_addrs_3_lpi_1_dfm_2[3:0];
  wire [3:0] nl_weight_mem_read_arbxbar_xbar_for_6_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_for_6_lshift_rg_s = weight_read_addrs_5_lpi_1_dfm_2[3:0];
  wire [3:0] nl_weight_mem_read_arbxbar_xbar_for_10_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_for_10_lshift_rg_s = weight_read_addrs_9_lpi_1_dfm_3[3:0];
  wire [3:0] nl_weight_mem_read_arbxbar_xbar_for_2_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_for_2_lshift_rg_s = weight_read_addrs_1_lpi_1_dfm_2[3:0];
  wire [31:0] nl_PECore_RunBias_if_for_14_PECore_RunBias_if_for_rshift_1_rg_a;
  assign nl_PECore_RunBias_if_for_14_PECore_RunBias_if_for_rshift_1_rg_a = MUX1HOT_v_32_4_2(accum_vector_data_13_sva,
      accum_vector_data_2_sva, accum_vector_data_8_sva, accum_vector_data_6_sva,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[2]) , (fsm_output[4])});
  wire PECore_RunBias_if_for_or_14_nl;
  wire [3:0] nl_PECore_RunBias_if_for_14_PECore_RunBias_if_for_rshift_1_rg_s;
  assign PECore_RunBias_if_for_or_14_nl = (fsm_output[4:2]!=3'b000);
  assign nl_PECore_RunBias_if_for_14_PECore_RunBias_if_for_rshift_1_rg_s = MUX_v_4_2_2(z_out_50,
      reg_PECore_RunMac_if_mux_122_ftd_1, PECore_RunBias_if_for_or_14_nl);
  wire [31:0] nl_PECore_RunBias_if_for_11_PECore_RunBias_if_for_rshift_1_rg_a;
  assign nl_PECore_RunBias_if_for_11_PECore_RunBias_if_for_rshift_1_rg_a = MUX1HOT_v_32_4_2(PECore_RunBias_if_accum_vector_out_data_lpi_1_dfm,
      PECore_RunBias_if_accum_vector_out_data_15_lpi_1_dfm, accum_vector_data_12_sva,
      PECore_RunBias_if_accum_vector_out_data_14_lpi_1_dfm, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[1]) , (fsm_output[3])});
  wire [3:0] nl_PECore_RunBias_if_for_11_PECore_RunBias_if_for_rshift_1_rg_s;
  assign nl_PECore_RunBias_if_for_11_PECore_RunBias_if_for_rshift_1_rg_s = MUX_v_4_2_2(reg_PECore_RunMac_if_mux_122_ftd_1,
      z_out_50, fsm_output[1]);
  wire [31:0] nl_PECore_RunBias_if_for_10_PECore_RunBias_if_for_rshift_1_rg_a;
  assign nl_PECore_RunBias_if_for_10_PECore_RunBias_if_for_rshift_1_rg_a = MUX1HOT_v_32_4_2(accum_vector_data_9_sva,
      accum_vector_data_14_sva, accum_vector_data_7_sva, accum_vector_data_4_sva,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])});
  wire [3:0] nl_PECore_RunBias_if_for_10_PECore_RunBias_if_for_rshift_1_rg_s;
  assign nl_PECore_RunBias_if_for_10_PECore_RunBias_if_for_rshift_1_rg_s = MUX_v_4_2_2(reg_PECore_RunMac_if_mux_122_ftd_1,
      z_out_50, fsm_output[1]);
  wire [31:0] nl_PECore_RunBias_if_for_16_PECore_RunBias_if_for_rshift_1_rg_a;
  assign nl_PECore_RunBias_if_for_16_PECore_RunBias_if_for_rshift_1_rg_a = MUX1HOT_v_32_4_2(PECore_RunBias_if_accum_vector_out_data_13_lpi_1_dfm,
      accum_vector_data_3_sva, accum_vector_data_5_sva, accum_vector_data_15_sva,
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[1])});
  wire [3:0] nl_PECore_RunBias_if_for_16_PECore_RunBias_if_for_rshift_1_rg_s;
  assign nl_PECore_RunBias_if_for_16_PECore_RunBias_if_for_rshift_1_rg_s = MUX_v_4_2_2(reg_PECore_RunMac_if_mux_122_ftd_1,
      z_out_50, fsm_output[1]);
  wire[3:0] adpfloat_tmp_to_fixed_20U_14U_mux1h_20_nl;
  wire [4:0] nl_PECore_RunBias_if_for_13_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_a;
  assign adpfloat_tmp_to_fixed_20U_14U_mux1h_20_nl = MUX1HOT_v_4_4_2((input_mem_banks_read_read_data_lpi_1[43:40]),
      (input_mem_banks_write_if_for_if_mux_cse[99:96]), (input_mem_banks_read_read_data_lpi_1[3:0]),
      (input_mem_banks_read_read_data_lpi_1[35:32]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4])});
  assign nl_PECore_RunBias_if_for_13_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_a =
      {1'b1 , adpfloat_tmp_to_fixed_20U_14U_mux1h_20_nl};
  wire[4:0] adpfloat_tmp_to_fixed_20U_14U_mux1h_13_nl;
  wire[4:0] PECore_RunBias_if_for_13_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_13_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_13_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_13_operator_33_true_acc_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_mux1h_21_nl;
  wire [5:0] nl_PECore_RunBias_if_for_13_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_s;
  assign nl_PECore_RunBias_if_for_13_operator_33_true_acc_nl = (operator_4_false_acc_psp_13_sva_1[3:1])
      + 3'b111;
  assign PECore_RunBias_if_for_13_operator_33_true_acc_nl = nl_PECore_RunBias_if_for_13_operator_33_true_acc_nl[2:0];
  assign nl_PECore_RunBias_if_for_13_operator_34_true_acc_nl = conv_s2s_4_5({PECore_RunBias_if_for_13_operator_33_true_acc_nl
      , (operator_4_false_acc_psp_13_sva_1[0])}) + 5'b00111;
  assign PECore_RunBias_if_for_13_operator_34_true_acc_nl = nl_PECore_RunBias_if_for_13_operator_34_true_acc_nl[4:0];
  assign adpfloat_tmp_to_fixed_20U_14U_mux1h_13_nl = MUX1HOT_v_5_4_2(reg_PECore_RunMac_if_mux_103_ftd_1,
      PECore_RunBias_if_for_13_operator_34_true_acc_nl, reg_PECore_RunMac_if_mux_14_ftd_1,
      reg_PECore_RunMac_if_mux_102_ftd_1, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4])});
  assign adpfloat_tmp_to_fixed_20U_14U_mux1h_21_nl = MUX1HOT_s_1_4_2(PECore_RunBias_if_for_6_operator_4_false_slc_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_0_itm,
      (z_out_50[0]), (reg_PECore_RunMac_if_mux_123_ftd_1[0]), (reg_PECore_RunMac_if_mux_127_ftd_1[0]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])});
  assign nl_PECore_RunBias_if_for_13_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_s =
      {adpfloat_tmp_to_fixed_20U_14U_mux1h_13_nl , adpfloat_tmp_to_fixed_20U_14U_mux1h_21_nl};
  wire[3:0] adpfloat_tmp_to_fixed_20U_14U_mux1h_22_nl;
  wire [4:0] nl_PECore_RunBias_if_for_16_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_a;
  assign adpfloat_tmp_to_fixed_20U_14U_mux1h_22_nl = MUX1HOT_v_4_4_2((input_mem_banks_read_read_data_lpi_1[51:48]),
      (input_mem_banks_write_if_for_if_mux_cse[123:120]), (input_mem_banks_read_read_data_lpi_1[59:56]),
      (input_mem_banks_read_read_data_lpi_1[11:8]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4])});
  assign nl_PECore_RunBias_if_for_16_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_a =
      {1'b1 , adpfloat_tmp_to_fixed_20U_14U_mux1h_22_nl};
  wire[4:0] adpfloat_tmp_to_fixed_20U_14U_mux1h_15_nl;
  wire[4:0] PECore_RunBias_if_for_16_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_16_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_16_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_16_operator_33_true_acc_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_mux1h_23_nl;
  wire [5:0] nl_PECore_RunBias_if_for_16_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_s;
  assign nl_PECore_RunBias_if_for_16_operator_33_true_acc_nl = (operator_4_false_acc_psp_sva_1[3:1])
      + 3'b111;
  assign PECore_RunBias_if_for_16_operator_33_true_acc_nl = nl_PECore_RunBias_if_for_16_operator_33_true_acc_nl[2:0];
  assign nl_PECore_RunBias_if_for_16_operator_34_true_acc_nl = conv_s2s_4_5({PECore_RunBias_if_for_16_operator_33_true_acc_nl
      , (operator_4_false_acc_psp_sva_1[0])}) + 5'b00111;
  assign PECore_RunBias_if_for_16_operator_34_true_acc_nl = nl_PECore_RunBias_if_for_16_operator_34_true_acc_nl[4:0];
  assign adpfloat_tmp_to_fixed_20U_14U_mux1h_15_nl = MUX1HOT_v_5_4_2(reg_PECore_RunMac_if_mux_104_ftd_1,
      PECore_RunBias_if_for_16_operator_34_true_acc_nl, (PECore_RunMac_if_mux_105_itm[4:0]),
      reg_PECore_RunMac_if_mux_141_ftd_1, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4])});
  assign adpfloat_tmp_to_fixed_20U_14U_mux1h_23_nl = MUX1HOT_s_1_4_2(PECore_RunBias_if_for_7_operator_4_false_slc_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_0_itm,
      (adpfloat_tmp_to_fixed_20U_14U_acc_sdt_sva_1[0]), (reg_PECore_RunMac_if_mux_128_ftd_1[0]),
      (reg_PECore_RunMac_if_mux_124_ftd_1[0]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4])});
  assign nl_PECore_RunBias_if_for_16_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_s =
      {adpfloat_tmp_to_fixed_20U_14U_mux1h_15_nl , adpfloat_tmp_to_fixed_20U_14U_mux1h_23_nl};
  wire[3:0] adpfloat_tmp_to_fixed_20U_14U_mux1h_24_nl;
  wire [4:0] nl_PECore_RunBias_if_for_10_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_a;
  assign adpfloat_tmp_to_fixed_20U_14U_mux1h_24_nl = MUX1HOT_v_4_4_2((input_mem_banks_read_read_data_lpi_1[75:72]),
      (input_mem_banks_write_if_for_if_mux_cse[115:112]), (input_mem_banks_read_read_data_lpi_1[67:64]),
      (input_mem_banks_read_read_data_lpi_1[19:16]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4])});
  assign nl_PECore_RunBias_if_for_10_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_a =
      {1'b1 , adpfloat_tmp_to_fixed_20U_14U_mux1h_24_nl};
  wire[4:0] adpfloat_tmp_to_fixed_20U_14U_mux1h_17_nl;
  wire[4:0] PECore_RunBias_if_for_15_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_15_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_15_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_15_operator_33_true_acc_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_mux1h_25_nl;
  wire [5:0] nl_PECore_RunBias_if_for_10_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_s;
  assign nl_PECore_RunBias_if_for_15_operator_33_true_acc_nl = (operator_4_false_acc_psp_15_sva_1[3:1])
      + 3'b111;
  assign PECore_RunBias_if_for_15_operator_33_true_acc_nl = nl_PECore_RunBias_if_for_15_operator_33_true_acc_nl[2:0];
  assign nl_PECore_RunBias_if_for_15_operator_34_true_acc_nl = conv_s2s_4_5({PECore_RunBias_if_for_15_operator_33_true_acc_nl
      , (operator_4_false_acc_psp_15_sva_1[0])}) + 5'b00111;
  assign PECore_RunBias_if_for_15_operator_34_true_acc_nl = nl_PECore_RunBias_if_for_15_operator_34_true_acc_nl[4:0];
  assign adpfloat_tmp_to_fixed_20U_14U_mux1h_17_nl = MUX1HOT_v_5_4_2(reg_PECore_RunMac_if_mux_100_ftd_1,
      PECore_RunBias_if_for_15_operator_34_true_acc_nl, (PECore_RunMac_if_mux_106_itm[4:0]),
      reg_PECore_RunMac_if_mux_1_ftd_1, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4])});
  assign adpfloat_tmp_to_fixed_20U_14U_mux1h_25_nl = MUX1HOT_s_1_4_2(PECore_RunBias_if_for_10_operator_4_false_slc_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_0_itm,
      (adpfloat_tmp_to_fixed_20U_14U_acc_sdt_15_sva_1[0]), (reg_PECore_RunMac_if_mux_129_ftd_1[0]),
      (reg_PECore_RunMac_if_mux_125_ftd_1[0]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4])});
  assign nl_PECore_RunBias_if_for_10_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_s =
      {adpfloat_tmp_to_fixed_20U_14U_mux1h_17_nl , adpfloat_tmp_to_fixed_20U_14U_mux1h_25_nl};
  wire[3:0] adpfloat_tmp_to_fixed_20U_14U_mux1h_26_nl;
  wire [4:0] nl_PECore_RunBias_if_for_11_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_a;
  assign adpfloat_tmp_to_fixed_20U_14U_mux1h_26_nl = MUX1HOT_v_4_4_2((input_mem_banks_read_read_data_lpi_1[83:80]),
      (input_mem_banks_write_if_for_if_mux_cse[107:104]), (input_mem_banks_read_read_data_lpi_1[91:88]),
      (input_mem_banks_read_read_data_lpi_1[27:24]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4])});
  assign nl_PECore_RunBias_if_for_11_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_a =
      {1'b1 , adpfloat_tmp_to_fixed_20U_14U_mux1h_26_nl};
  wire[4:0] adpfloat_tmp_to_fixed_20U_14U_mux1h_19_nl;
  wire[4:0] PECore_RunBias_if_for_14_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_14_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_14_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_14_operator_33_true_acc_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_mux1h_27_nl;
  wire [5:0] nl_PECore_RunBias_if_for_11_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_s;
  assign nl_PECore_RunBias_if_for_14_operator_33_true_acc_nl = (operator_4_false_acc_psp_14_sva_1[3:1])
      + 3'b111;
  assign PECore_RunBias_if_for_14_operator_33_true_acc_nl = nl_PECore_RunBias_if_for_14_operator_33_true_acc_nl[2:0];
  assign nl_PECore_RunBias_if_for_14_operator_34_true_acc_nl = conv_s2s_4_5({PECore_RunBias_if_for_14_operator_33_true_acc_nl
      , (operator_4_false_acc_psp_14_sva_1[0])}) + 5'b00111;
  assign PECore_RunBias_if_for_14_operator_34_true_acc_nl = nl_PECore_RunBias_if_for_14_operator_34_true_acc_nl[4:0];
  assign adpfloat_tmp_to_fixed_20U_14U_mux1h_19_nl = MUX1HOT_v_5_4_2(reg_PECore_RunMac_if_mux_101_ftd_1,
      PECore_RunBias_if_for_14_operator_34_true_acc_nl, reg_PECore_RunMac_if_mux_138_ftd_1,
      reg_PECore_RunMac_if_mux_10_ftd_1, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4])});
  assign adpfloat_tmp_to_fixed_20U_14U_mux1h_27_nl = MUX1HOT_s_1_4_2(PECore_RunBias_if_for_11_operator_4_false_slc_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_0_itm,
      (adpfloat_tmp_to_fixed_20U_14U_acc_sdt_14_sva_1[0]), (reg_PECore_RunMac_if_mux_11_ftd_1[0]),
      (reg_PECore_RunMac_if_mux_126_ftd_1[0]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4])});
  assign nl_PECore_RunBias_if_for_11_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_s =
      {adpfloat_tmp_to_fixed_20U_14U_mux1h_19_nl , adpfloat_tmp_to_fixed_20U_14U_mux1h_27_nl};
  wire [319:0] nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_idat;
  assign nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_idat = {act_port_Push_mioi_idat_319_300
      , act_port_Push_mioi_idat_299_280 , act_port_Push_mioi_idat_279_260 , act_port_Push_mioi_idat_259_240
      , act_port_Push_mioi_idat_239_220 , act_port_Push_mioi_idat_219_200 , act_port_Push_mioi_idat_199_180
      , act_port_Push_mioi_idat_179_160 , act_port_Push_mioi_idat_159_140 , act_port_Push_mioi_idat_139_120
      , act_port_Push_mioi_idat_119_100 , act_port_Push_mioi_idat_99_80 , act_port_Push_mioi_idat_79_60
      , act_port_Push_mioi_idat_59_40 , act_port_Push_mioi_idat_39_20 , act_port_Push_mioi_idat_19_0};
  wire [127:0] nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_idat;
  assign nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_idat = {rva_out_Push_mioi_idat_127_120
      , rva_out_Push_mioi_idat_119_112 , rva_out_Push_mioi_idat_111_104 , rva_out_Push_mioi_idat_103_96
      , rva_out_Push_mioi_idat_95_88 , rva_out_Push_mioi_idat_87_80 , rva_out_Push_mioi_idat_79_72
      , rva_out_Push_mioi_idat_71_64 , rva_out_Push_mioi_idat_63_56 , rva_out_Push_mioi_idat_55_48
      , rva_out_Push_mioi_idat_47_40 , rva_out_Push_mioi_idat_39_36 , rva_out_Push_mioi_idat_35_32
      , rva_out_Push_mioi_idat_31_27 , rva_out_Push_mioi_idat_26_25 , rva_out_Push_mioi_idat_24
      , rva_out_Push_mioi_idat_23_19 , rva_out_Push_mioi_idat_18_17 , rva_out_Push_mioi_idat_16
      , rva_out_Push_mioi_idat_15_11 , rva_out_Push_mioi_idat_10_9 , rva_out_Push_mioi_idat_8
      , rva_out_Push_mioi_idat_7_1 , rva_out_Push_mioi_idat_0};
  PECore_ProductSum  Datapath_for_1_ProductSum_cmp (
      .in_1_data_rsc_dat(nl_Datapath_for_1_ProductSum_cmp_in_1_data_rsc_dat[127:0]),
      .in_2_data_rsc_dat(input_mem_banks_read_read_data_mux_rmff),
      .out_rsc_z(Datapath_for_1_ProductSum_cmp_out_rsc_z),
      .ccs_ccore_start_rsc_dat(or_2419_rmff),
      .ccs_ccore_clk(clk),
      .ccs_ccore_arst(rst),
      .ccs_ccore_en(Datapath_for_1_ProductSum_cmp_ccs_ccore_en)
    );
  PECore_ProductSum  Datapath_for_1_ProductSum_cmp_1 (
      .in_1_data_rsc_dat(nl_Datapath_for_1_ProductSum_cmp_1_in_1_data_rsc_dat[127:0]),
      .in_2_data_rsc_dat(input_mem_banks_read_read_data_mux_rmff),
      .out_rsc_z(Datapath_for_1_ProductSum_cmp_1_out_rsc_z),
      .ccs_ccore_start_rsc_dat(or_2419_rmff),
      .ccs_ccore_clk(clk),
      .ccs_ccore_arst(rst),
      .ccs_ccore_en(Datapath_for_1_ProductSum_cmp_ccs_ccore_en)
    );
  PECore_ProductSum  Datapath_for_1_ProductSum_cmp_2 (
      .in_1_data_rsc_dat(nl_Datapath_for_1_ProductSum_cmp_2_in_1_data_rsc_dat[127:0]),
      .in_2_data_rsc_dat(input_mem_banks_read_read_data_mux_rmff),
      .out_rsc_z(Datapath_for_1_ProductSum_cmp_2_out_rsc_z),
      .ccs_ccore_start_rsc_dat(or_2419_rmff),
      .ccs_ccore_clk(clk),
      .ccs_ccore_arst(rst),
      .ccs_ccore_en(Datapath_for_1_ProductSum_cmp_ccs_ccore_en)
    );
  PECore_ProductSum  Datapath_for_1_ProductSum_cmp_3 (
      .in_1_data_rsc_dat(nl_Datapath_for_1_ProductSum_cmp_3_in_1_data_rsc_dat[127:0]),
      .in_2_data_rsc_dat(input_mem_banks_read_read_data_mux_rmff),
      .out_rsc_z(Datapath_for_1_ProductSum_cmp_3_out_rsc_z),
      .ccs_ccore_start_rsc_dat(or_2419_rmff),
      .ccs_ccore_clk(clk),
      .ccs_ccore_arst(rst),
      .ccs_ccore_en(Datapath_for_1_ProductSum_cmp_ccs_ccore_en)
    );
  PECore_mgc_muladd1 #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_cst(32'sd1),
  .signd_cst(32'sd0),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd13),
  .add_axb(32'sd1),
  .add_c(32'sd1),
  .add_d(32'sd1),
  .use_const(32'sd1)) PEManager_16U_GetWeightAddr_if_acc_4_cmp (
      .a(nl_PEManager_16U_GetWeightAddr_if_acc_4_cmp_a[7:0]),
      .b(nl_PEManager_16U_GetWeightAddr_if_acc_4_cmp_b[7:0]),
      .c(nl_PEManager_16U_GetWeightAddr_if_acc_4_cmp_c[7:0]),
      .cst(1'b0),
      .z(PEManager_16U_GetWeightAddr_if_acc_4_cmp_z)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd16)) weight_mem_write_arbxbar_xbar_for_lshift_rg (
      .a(nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a),
      .s(nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s[3:0]),
      .z(weight_mem_write_arbxbar_xbar_for_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd16)) weight_mem_read_arbxbar_xbar_for_15_lshift_rg (
      .a(weight_read_req_valid_8_lpi_1_dfm_1),
      .s(nl_weight_mem_read_arbxbar_xbar_for_15_lshift_rg_s[3:0]),
      .z(weight_mem_read_arbxbar_xbar_for_15_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd16)) weight_mem_read_arbxbar_xbar_for_1_lshift_rg (
      .a(weight_read_req_valid_0_lpi_1_dfm_4_mx0),
      .s(nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s[3:0]),
      .z(weight_mem_read_arbxbar_xbar_for_1_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd16)) weight_mem_read_arbxbar_xbar_for_11_lshift_rg (
      .a(weight_read_req_valid_8_lpi_1_dfm_1),
      .s(nl_weight_mem_read_arbxbar_xbar_for_11_lshift_rg_s[3:0]),
      .z(weight_mem_read_arbxbar_xbar_for_11_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd16)) weight_mem_read_arbxbar_xbar_for_13_lshift_rg (
      .a(weight_read_req_valid_8_lpi_1_dfm_1),
      .s(nl_weight_mem_read_arbxbar_xbar_for_13_lshift_rg_s[3:0]),
      .z(weight_mem_read_arbxbar_xbar_for_13_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd16)) weight_mem_read_arbxbar_xbar_for_16_lshift_rg (
      .a(weight_read_req_valid_8_lpi_1_dfm_1),
      .s(nl_weight_mem_read_arbxbar_xbar_for_16_lshift_rg_s[3:0]),
      .z(weight_mem_read_arbxbar_xbar_for_16_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd16)) weight_mem_read_arbxbar_xbar_for_12_lshift_rg (
      .a(weight_read_req_valid_8_lpi_1_dfm_1),
      .s(nl_weight_mem_read_arbxbar_xbar_for_12_lshift_rg_s[3:0]),
      .z(weight_mem_read_arbxbar_xbar_for_12_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd16)) weight_mem_read_arbxbar_xbar_for_14_lshift_rg (
      .a(weight_read_req_valid_8_lpi_1_dfm_1),
      .s(nl_weight_mem_read_arbxbar_xbar_for_14_lshift_rg_s[3:0]),
      .z(weight_mem_read_arbxbar_xbar_for_14_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd16)) weight_mem_read_arbxbar_xbar_for_7_lshift_rg (
      .a(PECore_RunFSM_switch_lp_equal_tmp_5),
      .s(nl_weight_mem_read_arbxbar_xbar_for_7_lshift_rg_s[3:0]),
      .z(weight_mem_read_arbxbar_xbar_for_7_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd16)) weight_mem_read_arbxbar_xbar_for_9_lshift_rg (
      .a(weight_read_req_valid_8_lpi_1_dfm_1),
      .s(nl_weight_mem_read_arbxbar_xbar_for_9_lshift_rg_s[3:0]),
      .z(weight_mem_read_arbxbar_xbar_for_9_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd16)) weight_mem_read_arbxbar_xbar_for_3_lshift_rg (
      .a(PECore_RunFSM_switch_lp_equal_tmp_5),
      .s(nl_weight_mem_read_arbxbar_xbar_for_3_lshift_rg_s[3:0]),
      .z(weight_mem_read_arbxbar_xbar_for_3_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd16)) weight_mem_read_arbxbar_xbar_for_5_lshift_rg (
      .a(PECore_RunFSM_switch_lp_equal_tmp_5),
      .s(nl_weight_mem_read_arbxbar_xbar_for_5_lshift_rg_s[3:0]),
      .z(weight_mem_read_arbxbar_xbar_for_5_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd16)) weight_mem_read_arbxbar_xbar_for_8_lshift_rg (
      .a(PECore_RunFSM_switch_lp_equal_tmp_5),
      .s(nl_weight_mem_read_arbxbar_xbar_for_8_lshift_rg_s[3:0]),
      .z(weight_mem_read_arbxbar_xbar_for_8_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd16)) weight_mem_read_arbxbar_xbar_for_4_lshift_rg (
      .a(PECore_RunFSM_switch_lp_equal_tmp_5),
      .s(nl_weight_mem_read_arbxbar_xbar_for_4_lshift_rg_s[3:0]),
      .z(weight_mem_read_arbxbar_xbar_for_4_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd16)) weight_mem_read_arbxbar_xbar_for_6_lshift_rg (
      .a(PECore_RunFSM_switch_lp_equal_tmp_5),
      .s(nl_weight_mem_read_arbxbar_xbar_for_6_lshift_rg_s[3:0]),
      .z(weight_mem_read_arbxbar_xbar_for_6_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd16)) weight_mem_read_arbxbar_xbar_for_10_lshift_rg (
      .a(weight_read_req_valid_8_lpi_1_dfm_1),
      .s(nl_weight_mem_read_arbxbar_xbar_for_10_lshift_rg_s[3:0]),
      .z(weight_mem_read_arbxbar_xbar_for_10_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd16)) weight_mem_read_arbxbar_xbar_for_2_lshift_rg (
      .a(PECore_RunFSM_switch_lp_equal_tmp_5),
      .s(nl_weight_mem_read_arbxbar_xbar_for_2_lshift_rg_s[3:0]),
      .z(weight_mem_read_arbxbar_xbar_for_2_lshift_tmp)
    );
  PECore_mgc_shift_r_v5 #(.width_a(32'sd32),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd32)) PECore_RunBias_if_for_14_PECore_RunBias_if_for_rshift_1_rg (
      .a(nl_PECore_RunBias_if_for_14_PECore_RunBias_if_for_rshift_1_rg_a[31:0]),
      .s(nl_PECore_RunBias_if_for_14_PECore_RunBias_if_for_rshift_1_rg_s[3:0]),
      .z(z_out_37)
    );
  PECore_mgc_shift_r_v5 #(.width_a(32'sd32),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd32)) PECore_RunBias_if_for_11_PECore_RunBias_if_for_rshift_1_rg (
      .a(nl_PECore_RunBias_if_for_11_PECore_RunBias_if_for_rshift_1_rg_a[31:0]),
      .s(nl_PECore_RunBias_if_for_11_PECore_RunBias_if_for_rshift_1_rg_s[3:0]),
      .z(z_out_38)
    );
  PECore_mgc_shift_r_v5 #(.width_a(32'sd32),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd32)) PECore_RunBias_if_for_10_PECore_RunBias_if_for_rshift_1_rg (
      .a(nl_PECore_RunBias_if_for_10_PECore_RunBias_if_for_rshift_1_rg_a[31:0]),
      .s(nl_PECore_RunBias_if_for_10_PECore_RunBias_if_for_rshift_1_rg_s[3:0]),
      .z(z_out_39)
    );
  PECore_mgc_shift_r_v5 #(.width_a(32'sd32),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd32)) PECore_RunBias_if_for_16_PECore_RunBias_if_for_rshift_1_rg (
      .a(nl_PECore_RunBias_if_for_16_PECore_RunBias_if_for_rshift_1_rg_a[31:0]),
      .s(nl_PECore_RunBias_if_for_16_PECore_RunBias_if_for_rshift_1_rg_s[3:0]),
      .z(z_out_40)
    );
  PECore_mgc_shift_bl_v5 #(.width_a(32'sd5),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd20)) PECore_RunBias_if_for_13_adpfloat_tmp_to_fixed_20U_14U_lshift_rg
      (
      .a(nl_PECore_RunBias_if_for_13_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_a[4:0]),
      .s(nl_PECore_RunBias_if_for_13_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_s[5:0]),
      .z(z_out_46)
    );
  PECore_mgc_shift_bl_v5 #(.width_a(32'sd5),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd20)) PECore_RunBias_if_for_16_adpfloat_tmp_to_fixed_20U_14U_lshift_rg
      (
      .a(nl_PECore_RunBias_if_for_16_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_a[4:0]),
      .s(nl_PECore_RunBias_if_for_16_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_s[5:0]),
      .z(z_out_47)
    );
  PECore_mgc_shift_bl_v5 #(.width_a(32'sd5),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd20)) PECore_RunBias_if_for_10_adpfloat_tmp_to_fixed_20U_14U_lshift_rg
      (
      .a(nl_PECore_RunBias_if_for_10_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_a[4:0]),
      .s(nl_PECore_RunBias_if_for_10_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_s[5:0]),
      .z(z_out_48)
    );
  PECore_mgc_shift_bl_v5 #(.width_a(32'sd5),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd20)) PECore_RunBias_if_for_11_adpfloat_tmp_to_fixed_20U_14U_lshift_rg
      (
      .a(nl_PECore_RunBias_if_for_11_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_a[4:0]),
      .s(nl_PECore_RunBias_if_for_11_adpfloat_tmp_to_fixed_20U_14U_lshift_rg_s[5:0]),
      .z(z_out_49)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi PECore_PECoreRun_input_port_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .input_port_val(input_port_val),
      .input_port_rdy(input_port_rdy),
      .input_port_msg(input_port_msg),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .input_port_PopNB_mioi_oswt(reg_input_port_PopNB_mioi_oswt_cse),
      .input_port_PopNB_mioi_idat_mxwt(input_port_PopNB_mioi_idat_mxwt),
      .input_port_PopNB_mioi_ivld_mxwt(input_port_PopNB_mioi_ivld_mxwt)
    );
  PECore_PECore_PECoreRun_wait_dp PECore_PECoreRun_wait_dp_inst (
      .weight_mem_banks_bank_array_impl_data0_rsci_clken_d(weight_mem_banks_bank_array_impl_data0_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data1_rsci_clken_d(weight_mem_banks_bank_array_impl_data1_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data2_rsci_clken_d(weight_mem_banks_bank_array_impl_data2_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data3_rsci_clken_d(weight_mem_banks_bank_array_impl_data3_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data4_rsci_clken_d(weight_mem_banks_bank_array_impl_data4_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data5_rsci_clken_d(weight_mem_banks_bank_array_impl_data5_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data6_rsci_clken_d(weight_mem_banks_bank_array_impl_data6_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data7_rsci_clken_d(weight_mem_banks_bank_array_impl_data7_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data8_rsci_clken_d(weight_mem_banks_bank_array_impl_data8_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data9_rsci_clken_d(weight_mem_banks_bank_array_impl_data9_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data10_rsci_clken_d(weight_mem_banks_bank_array_impl_data10_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data11_rsci_clken_d(weight_mem_banks_bank_array_impl_data11_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data12_rsci_clken_d(weight_mem_banks_bank_array_impl_data12_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data13_rsci_clken_d(weight_mem_banks_bank_array_impl_data13_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data14_rsci_clken_d(weight_mem_banks_bank_array_impl_data14_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data15_rsci_clken_d(weight_mem_banks_bank_array_impl_data15_rsci_clken_d),
      .input_mem_banks_bank_array_impl_data0_rsci_clken_d(input_mem_banks_bank_array_impl_data0_rsci_clken_d),
      .PECoreRun_wen(PECoreRun_wen),
      .weight_mem_banks_bank_array_impl_data0_rsci_cgo(reg_weight_mem_banks_bank_array_impl_data0_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_array_impl_data0_rsci_cgo_ir_unreg(or_2438_rmff),
      .weight_mem_banks_bank_array_impl_data1_rsci_cgo(reg_weight_mem_banks_bank_array_impl_data1_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_array_impl_data1_rsci_cgo_ir_unreg(or_2437_rmff),
      .weight_mem_banks_bank_array_impl_data2_rsci_cgo(reg_weight_mem_banks_bank_array_impl_data2_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_array_impl_data2_rsci_cgo_ir_unreg(or_2436_rmff),
      .weight_mem_banks_bank_array_impl_data3_rsci_cgo(reg_weight_mem_banks_bank_array_impl_data3_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_array_impl_data3_rsci_cgo_ir_unreg(or_2435_rmff),
      .weight_mem_banks_bank_array_impl_data4_rsci_cgo(reg_weight_mem_banks_bank_array_impl_data4_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_array_impl_data4_rsci_cgo_ir_unreg(or_2434_rmff),
      .weight_mem_banks_bank_array_impl_data5_rsci_cgo(reg_weight_mem_banks_bank_array_impl_data5_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_array_impl_data5_rsci_cgo_ir_unreg(or_2433_rmff),
      .weight_mem_banks_bank_array_impl_data6_rsci_cgo(reg_weight_mem_banks_bank_array_impl_data6_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_array_impl_data6_rsci_cgo_ir_unreg(or_2432_rmff),
      .weight_mem_banks_bank_array_impl_data7_rsci_cgo(reg_weight_mem_banks_bank_array_impl_data7_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_array_impl_data7_rsci_cgo_ir_unreg(or_2431_rmff),
      .weight_mem_banks_bank_array_impl_data8_rsci_cgo(reg_weight_mem_banks_bank_array_impl_data8_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_array_impl_data8_rsci_cgo_ir_unreg(or_2430_rmff),
      .weight_mem_banks_bank_array_impl_data9_rsci_cgo(reg_weight_mem_banks_bank_array_impl_data9_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_array_impl_data9_rsci_cgo_ir_unreg(or_2429_rmff),
      .weight_mem_banks_bank_array_impl_data10_rsci_cgo(reg_weight_mem_banks_bank_array_impl_data10_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_array_impl_data10_rsci_cgo_ir_unreg(or_2428_rmff),
      .weight_mem_banks_bank_array_impl_data11_rsci_cgo(reg_weight_mem_banks_bank_array_impl_data11_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_array_impl_data11_rsci_cgo_ir_unreg(or_2427_rmff),
      .weight_mem_banks_bank_array_impl_data12_rsci_cgo(reg_weight_mem_banks_bank_array_impl_data12_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_array_impl_data12_rsci_cgo_ir_unreg(or_2426_rmff),
      .weight_mem_banks_bank_array_impl_data13_rsci_cgo(reg_weight_mem_banks_bank_array_impl_data13_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_array_impl_data13_rsci_cgo_ir_unreg(or_2425_rmff),
      .weight_mem_banks_bank_array_impl_data14_rsci_cgo(reg_weight_mem_banks_bank_array_impl_data14_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_array_impl_data14_rsci_cgo_ir_unreg(or_2424_rmff),
      .weight_mem_banks_bank_array_impl_data15_rsci_cgo(reg_weight_mem_banks_bank_array_impl_data15_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_array_impl_data15_rsci_cgo_ir_unreg(or_2423_rmff),
      .input_mem_banks_bank_array_impl_data0_rsci_cgo(reg_input_mem_banks_bank_array_impl_data0_rsci_cgo_ir_cse),
      .input_mem_banks_bank_array_impl_data0_rsci_cgo_ir_unreg(or_2422_rmff),
      .Datapath_for_1_ProductSum_cmp_cgo(reg_Datapath_for_1_ProductSum_cmp_cgo_ir_3_cse),
      .Datapath_for_1_ProductSum_cmp_cgo_ir_unreg(or_2421_rmff),
      .Datapath_for_1_ProductSum_cmp_ccs_ccore_en(Datapath_for_1_ProductSum_cmp_ccs_ccore_en)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi PECore_PECoreRun_rva_in_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_val(rva_in_val),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_msg(rva_in_msg),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .rva_in_PopNB_mioi_oswt(reg_rva_in_PopNB_mioi_oswt_cse),
      .rva_in_PopNB_mioi_idat_mxwt(rva_in_PopNB_mioi_idat_mxwt),
      .rva_in_PopNB_mioi_ivld_mxwt(rva_in_PopNB_mioi_ivld_mxwt)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi PECore_PECoreRun_act_port_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .act_port_val(act_port_val),
      .act_port_rdy(act_port_rdy),
      .act_port_msg(act_port_msg),
      .PECoreRun_wen(PECoreRun_wen),
      .act_port_Push_mioi_oswt(reg_act_port_Push_mioi_iswt0_cse),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .act_port_Push_mioi_idat(nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_idat[319:0])
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi PECore_PECoreRun_rva_out_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_val(rva_out_val),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_msg(rva_out_msg),
      .PECoreRun_wen(PECoreRun_wen),
      .rva_out_Push_mioi_oswt(reg_rva_out_Push_mioi_iswt0_cse),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_idat(nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_idat[127:0])
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi PECore_PECoreRun_start_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .start_val(start_val),
      .start_rdy(start_rdy),
      .start_msg(start_msg),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .start_PopNB_mioi_oswt(reg_start_PopNB_mioi_iswt0_cse),
      .start_PopNB_mioi_idat_mxwt(start_PopNB_mioi_idat_mxwt),
      .start_PopNB_mioi_ivld_mxwt(start_PopNB_mioi_ivld_mxwt)
    );
  PECore_PECore_PECoreRun_staller PECore_PECoreRun_staller_inst (
      .clk(clk),
      .rst(rst),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp)
    );
  PECore_PECore_PECoreRun_PECoreRun_fsm PECore_PECoreRun_PECoreRun_fsm_inst (
      .clk(clk),
      .rst(rst),
      .PECoreRun_wen(PECoreRun_wen),
      .fsm_output(fsm_output)
    );
  assign weight_mem_banks_write_if_for_if_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_3039_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb = weight_mem_banks_write_if_for_if_mux_cse;
  assign weight_mem_banks_write_if_for_if_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_3039_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb = weight_mem_banks_write_if_for_if_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb = weight_mem_banks_write_if_for_if_mux_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb = weight_mem_banks_write_if_for_if_mux_1_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb
      = weight_mem_banks_write_if_for_if_mux_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb
      = weight_mem_banks_write_if_for_if_mux_1_cse;
  assign weight_mem_banks_read_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, or_1405_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 = weight_mem_banks_read_for_mux_cse;
  assign weight_mem_banks_read_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, or_1405_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1 = weight_mem_banks_read_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 = weight_mem_banks_read_for_mux_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1 = weight_mem_banks_read_for_mux_1_cse;
  assign weight_mem_banks_write_if_for_if_mux_4_cse = MUX1HOT_s_1_1_2(1'b1, and_3035_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2 = weight_mem_banks_write_if_for_if_mux_4_cse;
  assign weight_mem_banks_write_if_for_if_mux_5_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_3035_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2 = weight_mem_banks_write_if_for_if_mux_5_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2 = weight_mem_banks_write_if_for_if_mux_4_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2 = weight_mem_banks_write_if_for_if_mux_5_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1
      = weight_mem_banks_write_if_for_if_mux_4_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1
      = weight_mem_banks_write_if_for_if_mux_5_cse;
  assign weight_mem_banks_read_for_mux_4_cse = MUX1HOT_s_1_1_2(1'b1, or_1409_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3 = weight_mem_banks_read_for_mux_4_cse;
  assign weight_mem_banks_read_for_mux_5_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, or_1409_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3 = weight_mem_banks_read_for_mux_5_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3 = weight_mem_banks_read_for_mux_4_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3 = weight_mem_banks_read_for_mux_5_cse;
  assign weight_mem_banks_write_if_for_if_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_3031_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4 = weight_mem_banks_write_if_for_if_mux_8_cse;
  assign weight_mem_banks_write_if_for_if_mux_9_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_3031_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4 = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4 = weight_mem_banks_write_if_for_if_mux_8_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4 = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2
      = weight_mem_banks_write_if_for_if_mux_8_cse;
   assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2
      = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign weight_mem_banks_read_for_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, or_1413_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5 = weight_mem_banks_read_for_mux_8_cse;
  assign weight_mem_banks_read_for_mux_9_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, or_1413_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5 = weight_mem_banks_read_for_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5 = weight_mem_banks_read_for_mux_8_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5 = weight_mem_banks_read_for_mux_9_cse;
  assign weight_mem_banks_write_if_for_if_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_3027_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6 = weight_mem_banks_write_if_for_if_mux_12_cse;
  assign weight_mem_banks_write_if_for_if_mux_13_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_3027_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6 = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6 = weight_mem_banks_write_if_for_if_mux_12_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6 = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3
      = weight_mem_banks_write_if_for_if_mux_12_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3
      = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign weight_mem_banks_read_for_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, or_1417_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7 = weight_mem_banks_read_for_mux_12_cse;
  assign weight_mem_banks_read_for_mux_13_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, or_1417_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7 = weight_mem_banks_read_for_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7 = weight_mem_banks_read_for_mux_12_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7 = weight_mem_banks_read_for_mux_13_cse;
  assign weight_mem_banks_write_if_for_if_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_3023_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8 = weight_mem_banks_write_if_for_if_mux_16_cse;
  assign weight_mem_banks_write_if_for_if_mux_17_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_3023_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8 = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8 = weight_mem_banks_write_if_for_if_mux_16_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8 = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4
      = weight_mem_banks_write_if_for_if_mux_16_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4
      = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign weight_mem_banks_read_for_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, or_1421_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9 = weight_mem_banks_read_for_mux_16_cse;
  assign weight_mem_banks_read_for_mux_17_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, or_1421_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9 = weight_mem_banks_read_for_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9 = weight_mem_banks_read_for_mux_16_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9 = weight_mem_banks_read_for_mux_17_cse;
  assign weight_mem_banks_write_if_for_if_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_3019_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10 = weight_mem_banks_write_if_for_if_mux_20_cse;
  assign weight_mem_banks_write_if_for_if_mux_21_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_3019_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10 = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10 = weight_mem_banks_write_if_for_if_mux_20_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10 = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5
      = weight_mem_banks_write_if_for_if_mux_20_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5
      = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign weight_mem_banks_read_for_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, or_1425_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11 = weight_mem_banks_read_for_mux_20_cse;
  assign weight_mem_banks_read_for_mux_21_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, or_1425_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11 = weight_mem_banks_read_for_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11 = weight_mem_banks_read_for_mux_20_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11 = weight_mem_banks_read_for_mux_21_cse;
  assign weight_mem_banks_write_if_for_if_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_3015_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12 = weight_mem_banks_write_if_for_if_mux_24_cse;
  assign weight_mem_banks_write_if_for_if_mux_25_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_3015_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12 = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12 = weight_mem_banks_write_if_for_if_mux_24_cse;
   assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12 = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6
      = weight_mem_banks_write_if_for_if_mux_24_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6
      = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign weight_mem_banks_read_for_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, or_1429_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13 = weight_mem_banks_read_for_mux_24_cse;
  assign weight_mem_banks_read_for_mux_25_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, or_1429_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13 = weight_mem_banks_read_for_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13 = weight_mem_banks_read_for_mux_24_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13 = weight_mem_banks_read_for_mux_25_cse;
  assign weight_mem_banks_write_if_for_if_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_3011_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14 = weight_mem_banks_write_if_for_if_mux_28_cse;
  assign weight_mem_banks_write_if_for_if_mux_29_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_3011_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14 = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14 = weight_mem_banks_write_if_for_if_mux_28_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14 = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7
      = weight_mem_banks_write_if_for_if_mux_28_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7
      = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign weight_mem_banks_read_for_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, or_1433_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15 = weight_mem_banks_read_for_mux_28_cse;
  assign weight_mem_banks_read_for_mux_29_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, or_1433_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15 = weight_mem_banks_read_for_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15 = weight_mem_banks_read_for_mux_28_cse;
   assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15 = weight_mem_banks_read_for_mux_29_cse;
  assign weight_mem_banks_write_if_for_if_mux_32_cse = MUX1HOT_s_1_1_2(1'b1, and_3007_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16 = weight_mem_banks_write_if_for_if_mux_32_cse;
  assign weight_mem_banks_write_if_for_if_mux_33_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_3007_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16 = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16 = weight_mem_banks_write_if_for_if_mux_32_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16 = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8
      = weight_mem_banks_write_if_for_if_mux_32_cse;
   assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8
      = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign weight_mem_banks_read_for_mux_32_cse = MUX1HOT_s_1_1_2(1'b1, or_1437_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17 = weight_mem_banks_read_for_mux_32_cse;
  assign weight_mem_banks_read_for_mux_33_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, or_1437_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17 = weight_mem_banks_read_for_mux_33_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17 = weight_mem_banks_read_for_mux_32_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17 = weight_mem_banks_read_for_mux_33_cse;
  assign weight_mem_banks_write_if_for_if_mux_36_cse = MUX1HOT_s_1_1_2(1'b1, and_3003_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18 = weight_mem_banks_write_if_for_if_mux_36_cse;
  assign weight_mem_banks_write_if_for_if_mux_37_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_3003_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18 = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18 = weight_mem_banks_write_if_for_if_mux_36_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18 = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9
      = weight_mem_banks_write_if_for_if_mux_36_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9
      = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign weight_mem_banks_read_for_mux_36_cse = MUX1HOT_s_1_1_2(1'b1, or_1441_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19 = weight_mem_banks_read_for_mux_36_cse;
  assign weight_mem_banks_read_for_mux_37_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, or_1441_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19 = weight_mem_banks_read_for_mux_37_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19 = weight_mem_banks_read_for_mux_36_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19 = weight_mem_banks_read_for_mux_37_cse;
  assign weight_mem_banks_write_if_for_if_mux_40_cse = MUX1HOT_s_1_1_2(1'b1, and_2999_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20 = weight_mem_banks_write_if_for_if_mux_40_cse;
  assign weight_mem_banks_write_if_for_if_mux_41_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_2999_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20 = weight_mem_banks_write_if_for_if_mux_41_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20 = weight_mem_banks_write_if_for_if_mux_40_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20 = weight_mem_banks_write_if_for_if_mux_41_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_10
      = weight_mem_banks_write_if_for_if_mux_40_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_10
      = weight_mem_banks_write_if_for_if_mux_41_cse;
  assign weight_mem_banks_read_for_mux_40_cse = MUX1HOT_s_1_1_2(1'b1, or_1445_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21 = weight_mem_banks_read_for_mux_40_cse;
  assign weight_mem_banks_read_for_mux_41_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, or_1445_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21 = weight_mem_banks_read_for_mux_41_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21 = weight_mem_banks_read_for_mux_40_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21 = weight_mem_banks_read_for_mux_41_cse;
  assign weight_mem_banks_write_if_for_if_mux_44_cse = MUX1HOT_s_1_1_2(1'b1, and_2995_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22 = weight_mem_banks_write_if_for_if_mux_44_cse;
   assign weight_mem_banks_write_if_for_if_mux_45_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_2995_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22 = weight_mem_banks_write_if_for_if_mux_45_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22 = weight_mem_banks_write_if_for_if_mux_44_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22 = weight_mem_banks_write_if_for_if_mux_45_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_11
      = weight_mem_banks_write_if_for_if_mux_44_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_11
      = weight_mem_banks_write_if_for_if_mux_45_cse;
  assign weight_mem_banks_read_for_mux_44_cse = MUX1HOT_s_1_1_2(1'b1, or_1449_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23 = weight_mem_banks_read_for_mux_44_cse;
  assign weight_mem_banks_read_for_mux_45_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, or_1449_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23 = weight_mem_banks_read_for_mux_45_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23 = weight_mem_banks_read_for_mux_44_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23 = weight_mem_banks_read_for_mux_45_cse;
  assign weight_mem_banks_write_if_for_if_mux_48_cse = MUX1HOT_s_1_1_2(1'b1, and_2991_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24 = weight_mem_banks_write_if_for_if_mux_48_cse;
  assign weight_mem_banks_write_if_for_if_mux_49_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_2991_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24 = weight_mem_banks_write_if_for_if_mux_49_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24 = weight_mem_banks_write_if_for_if_mux_48_cse;
 assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24 = weight_mem_banks_write_if_for_if_mux_49_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_12
      = weight_mem_banks_write_if_for_if_mux_48_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_12
      = weight_mem_banks_write_if_for_if_mux_49_cse;
  assign weight_mem_banks_read_for_mux_48_cse = MUX1HOT_s_1_1_2(1'b1, or_1453_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25 = weight_mem_banks_read_for_mux_48_cse;
  assign weight_mem_banks_read_for_mux_49_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, or_1453_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25 = weight_mem_banks_read_for_mux_49_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25 = weight_mem_banks_read_for_mux_48_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25 = weight_mem_banks_read_for_mux_49_cse;
  assign weight_mem_banks_write_if_for_if_mux_52_cse = MUX1HOT_s_1_1_2(1'b1, and_2987_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26 = weight_mem_banks_write_if_for_if_mux_52_cse;
  assign weight_mem_banks_write_if_for_if_mux_53_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_2987_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26 = weight_mem_banks_write_if_for_if_mux_53_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26 = weight_mem_banks_write_if_for_if_mux_52_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26 = weight_mem_banks_write_if_for_if_mux_53_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_13
      = weight_mem_banks_write_if_for_if_mux_52_cse;
    assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_13
      = weight_mem_banks_write_if_for_if_mux_53_cse;
  assign weight_mem_banks_read_for_mux_52_cse = MUX1HOT_s_1_1_2(1'b1, or_1457_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27 = weight_mem_banks_read_for_mux_52_cse;
  assign weight_mem_banks_read_for_mux_53_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, or_1457_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27 = weight_mem_banks_read_for_mux_53_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27 = weight_mem_banks_read_for_mux_52_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27 = weight_mem_banks_read_for_mux_53_cse;
  assign weight_mem_banks_write_if_for_if_mux_56_cse = MUX1HOT_s_1_1_2(1'b1, and_2983_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_28 = weight_mem_banks_write_if_for_if_mux_56_cse;
  assign weight_mem_banks_write_if_for_if_mux_57_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_2983_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_28 = weight_mem_banks_write_if_for_if_mux_57_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_28 = weight_mem_banks_write_if_for_if_mux_56_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_28 = weight_mem_banks_write_if_for_if_mux_57_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_14
      = weight_mem_banks_write_if_for_if_mux_56_cse;
 assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_14
      = weight_mem_banks_write_if_for_if_mux_57_cse;
  assign weight_mem_banks_read_for_mux_56_cse = MUX1HOT_s_1_1_2(1'b1, or_1461_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_29 = weight_mem_banks_read_for_mux_56_cse;
  assign weight_mem_banks_read_for_mux_57_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, or_1461_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_29 = weight_mem_banks_read_for_mux_57_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_29 = weight_mem_banks_read_for_mux_56_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_29 = weight_mem_banks_read_for_mux_57_cse;
  assign weight_mem_banks_write_if_for_if_mux_60_cse = MUX1HOT_s_1_1_2(1'b1, and_2979_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_30 = weight_mem_banks_write_if_for_if_mux_60_cse;
  assign weight_mem_banks_write_if_for_if_mux_61_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_2979_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_30 = weight_mem_banks_write_if_for_if_mux_61_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_30 = weight_mem_banks_write_if_for_if_mux_60_cse;
 
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_30 = weight_mem_banks_write_if_for_if_mux_61_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_15
      = weight_mem_banks_write_if_for_if_mux_60_cse;
  
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_15
      = weight_mem_banks_write_if_for_if_mux_61_cse;
  assign weight_mem_banks_read_for_mux_60_cse = MUX1HOT_s_1_1_2(1'b1, or_1465_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_31 = weight_mem_banks_read_for_mux_60_cse;
  
  assign weight_mem_banks_read_for_mux_61_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, or_1465_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_31 = weight_mem_banks_read_for_mux_61_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_31 = weight_mem_banks_read_for_mux_60_cse;
  
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_31 = weight_mem_banks_read_for_mux_61_cse;
  assign input_mem_banks_write_if_for_if_mux_1_cse = MUX1HOT_s_1_1_2(1'b1, or_1183_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_32 = input_mem_banks_write_if_for_if_mux_1_cse;
  
  assign input_mem_banks_write_if_for_if_mux_2_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      or_1183_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_32 = input_mem_banks_write_if_for_if_mux_2_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_32 = input_mem_banks_write_if_for_if_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_32 = input_mem_banks_write_if_for_if_mux_2_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_16
      = input_mem_banks_write_if_for_if_mux_1_cse;
 
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_16
      = input_mem_banks_write_if_for_if_mux_2_cse;
  assign input_mem_banks_read_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_2973_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_33 = input_mem_banks_read_for_mux_cse;
  
  assign input_mem_banks_read_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_2973_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_33 = input_mem_banks_read_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_33 = input_mem_banks_read_for_mux_cse;
  
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_33 = input_mem_banks_read_for_mux_1_cse;
  assign or_1521_cse = and_5345_cse | is_start_sva;
  assign PECore_RunMac_if_and_208_cse = (~ crossbar_spec_PE_Weight_WordType_16U_16U_for_land_13_lpi_1_dfm)
      & PECore_RunMac_if_and_433_cse;
  assign PECore_RunMac_if_and_209_cse = crossbar_spec_PE_Weight_WordType_16U_16U_for_land_13_lpi_1_dfm
      & PECore_RunMac_if_and_433_cse;
  assign PECore_RunMac_if_and_176_cse = (~ crossbar_spec_PE_Weight_WordType_16U_16U_for_land_15_lpi_1_dfm)
      & PECore_RunMac_if_and_433_cse;
  assign PECore_RunMac_if_and_177_cse = crossbar_spec_PE_Weight_WordType_16U_16U_for_land_15_lpi_1_dfm
      & PECore_RunMac_if_and_433_cse;
  assign PECore_RunMac_if_and_144_cse = (~ crossbar_spec_PE_Weight_WordType_16U_16U_for_land_14_lpi_1_dfm)
      & PECore_RunMac_if_and_433_cse;
  assign PECore_RunMac_if_and_145_cse = crossbar_spec_PE_Weight_WordType_16U_16U_for_land_14_lpi_1_dfm
      & PECore_RunMac_if_and_433_cse;
  assign PECore_RunMac_if_and_112_cse = (~ crossbar_spec_PE_Weight_WordType_16U_16U_for_land_lpi_1_dfm)
      & PECore_RunMac_if_and_433_cse;
  assign PECore_RunMac_if_and_113_cse = crossbar_spec_PE_Weight_WordType_16U_16U_for_land_lpi_1_dfm
      & PECore_RunMac_if_and_433_cse;
  assign PECore_PushAxiRsp_if_and_cse = PECoreRun_wen & ((w_axi_rsp_lpi_1_dfm_1 &
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm & (~ is_start_sva)
      & (fsm_output[3])) | or_tmp_1655);
  assign PECore_PushAxiRsp_if_and_10_cse = PECoreRun_wen & (~((~ w_axi_rsp_lpi_1_dfm_1)
      | is_start_sva | (~ (fsm_output[3]))));
  assign PECore_PushAxiRsp_if_and_45_cse = (~ or_tmp_545) & PECore_PushAxiRsp_if_asn_70;
  assign and_5501_cse = PECore_PushAxiRsp_if_and_45_cse & (~ or_dcpl_717);
  assign and_5502_cse = input_mem_banks_load_store_for_else_and_cse & (~ crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm);
  assign PECore_PushAxiRsp_if_and_47_enex5 = PECore_PushAxiRsp_if_and_10_cse & reg_PECore_RunMac_if_mux_123_1_enexo;
  assign PECore_PushAxiRsp_if_and_48_enex5 = PECore_PushAxiRsp_if_and_10_cse & reg_PECore_RunMac_if_mux_142_1_enexo;
  assign PECore_PushAxiRsp_if_and_49_enex5 = PECore_PushAxiRsp_if_and_10_cse & reg_rva_out_reg_data_47_40_sva_dfm_4_enexo;
  assign PECore_PushAxiRsp_if_and_50_enex5 = PECore_PushAxiRsp_if_and_10_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_enexo;
  assign PECore_PushAxiRsp_if_and_51_enex5 = PECore_PushAxiRsp_if_and_10_cse & reg_rva_out_reg_data_63_56_sva_dfm_4_enexo;
  assign PECore_PushAxiRsp_if_and_52_enex5 = PECore_PushAxiRsp_if_and_10_cse & reg_rva_out_reg_data_71_64_sva_dfm_4_enexo;
  assign PECore_PushAxiRsp_if_and_53_enex5 = PECore_PushAxiRsp_if_and_10_cse & reg_rva_out_reg_data_79_72_sva_dfm_4_enexo;
  assign PECore_PushAxiRsp_if_and_54_enex5 = PECore_PushAxiRsp_if_and_10_cse & reg_rva_out_reg_data_87_80_sva_dfm_4_enexo;
  assign PECore_PushAxiRsp_if_and_55_enex5 = PECore_PushAxiRsp_if_and_10_cse & reg_rva_out_reg_data_95_88_sva_dfm_4_enexo;
  assign PECore_PushAxiRsp_if_and_56_enex5 = PECore_PushAxiRsp_if_and_10_cse & reg_rva_out_reg_data_103_96_sva_dfm_4_enexo;
  assign PECore_PushAxiRsp_if_and_57_enex5 = PECore_PushAxiRsp_if_and_10_cse & reg_rva_out_reg_data_111_104_sva_dfm_4_enexo;
  assign PECore_PushAxiRsp_if_and_58_enex5 = PECore_PushAxiRsp_if_and_10_cse & reg_rva_out_reg_data_119_112_sva_dfm_4_enexo;
  assign PECore_PushAxiRsp_if_and_59_enex5 = PECore_PushAxiRsp_if_and_10_cse & reg_rva_out_reg_data_127_120_sva_dfm_4_enexo;
  assign PECore_PushOutput_if_and_cse = PECoreRun_wen & (~((~ state_2_0_sva_2) |
      state_2_0_sva_1 | or_dcpl_247 | (~ (fsm_output[3]))));
  assign PECore_PushOutput_if_and_16_enex5 = PECore_PushOutput_if_and_cse & reg_act_port_reg_data_0_enexo;
  assign PECore_PushOutput_if_and_17_enex5 = PECore_PushOutput_if_and_cse & reg_act_port_reg_data_1_enexo;
  assign PECore_PushOutput_if_and_18_enex5 = PECore_PushOutput_if_and_cse & reg_act_port_reg_data_2_enexo;
  assign PECore_PushOutput_if_and_19_enex5 = PECore_PushOutput_if_and_cse & reg_act_port_reg_data_3_enexo;
  assign PECore_PushOutput_if_and_20_enex5 = PECore_PushOutput_if_and_cse & reg_act_port_reg_data_4_enexo;
  assign PECore_PushOutput_if_and_21_enex5 = PECore_PushOutput_if_and_cse & reg_act_port_reg_data_5_enexo;
  assign PECore_PushOutput_if_and_22_enex5 = PECore_PushOutput_if_and_cse & reg_act_port_reg_data_6_enexo;
  assign PECore_PushOutput_if_and_25_enex5 = PECore_PushOutput_if_and_cse & reg_act_port_reg_data_9_enexo;
  assign PECore_PushOutput_if_and_26_enex5 = PECore_PushOutput_if_and_cse & reg_act_port_reg_data_10_enexo;
  assign PECore_PushOutput_if_and_28_enex5 = PECore_PushOutput_if_and_cse & reg_act_port_reg_data_asn_3_enexo;
  assign PECore_PushOutput_if_and_29_enex5 = PECore_PushOutput_if_and_cse & reg_act_port_reg_data_asn_2_enexo;
  assign PECore_PushOutput_if_and_30_enex5 = PECore_PushOutput_if_and_cse & reg_act_port_reg_data_asn_1_enexo;
  assign PECore_PushOutput_if_and_31_enex5 = PECore_PushOutput_if_and_cse & reg_act_port_reg_data_asn_enexo;
  assign or_2419_rmff = (and_dcpl_211 & nor_499_cse) | and_2907_cse;
  assign input_mem_banks_read_read_data_and_nl = (~ or_796_cse) & (fsm_output[2]);
  assign input_mem_banks_read_read_data_mux_rmff = MUX_v_128_2_2(input_mem_banks_read_read_data_lpi_1,
      input_mem_banks_bank_array_impl_data0_rsci_q_d, input_mem_banks_read_read_data_and_nl);
  assign or_1534_cse = state_2_0_sva_0 | (~ state_2_0_sva_1) | state_2_0_sva_2;
  assign or_1536_nl = (~ while_stage_0_2) | reg_PECore_RunMac_asn_15_itm_1_ftd_2
      | reg_PECore_RunMac_asn_15_itm_1_ftd | (~ and_5335_cse);
  assign nor_244_nl = ~(and_5335_cse | and_dcpl_135);
  assign or_1531_nl = reg_PECore_RunMac_asn_15_itm_1_ftd_2 | reg_PECore_RunMac_asn_15_itm_1_ftd;
  assign mux_591_nl = MUX_s_1_2_2(nor_244_nl, or_500_cse, or_1531_nl);
  assign or_1530_nl = reg_PECore_RunMac_asn_15_itm_1_ftd_2 | reg_PECore_RunMac_asn_15_itm_1_ftd
      | (~ and_5335_cse);
  assign mux_592_nl = MUX_s_1_2_2(mux_591_nl, or_1530_nl, state_2_0_sva_0);
  assign mux_593_nl = MUX_s_1_2_2(or_1534_cse, mux_592_nl, while_stage_0_2);
  assign mux_594_nl = MUX_s_1_2_2(or_1536_nl, mux_593_nl, is_start_sva);
  assign or_2421_rmff = (and_dcpl_211 & or_dcpl_251) | and_2907_cse | ((~ mux_594_nl)
      & (fsm_output[2]));
  assign nor_242_nl = ~(state_2_0_sva_1 | input_port_PopNB_mioi_ivld_mxwt | (~ or_tmp_1286));
  assign nor_243_nl = ~(and_cse | (~ or_tmp_1286));
  assign mux_595_nl = MUX_s_1_2_2(nor_242_nl, nor_243_nl, state_2_0_sva_0);
  assign mux_596_nl = MUX_s_1_2_2(mux_595_nl, or_tmp_1286, state_2_0_sva_2);
  assign or_2422_rmff = ((~ mux_596_nl) & (fsm_output[1])) | ((input_read_req_valid_lpi_1_dfm_5
      | input_write_req_valid_lpi_1_dfm_5) & (fsm_output[2]));
  assign or_2423_rmff = (((weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]) | weight_mem_read_arbxbar_xbar_for_3_16_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp)
      & (fsm_output[1])) | (((weight_mem_write_arbxbar_xbar_for_empty_sva[15]) |
      weight_mem_read_arbxbar_xbar_for_3_16_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva)
      & (fsm_output[2]));
  assign or_2424_rmff = ((weight_mem_read_arbxbar_xbar_for_3_15_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      | (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14])) & (fsm_output[1])) |
      (((weight_mem_write_arbxbar_xbar_for_empty_sva[14]) | weight_mem_read_arbxbar_xbar_for_3_15_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva)
      & (fsm_output[2]));
  assign or_2425_rmff = ((weight_mem_read_arbxbar_xbar_for_3_14_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      | (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13])) & (fsm_output[1])) |
      (((weight_mem_write_arbxbar_xbar_for_empty_sva[13]) | weight_mem_read_arbxbar_xbar_for_3_14_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva)
      & (fsm_output[2]));
  assign or_2426_rmff = ((weight_mem_read_arbxbar_xbar_for_3_13_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      | (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12])) & (fsm_output[1])) |
      (((weight_mem_write_arbxbar_xbar_for_empty_sva[12]) | weight_mem_read_arbxbar_xbar_for_3_13_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva)
      & (fsm_output[2]));
  assign or_2427_rmff = ((weight_mem_read_arbxbar_xbar_for_3_12_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      | (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11])) & (fsm_output[1])) |
      (((weight_mem_write_arbxbar_xbar_for_empty_sva[11]) | weight_mem_read_arbxbar_xbar_for_3_12_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva)
      & (fsm_output[2]));
  assign or_2428_rmff = (((weight_mem_write_arbxbar_xbar_for_lshift_tmp[10]) | weight_mem_read_arbxbar_xbar_for_3_11_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp)
      & (fsm_output[1])) | (((weight_mem_write_arbxbar_xbar_for_empty_sva[10]) |
      weight_mem_read_arbxbar_xbar_for_3_11_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva)
      & (fsm_output[2]));
  assign or_2429_rmff = (((weight_mem_write_arbxbar_xbar_for_lshift_tmp[9]) | weight_mem_read_arbxbar_xbar_for_3_10_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp)
      & (fsm_output[1])) | (((weight_mem_write_arbxbar_xbar_for_empty_sva[9]) | weight_mem_read_arbxbar_xbar_for_3_10_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva)
      & (fsm_output[2]));
  assign or_2430_rmff = ((weight_mem_read_arbxbar_xbar_for_3_9_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      | (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8])) & (fsm_output[1])) | ((weight_mem_read_arbxbar_xbar_for_3_9_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
      | (weight_mem_write_arbxbar_xbar_for_empty_sva[8])) & (fsm_output[2]));
  assign or_2431_rmff = ((weight_mem_read_arbxbar_xbar_for_3_8_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      | (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7])) & (fsm_output[1])) | ((weight_mem_read_arbxbar_xbar_for_3_8_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
      | (weight_mem_write_arbxbar_xbar_for_empty_sva[7])) & (fsm_output[2]));
  assign or_2432_rmff = (((weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]) | weight_mem_read_arbxbar_xbar_for_3_7_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp)
      & (fsm_output[1])) | ((weight_mem_read_arbxbar_xbar_for_3_7_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
      | (weight_mem_write_arbxbar_xbar_for_empty_sva[6])) & (fsm_output[2]));
  assign or_2433_rmff = (((weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]) | weight_mem_read_arbxbar_xbar_for_3_6_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp)
      & (fsm_output[1])) | ((weight_mem_read_arbxbar_xbar_for_3_6_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
      | (weight_mem_write_arbxbar_xbar_for_empty_sva[5])) & (fsm_output[2]));
  assign or_2434_rmff = ((weight_mem_read_arbxbar_xbar_for_3_5_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      | (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4])) & (fsm_output[1])) | ((weight_mem_read_arbxbar_xbar_for_3_5_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
      | (weight_mem_write_arbxbar_xbar_for_empty_sva[4])) & (fsm_output[2]));
  assign or_2435_rmff = (((weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]) | weight_mem_read_arbxbar_xbar_for_3_4_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp)
      & (fsm_output[1])) | ((weight_mem_read_arbxbar_xbar_for_3_4_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
      | (weight_mem_write_arbxbar_xbar_for_empty_sva[3])) & (fsm_output[2]));
  assign or_2436_rmff = (((weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]) | weight_mem_read_arbxbar_xbar_for_3_3_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp)
      & (fsm_output[1])) | ((weight_mem_read_arbxbar_xbar_for_3_3_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
      | (weight_mem_write_arbxbar_xbar_for_empty_sva[2])) & (fsm_output[2]));
  assign or_2437_rmff = (((weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]) | weight_mem_read_arbxbar_xbar_for_3_2_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp)
      & (fsm_output[1])) | ((weight_mem_read_arbxbar_xbar_for_3_2_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
      | (weight_mem_write_arbxbar_xbar_for_empty_sva[1])) & (fsm_output[2]));
  assign or_2438_rmff = (((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]) | weight_mem_read_arbxbar_xbar_for_3_1_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp)
      & (fsm_output[1])) | ((weight_mem_read_arbxbar_xbar_for_3_1_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
      | (weight_mem_write_arbxbar_xbar_for_empty_sva[0])) & (fsm_output[2]));
  assign and_2966_cse = (~ is_start_sva) & (fsm_output[3]);
  assign nor_241_nl = ~((rva_in_PopNB_mioi_idat_mxwt[168]) | input_port_PopNB_mioi_ivld_mxwt
      | is_start_sva | (rva_in_PopNB_mioi_idat_mxwt[151:148]!=4'b0110) | (~ rva_in_PopNB_mioi_ivld_mxwt));
  assign mux_598_nl = MUX_s_1_2_2(nor_241_nl, or_tmp_20, state_2_0_sva_1);
  assign mux_597_nl = MUX_s_1_2_2((~ or_tmp_18), or_tmp_20, and_cse);
  assign mux_599_nl = MUX_s_1_2_2(mux_598_nl, mux_597_nl, state_2_0_sva_0);
  assign mux_600_nl = MUX_s_1_2_2(mux_599_nl, (~ or_tmp_18), state_2_0_sva_2);
  assign and_2973_cse = mux_600_nl & (fsm_output[1]);
  assign or_1584_cse = (~ (rva_in_PopNB_mioi_idat_mxwt[168])) | (rva_in_PopNB_mioi_idat_mxwt[148])
      | (~ (rva_in_PopNB_mioi_idat_mxwt[149])) | (rva_in_PopNB_mioi_idat_mxwt[151])
      | nand_199_cse;
  assign weight_write_data_data_mux1h_rmff = (rva_in_PopNB_mioi_idat_mxwt[7:0]) &
      ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
      & (signext_8_1(rva_in_PopNB_mioi_idat_mxwt[168])) & ({{7{rva_in_PopNB_mioi_ivld_mxwt}},
      rva_in_PopNB_mioi_ivld_mxwt}) & (signext_8_1(~ is_start_sva));
  assign weight_write_data_data_mux1h_1_rmff = (rva_in_PopNB_mioi_idat_mxwt[15:8])
      & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
      & (signext_8_1(rva_in_PopNB_mioi_idat_mxwt[168])) & ({{7{rva_in_PopNB_mioi_ivld_mxwt}},
      rva_in_PopNB_mioi_ivld_mxwt}) & (signext_8_1(~ is_start_sva));
  assign weight_write_data_data_mux1h_2_rmff = (rva_in_PopNB_mioi_idat_mxwt[23:16])
      & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
      & (signext_8_1(rva_in_PopNB_mioi_idat_mxwt[168])) & ({{7{rva_in_PopNB_mioi_ivld_mxwt}},
      rva_in_PopNB_mioi_ivld_mxwt}) & (signext_8_1(~ is_start_sva));
  assign weight_write_data_data_mux1h_3_rmff = (rva_in_PopNB_mioi_idat_mxwt[31:24])
      & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
      & (signext_8_1(rva_in_PopNB_mioi_idat_mxwt[168])) & ({{7{rva_in_PopNB_mioi_ivld_mxwt}},
      rva_in_PopNB_mioi_ivld_mxwt}) & (signext_8_1(~ is_start_sva));
  assign weight_write_data_data_mux1h_4_rmff = (rva_in_PopNB_mioi_idat_mxwt[39:32])
      & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
      & (signext_8_1(rva_in_PopNB_mioi_idat_mxwt[168])) & ({{7{rva_in_PopNB_mioi_ivld_mxwt}},
      rva_in_PopNB_mioi_ivld_mxwt}) & (signext_8_1(~ is_start_sva));
  assign weight_write_data_data_mux1h_5_rmff = (rva_in_PopNB_mioi_idat_mxwt[47:40])
      & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
      & (signext_8_1(rva_in_PopNB_mioi_idat_mxwt[168])) & ({{7{rva_in_PopNB_mioi_ivld_mxwt}},
      rva_in_PopNB_mioi_ivld_mxwt}) & (signext_8_1(~ is_start_sva));
  assign weight_write_data_data_mux1h_6_rmff = (rva_in_PopNB_mioi_idat_mxwt[55:48])
      & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
      & (signext_8_1(rva_in_PopNB_mioi_idat_mxwt[168])) & ({{7{rva_in_PopNB_mioi_ivld_mxwt}},
      rva_in_PopNB_mioi_ivld_mxwt}) & (signext_8_1(~ is_start_sva));
  assign weight_write_data_data_mux1h_7_rmff = (rva_in_PopNB_mioi_idat_mxwt[63:56])
      & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
      & (signext_8_1(rva_in_PopNB_mioi_idat_mxwt[168])) & ({{7{rva_in_PopNB_mioi_ivld_mxwt}},
      rva_in_PopNB_mioi_ivld_mxwt}) & (signext_8_1(~ is_start_sva));
  assign weight_write_data_data_mux1h_8_rmff = (rva_in_PopNB_mioi_idat_mxwt[71:64])
      & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
      & (signext_8_1(rva_in_PopNB_mioi_idat_mxwt[168])) & ({{7{rva_in_PopNB_mioi_ivld_mxwt}},
      rva_in_PopNB_mioi_ivld_mxwt}) & (signext_8_1(~ is_start_sva));
  assign weight_write_data_data_mux1h_9_rmff = (rva_in_PopNB_mioi_idat_mxwt[79:72])
      & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
      & (signext_8_1(rva_in_PopNB_mioi_idat_mxwt[168])) & ({{7{rva_in_PopNB_mioi_ivld_mxwt}},
      rva_in_PopNB_mioi_ivld_mxwt}) & (signext_8_1(~ is_start_sva));
  assign weight_write_data_data_mux1h_10_rmff = (rva_in_PopNB_mioi_idat_mxwt[87:80])
      & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
      & (signext_8_1(rva_in_PopNB_mioi_idat_mxwt[168])) & ({{7{rva_in_PopNB_mioi_ivld_mxwt}},
      rva_in_PopNB_mioi_ivld_mxwt}) & (signext_8_1(~ is_start_sva));
  assign weight_write_data_data_mux1h_11_rmff = (rva_in_PopNB_mioi_idat_mxwt[95:88])
      & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
      & (signext_8_1(rva_in_PopNB_mioi_idat_mxwt[168])) & ({{7{rva_in_PopNB_mioi_ivld_mxwt}},
      rva_in_PopNB_mioi_ivld_mxwt}) & (signext_8_1(~ is_start_sva));
  assign weight_write_data_data_mux1h_12_rmff = (rva_in_PopNB_mioi_idat_mxwt[103:96])
      & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
      & (signext_8_1(rva_in_PopNB_mioi_idat_mxwt[168])) & ({{7{rva_in_PopNB_mioi_ivld_mxwt}},
      rva_in_PopNB_mioi_ivld_mxwt}) & (signext_8_1(~ is_start_sva));
  assign weight_write_data_data_mux1h_13_rmff = (rva_in_PopNB_mioi_idat_mxwt[111:104])
      & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
      & (signext_8_1(rva_in_PopNB_mioi_idat_mxwt[168])) & ({{7{rva_in_PopNB_mioi_ivld_mxwt}},
      rva_in_PopNB_mioi_ivld_mxwt}) & (signext_8_1(~ is_start_sva));
  assign weight_write_data_data_mux1h_14_rmff = (rva_in_PopNB_mioi_idat_mxwt[119:112])
      & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
      & (signext_8_1(rva_in_PopNB_mioi_idat_mxwt[168])) & ({{7{rva_in_PopNB_mioi_ivld_mxwt}},
      rva_in_PopNB_mioi_ivld_mxwt}) & (signext_8_1(~ is_start_sva));
  assign while_while_and_18_itm = (rva_in_PopNB_mioi_idat_mxwt[127:120]) & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}},
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}) & (signext_8_1(rva_in_PopNB_mioi_idat_mxwt[168]))
      & ({{7{rva_in_PopNB_mioi_ivld_mxwt}}, rva_in_PopNB_mioi_ivld_mxwt}) & (signext_8_1(~
      is_start_sva));
  assign is_start_and_cse = PECoreRun_wen & (fsm_output[4]);
  assign PECore_UpdateFSM_switch_lp_not_47_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_1;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_4_cse
      = MUX_v_32_2_2(32'b00000000000000000000000000000000, z_out_25, PECore_UpdateFSM_switch_lp_not_47_nl);
  assign accum_vector_data_and_6_cse = PECoreRun_wen & (~(or_dcpl_718 | nor_499_cse));
  assign PECore_UpdateFSM_switch_lp_not_48_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_1;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_3_cse
      = MUX_v_32_2_2(32'b00000000000000000000000000000000, z_out_26, PECore_UpdateFSM_switch_lp_not_48_nl);
  assign PECore_UpdateFSM_switch_lp_not_49_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_1;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_2_cse
      = MUX_v_32_2_2(32'b00000000000000000000000000000000, z_out_27, PECore_UpdateFSM_switch_lp_not_49_nl);
  assign while_and_77_m1c = (~(z_out_24_32 | PECore_RunBias_if_for_11_operator_32_true_slc_operator_32_true_acc_13_svs_mx0))
      & while_and_46_tmp_1;
  assign while_and_221_nl = and_dcpl_437 & while_and_77_m1c;
  assign while_while_mux_9_m1c = MUX_s_1_2_2(while_and_221_nl, (~ while_and_46_tmp_1),
      or_dcpl_251);
  assign while_and_225_nl = or_dcpl_295 & while_and_77_m1c;
  assign while_and_226_nl = pe_config_is_bias_sva & while_and_61_m1c;
  assign while_and_227_nl = pe_config_is_bias_sva & while_and_79_m1c;
  assign while_mux1h_47_m1c = MUX1HOT_s_1_3_2(while_and_225_nl, while_and_226_nl,
      while_and_227_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign while_or_11_nl = ((fsm_output[1]) & while_while_mux_9_m1c) | (or_dcpl_251
      & while_mux1h_47_m1c);
  assign while_and_288_nl = (fsm_output[4]) & while_while_mux_9_m1c;
  assign while_and_289_nl = (fsm_output[3]) & while_while_mux_9_m1c;
  assign while_and_222_nl = and_dcpl_439 & while_and_77_m1c;
  assign while_and_223_nl = (~ pe_config_is_bias_sva) & while_and_61_m1c;
  assign while_and_224_nl = (~ pe_config_is_bias_sva) & while_and_79_m1c;
  assign while_mux1h_46_nl = MUX1HOT_s_1_3_2(while_and_222_nl, while_and_223_nl,
      while_and_224_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign while_and_290_nl = (~ or_dcpl_251) & while_mux1h_47_m1c;
  assign PECore_RunBias_if_for_and_55_nl = z_out_24_32 & (~ PECore_RunBias_if_for_11_operator_32_true_slc_operator_32_true_acc_13_svs_mx0)
      & while_and_46_tmp_1;
  assign PECore_RunBias_if_for_and_56_nl = z_out_22_32 & (~ z_out_11_13) & while_and_46_tmp_1;
  assign PECore_RunBias_if_for_and_57_nl = z_out_24_32 & (~ PECore_RunBias_if_for_12_operator_32_true_slc_operator_32_true_acc_13_svs_mx2)
      & while_and_46_tmp_1;
  assign while_mux1h_48_nl = MUX1HOT_s_1_3_2(PECore_RunBias_if_for_and_55_nl, PECore_RunBias_if_for_and_56_nl,
      PECore_RunBias_if_for_and_57_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign while_and_228_nl = PECore_RunBias_if_for_11_operator_32_true_slc_operator_32_true_acc_13_svs_mx0
      & while_and_46_tmp_1;
  assign while_and_229_nl = z_out_11_13 & while_and_46_tmp_1;
  assign while_and_230_nl = PECore_RunBias_if_for_12_operator_32_true_slc_operator_32_true_acc_13_svs_mx2
      & while_and_46_tmp_1;
  assign while_mux1h_49_nl = MUX1HOT_s_1_3_2(while_and_228_nl, while_and_229_nl,
      while_and_230_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign mux1h_12_nl = MUX1HOT_v_20_7_2((z_out_30[19:0]), act_port_reg_data_2_sva,
      act_port_reg_data_11_sva, (PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_11_sva[19:0]),
      reg_PECore_RunBias_if_accum_vector_out_data_11_lpi_1_dfm_ftd_12, 20'b10000000000000000001,
      20'b01111111111111111111, {while_or_11_nl , while_and_288_nl , while_and_289_nl
      , while_mux1h_46_nl , while_and_290_nl , while_mux1h_48_nl , while_mux1h_49_nl});
  assign PECore_UpdateFSM_switch_lp_not_65_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_1;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_26_cse
      = MUX_v_20_2_2(20'b00000000000000000000, mux1h_12_nl, PECore_UpdateFSM_switch_lp_not_65_nl);
  assign act_port_reg_data_and_8_cse = PECoreRun_wen & (~((~((PECore_UpdateFSM_switch_lp_equal_tmp_1
      | while_and_46_tmp_1) & while_stage_0_2)) | nor_499_cse));
  assign while_and_75_m1c = (~(z_out_23_32 | PECore_RunBias_if_for_10_operator_32_true_slc_operator_32_true_acc_13_svs_mx0))
      & while_and_46_tmp_1;
  assign while_and_231_nl = and_dcpl_437 & while_and_75_m1c;
  assign while_while_mux_11_m1c = MUX_s_1_2_2(while_and_231_nl, (~ while_and_46_tmp_1),
      or_dcpl_251);
  assign while_and_235_nl = or_dcpl_295 & while_and_75_m1c;
  assign while_and_236_nl = pe_config_is_bias_sva & while_and_57_m1c;
  assign while_and_237_nl = pe_config_is_bias_sva & while_and_59_m1c;
  assign while_mux1h_52_m1c = MUX1HOT_s_1_3_2(while_and_235_nl, while_and_236_nl,
      while_and_237_nl, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])});
  assign while_or_10_nl = ((fsm_output[1]) & while_while_mux_11_m1c) | (or_dcpl_251
      & while_mux1h_52_m1c);
  assign while_and_283_nl = (fsm_output[3]) & while_while_mux_11_m1c;
  assign while_and_284_nl = (fsm_output[4]) & while_while_mux_11_m1c;
  assign while_and_232_nl = and_dcpl_439 & while_and_75_m1c;
  assign while_and_233_nl = (~ pe_config_is_bias_sva) & while_and_57_m1c;
  assign while_and_234_nl = (~ pe_config_is_bias_sva) & while_and_59_m1c;
  assign while_mux1h_51_nl = MUX1HOT_s_1_3_2(while_and_232_nl, while_and_233_nl,
      while_and_234_nl, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])});
  assign while_and_285_nl = (~ or_dcpl_251) & while_mux1h_52_m1c;
  assign PECore_RunBias_if_for_and_58_nl = z_out_23_32 & (~ PECore_RunBias_if_for_10_operator_32_true_slc_operator_32_true_acc_13_svs_mx0)
      & while_and_46_tmp_1;
  assign PECore_RunBias_if_for_and_59_nl = z_out_21_32 & (~ PECore_RunBias_if_for_1_operator_32_true_slc_operator_32_true_acc_13_svs_mx2)
      & while_and_46_tmp_1;
  assign PECore_RunBias_if_for_and_60_nl = z_out_23_32 & (~ PECore_RunBias_if_for_2_operator_32_true_slc_operator_32_true_acc_13_svs_mx2)
      & while_and_46_tmp_1;
  assign while_mux1h_53_nl = MUX1HOT_s_1_3_2(PECore_RunBias_if_for_and_58_nl, PECore_RunBias_if_for_and_59_nl,
      PECore_RunBias_if_for_and_60_nl, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])});
  assign while_and_238_nl = PECore_RunBias_if_for_10_operator_32_true_slc_operator_32_true_acc_13_svs_mx0
      & while_and_46_tmp_1;
  assign while_and_239_nl = PECore_RunBias_if_for_1_operator_32_true_slc_operator_32_true_acc_13_svs_mx2
      & while_and_46_tmp_1;
  assign while_and_240_nl = PECore_RunBias_if_for_2_operator_32_true_slc_operator_32_true_acc_13_svs_mx2
      & while_and_46_tmp_1;
  assign while_mux1h_54_nl = MUX1HOT_s_1_3_2(while_and_238_nl, while_and_239_nl,
      while_and_240_nl, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])});
  assign mux1h_13_nl = MUX1HOT_v_20_7_2((z_out_29[19:0]), act_port_reg_data_0_sva,
      act_port_reg_data_1_sva, (PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_1_sva[19:0]),
      reg_PECore_RunBias_if_accum_vector_out_data_10_lpi_1_dfm_ftd_12, 20'b10000000000000000001,
      20'b01111111111111111111, {while_or_10_nl , while_and_283_nl , while_and_284_nl
      , while_mux1h_51_nl , while_and_285_nl , while_mux1h_53_nl , while_mux1h_54_nl});
  assign PECore_UpdateFSM_switch_lp_not_66_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_1;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_25_cse
      = MUX_v_20_2_2(20'b00000000000000000000, mux1h_13_nl, PECore_UpdateFSM_switch_lp_not_66_nl);
  assign while_and_69_m1c = (~(z_out_22_32 | PECore_RunBias_if_for_7_operator_32_true_slc_operator_32_true_acc_13_svs_mx0))
      & while_and_46_tmp_1;
  assign while_and_241_nl = and_dcpl_437 & while_and_69_m1c;
  assign while_while_mux_13_m1c = MUX_s_1_2_2(while_and_241_nl, (~ while_and_46_tmp_1),
      or_dcpl_251);
  assign while_and_245_nl = or_dcpl_295 & while_and_69_m1c;
  assign while_and_246_nl = pe_config_is_bias_sva & while_and_65_m1c;
  assign while_and_247_nl = pe_config_is_bias_sva & while_and_73_m1c;
  assign while_mux1h_57_m1c = MUX1HOT_s_1_3_2(while_and_245_nl, while_and_246_nl,
      while_and_247_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign while_or_9_nl = ((fsm_output[1]) & while_while_mux_13_m1c) | (or_dcpl_251
      & while_mux1h_57_m1c);
  assign while_and_278_nl = (fsm_output[4]) & while_while_mux_13_m1c;
  assign while_and_279_nl = (fsm_output[3]) & while_while_mux_13_m1c;
  assign while_and_242_nl = and_dcpl_439 & while_and_69_m1c;
  assign while_and_243_nl = (~ pe_config_is_bias_sva) & while_and_65_m1c;
  assign while_and_244_nl = (~ pe_config_is_bias_sva) & while_and_73_m1c;
  assign while_mux1h_56_nl = MUX1HOT_s_1_3_2(while_and_242_nl, while_and_243_nl,
      while_and_244_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign while_and_280_nl = (~ or_dcpl_251) & while_mux1h_57_m1c;
  assign PECore_RunBias_if_for_and_61_nl = z_out_22_32 & (~ PECore_RunBias_if_for_7_operator_32_true_slc_operator_32_true_acc_13_svs_mx0)
      & while_and_46_tmp_1;
  assign PECore_RunBias_if_for_and_62_nl = z_out_24_32 & (~ z_out_13_13) & while_and_46_tmp_1;
  assign PECore_RunBias_if_for_and_63_nl = z_out_22_32 & (~ z_out_12_13) & while_and_46_tmp_1;
  assign while_mux1h_58_nl = MUX1HOT_s_1_3_2(PECore_RunBias_if_for_and_61_nl, PECore_RunBias_if_for_and_62_nl,
      PECore_RunBias_if_for_and_63_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign while_and_248_nl = PECore_RunBias_if_for_7_operator_32_true_slc_operator_32_true_acc_13_svs_mx0
      & while_and_46_tmp_1;
  assign while_mux1h_59_nl = MUX1HOT_s_1_3_2(while_and_248_nl, while_and_66_cse,
      while_and_74_cse, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign mux1h_14_nl = MUX1HOT_v_20_7_2((z_out_32[19:0]), act_port_reg_data_4_sva,
      act_port_reg_data_8_sva, (PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_5_sva[19:0]),
      reg_PECore_RunBias_if_accum_vector_out_data_7_lpi_1_dfm_ftd_12, 20'b10000000000000000001,
      20'b01111111111111111111, {while_or_9_nl , while_and_278_nl , while_and_279_nl
      , while_mux1h_56_nl , while_and_280_nl , while_mux1h_58_nl , while_mux1h_59_nl});
  assign PECore_UpdateFSM_switch_lp_not_67_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_1;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_22_cse
      = MUX_v_20_2_2(20'b00000000000000000000, mux1h_14_nl, PECore_UpdateFSM_switch_lp_not_67_nl);
  assign while_and_67_m1c = (~(z_out_21_32 | PECore_RunBias_if_for_6_operator_32_true_slc_operator_32_true_acc_13_svs_mx0))
      & while_and_46_tmp_1;
  assign while_and_249_nl = and_dcpl_437 & while_and_67_m1c;
  assign while_while_mux_15_m1c = MUX_s_1_2_2(while_and_249_nl, (~ while_and_46_tmp_1),
      or_dcpl_251);
  assign while_and_253_nl = or_dcpl_295 & while_and_67_m1c;
  assign while_and_254_nl = pe_config_is_bias_sva & while_and_63_m1c;
  assign while_and_255_nl = pe_config_is_bias_sva & while_and_71_m1c;
  assign while_mux1h_62_m1c = MUX1HOT_s_1_3_2(while_and_253_nl, while_and_254_nl,
      while_and_255_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign while_or_nl = ((fsm_output[1]) & while_while_mux_15_m1c) | (or_dcpl_251
      & while_mux1h_62_m1c);
  assign while_and_273_nl = (fsm_output[4]) & while_while_mux_15_m1c;
  assign while_and_274_nl = (fsm_output[3]) & while_while_mux_15_m1c;
  assign while_and_250_nl = and_dcpl_439 & while_and_67_m1c;
  assign while_and_251_nl = (~ pe_config_is_bias_sva) & while_and_63_m1c;
  assign while_and_252_nl = (~ pe_config_is_bias_sva) & while_and_71_m1c;
  assign while_mux1h_61_nl = MUX1HOT_s_1_3_2(while_and_250_nl, while_and_251_nl,
      while_and_252_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign while_and_275_nl = (~ or_dcpl_251) & while_mux1h_62_m1c;
  assign PECore_RunBias_if_for_and_64_nl = z_out_21_32 & (~ PECore_RunBias_if_for_6_operator_32_true_slc_operator_32_true_acc_13_svs_mx0)
      & while_and_46_tmp_1;
  assign PECore_RunBias_if_for_and_65_nl = z_out_21_32 & (~ z_out_12_13) & while_and_46_tmp_1;
  assign PECore_RunBias_if_for_and_66_nl = z_out_23_32 & (~ z_out_13_13) & while_and_46_tmp_1;
  assign while_mux1h_63_nl = MUX1HOT_s_1_3_2(PECore_RunBias_if_for_and_64_nl, PECore_RunBias_if_for_and_65_nl,
      PECore_RunBias_if_for_and_66_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign while_and_256_nl = PECore_RunBias_if_for_6_operator_32_true_slc_operator_32_true_acc_13_svs_mx0
      & while_and_46_tmp_1;
  assign while_mux1h_64_nl = MUX1HOT_s_1_3_2(while_and_256_nl, while_and_74_cse,
      while_and_66_cse, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign mux1h_15_nl = MUX1HOT_v_20_7_2((z_out_31[19:0]), act_port_reg_data_3_sva,
      act_port_reg_data_7_sva, (PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_4_sva[19:0]),
      reg_PECore_RunBias_if_accum_vector_out_data_6_lpi_1_dfm_ftd_12, 20'b10000000000000000001,
      20'b01111111111111111111, {while_or_nl , while_and_273_nl , while_and_274_nl
      , while_mux1h_61_nl , while_and_275_nl , while_mux1h_63_nl , while_mux1h_64_nl});
  assign PECore_UpdateFSM_switch_lp_not_38_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_1;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_21_cse
      = MUX_v_20_2_2(20'b00000000000000000000, mux1h_15_nl, PECore_UpdateFSM_switch_lp_not_38_nl);
  assign and_cse = pe_config_is_bias_sva & state_2_0_sva_1;
  assign nor_499_cse = ~((fsm_output[1:0]!=2'b00));
  assign while_and_cse = PECoreRun_wen & (~ or_dcpl_251);
  assign pe_manager_adplfloat_bias_weight_and_cse = PECoreRun_wen & (~((~ (fsm_output[1]))
      | or_dcpl_306));
  assign pe_manager_adplfloat_bias_weight_and_1_cse = PECoreRun_wen & (~((~ (fsm_output[1]))
      | or_dcpl_310));
  assign pe_manager_cluster_lut_data_and_cse = PECoreRun_wen & (~((~ (fsm_output[1]))
      | (~ PECore_DecodeAxiWrite_case_4_switch_lp_nor_13_tmp) | (~ (rva_in_PopNB_mioi_idat_mxwt[133]))
      | (~ rva_in_PopNB_mioi_ivld_mxwt) | or_dcpl_302 | or_dcpl_313));
  assign pe_manager_cluster_lut_data_and_1_cse = PECoreRun_wen & (~((~ (fsm_output[1]))
      | (~ (rva_in_PopNB_mioi_idat_mxwt[134])) | (~ PECore_DecodeAxiWrite_case_4_switch_lp_nor_9_tmp)
      | (~ rva_in_PopNB_mioi_ivld_mxwt) | or_dcpl_302 | or_dcpl_313));
  assign pe_config_manager_counter_and_cse = PECoreRun_wen & (fsm_output[1]);
  assign and_5844_cse = state_2_0_sva_2 & (~ state_2_0_sva_1) & (~ state_2_0_sva_0);
  assign weight_port_read_out_data_and_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_16U_16U_for_land_lpi_1_dfm
      & (fsm_output[2]);
  assign weight_port_read_out_data_and_16_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_16U_16U_for_land_15_lpi_1_dfm
      & (fsm_output[2]);
  assign weight_port_read_out_data_and_32_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_16U_16U_for_land_14_lpi_1_dfm
      & (fsm_output[2]);
  assign weight_port_read_out_data_and_48_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_16U_16U_for_land_13_lpi_1_dfm
      & (fsm_output[2]);
  assign weight_port_read_out_data_and_64_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm
      & (fsm_output[2]);
  assign weight_port_read_out_data_and_80_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_16U_16U_for_land_9_lpi_1_dfm
      & (fsm_output[2]);
  assign weight_port_read_out_data_and_96_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm
      & (fsm_output[2]);
  assign weight_port_read_out_data_and_112_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm
      & (fsm_output[2]);
  assign weight_port_read_out_data_and_128_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm
      & (fsm_output[2]);
  assign weight_port_read_out_data_and_136_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm
      & (fsm_output[2]);
  assign weight_port_read_out_data_and_152_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm
      & (fsm_output[2]);
  assign weight_port_read_out_data_and_168_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm
      & (fsm_output[2]);
  assign weight_port_read_out_data_and_184_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm
      & (fsm_output[2]);
  assign weight_port_read_out_data_and_200_cse = PECoreRun_wen & rva_out_reg_data_and_2_cse;
  assign while_while_nor_cse = ~((fsm_output[4]) | while_mux_440_cse);
  assign while_and_268_cse = (fsm_output[4]) & (~ while_mux_440_cse);
  assign while_and_269_nl = (~ (fsm_output[4])) & while_mux_440_cse;
  assign while_and_270_nl = (fsm_output[4]) & while_mux_440_cse;
  assign while_mux1h_67_nl = MUX1HOT_v_32_4_2(accum_vector_data_15_sva, accum_vector_data_8_sva,
      z_out_28, z_out_26, {while_while_nor_cse , while_and_268_cse , while_and_269_nl
      , while_and_270_nl});
  assign PECore_UpdateFSM_switch_lp_not_55_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_1;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_15_cse
      = MUX_v_32_2_2(32'b00000000000000000000000000000000, while_mux1h_67_nl, PECore_UpdateFSM_switch_lp_not_55_nl);
  assign accum_vector_data_and_9_cse = PECoreRun_wen & (fsm_output[3]);
  assign while_mux_nl = MUX_v_32_4_2(accum_vector_data_14_sva, accum_vector_data_7_sva,
      z_out_26, z_out_27, {while_mux_440_cse , (fsm_output[4])});
  assign PECore_UpdateFSM_switch_lp_not_56_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_1;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_14_cse
      = MUX_v_32_2_2(32'b00000000000000000000000000000000, while_mux_nl, PECore_UpdateFSM_switch_lp_not_56_nl);
  assign while_mux1h_65_nl = MUX1HOT_v_32_3_2(accum_vector_data_13_sva, PECore_RunBias_if_accum_vector_out_data_lpi_1_dfm,
      z_out_25, {while_while_nor_cse , while_and_268_cse , while_mux_440_cse});
  assign PECore_UpdateFSM_switch_lp_not_57_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_1;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_13_cse
      = MUX_v_32_2_2(32'b00000000000000000000000000000000, while_mux1h_65_nl, PECore_UpdateFSM_switch_lp_not_57_nl);
  assign while_mux_449_nl = MUX_v_32_4_2(accum_vector_data_12_sva, PECore_RunBias_if_accum_vector_out_data_13_lpi_1_dfm,
      z_out_27, z_out_28, {while_mux_440_cse , (fsm_output[4])});
  assign PECore_UpdateFSM_switch_lp_not_58_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_1;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_12_cse
      = MUX_v_32_2_2(32'b00000000000000000000000000000000, while_mux_449_nl, PECore_UpdateFSM_switch_lp_not_58_nl);
  assign while_and_81_m1c = (~(z_out_21_32 | PECore_RunBias_if_for_13_operator_32_true_slc_operator_32_true_acc_13_svs_mx1))
      & while_and_48_tmp_1;
  assign and_5871_cse = (~(state_2_0_sva_1 | state_2_0_sva_2)) & state_2_0_sva_0;
  assign and_5872_cse = (and_5871_cse | while_and_48_tmp_1) & (fsm_output[2]) & PECoreRun_wen;
  assign while_and_83_m1c = (~(z_out_24_32 | PECore_RunBias_if_for_14_operator_32_true_slc_operator_32_true_acc_13_svs_mx1))
      & while_and_48_tmp_1;
  assign while_and_85_m1c = (~(z_out_23_32 | PECore_RunBias_if_for_15_operator_32_true_slc_operator_32_true_acc_13_svs_mx1))
      & while_and_48_tmp_1;
  assign while_and_87_m1c = (~(z_out_22_32 | PECore_RunBias_if_for_16_operator_32_true_slc_operator_32_true_acc_13_svs_mx1))
      & while_and_48_tmp_1;
  assign while_and_57_m1c = (~(z_out_21_32 | PECore_RunBias_if_for_1_operator_32_true_slc_operator_32_true_acc_13_svs_mx2))
      & while_and_46_tmp_1;
  assign while_and_59_m1c = (~(z_out_23_32 | PECore_RunBias_if_for_2_operator_32_true_slc_operator_32_true_acc_13_svs_mx2))
      & while_and_46_tmp_1;
  assign while_and_61_m1c = (~(z_out_22_32 | z_out_11_13)) & while_and_46_tmp_1;
  assign while_and_63_m1c = (~(z_out_21_32 | z_out_12_13)) & while_and_46_tmp_1;
  assign while_and_79_m1c = (~(z_out_24_32 | PECore_RunBias_if_for_12_operator_32_true_slc_operator_32_true_acc_13_svs_mx2))
      & while_and_46_tmp_1;
  assign while_and_65_m1c = (~(z_out_24_32 | z_out_13_13)) & while_and_46_tmp_1;
  assign while_and_73_m1c = (~(z_out_22_32 | z_out_12_13)) & while_and_46_tmp_1;
  assign while_and_71_m1c = (~(z_out_23_32 | z_out_13_13)) & while_and_46_tmp_1;
  assign PECore_DecodeAxi_if_and_3_cse = PECoreRun_wen & (~(is_start_sva | nor_499_cse));
  assign pe_config_is_valid_and_cse = PECoreRun_wen & (~(PECore_DecodeAxiWrite_case_4_switch_lp_or_6_cse_1
      | (~ PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_31)))
      & (rva_in_PopNB_mio_mrgout_dat_sva_1[168]) & rva_in_PopNB_mioi_ivld_mxwt &
      (~ or_tmp_2232);
  assign pe_config_num_output_and_cse = PECoreRun_wen & (~((~ (fsm_output[1])) |
      or_dcpl_334));
  assign and_4031_m1c = or_1534_cse & (fsm_output[1]);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_ssc
      = PECoreRun_wen & (fsm_output[1]) & weight_mem_read_arbxbar_xbar_for_3_1_operator_31_false_operator_31_false_operator_31_false_or_seb;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_1_ssc
      = PECoreRun_wen & (fsm_output[1]) & weight_mem_read_arbxbar_xbar_for_3_2_operator_31_false_operator_31_false_operator_31_false_or_seb;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_2_ssc
      = PECoreRun_wen & (fsm_output[1]) & weight_mem_read_arbxbar_xbar_for_3_3_operator_31_false_operator_31_false_operator_31_false_or_seb;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_3_ssc
      = PECoreRun_wen & (fsm_output[1]) & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_3_tmp;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_4_ssc
      = PECoreRun_wen & (fsm_output[1]) & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_4_tmp;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_5_ssc
      = PECoreRun_wen & (fsm_output[1]) & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_5_tmp;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_6_ssc
      = PECoreRun_wen & (fsm_output[1]) & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_6_tmp;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_7_ssc
      = PECoreRun_wen & (fsm_output[1]) & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_7_tmp;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_8_ssc
      = PECoreRun_wen & (fsm_output[1]) & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_8_tmp;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_9_ssc
      = PECoreRun_wen & (fsm_output[1]) & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_9_tmp;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_10_ssc
      = PECoreRun_wen & (fsm_output[1]) & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_10_tmp;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_11_ssc
      = PECoreRun_wen & (fsm_output[1]) & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_11_tmp;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_12_ssc
      = PECoreRun_wen & (fsm_output[1]) & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_12_tmp;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_13_ssc
      = PECoreRun_wen & (fsm_output[1]) & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_13_tmp;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_14_ssc
      = PECoreRun_wen & (fsm_output[1]) & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_14_tmp;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_15_cse
      = PECoreRun_wen & (fsm_output[1]) & weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse;
  assign PECore_DecodeAxiRead_switch_lp_and_2_cse = is_start_sva & (fsm_output[4]);
  assign PECore_DecodeAxiRead_switch_lp_and_3_rgt = (~ is_start_sva) & (fsm_output[4]);
  assign PECore_CheckStart_start_reg_and_cse = PECoreRun_wen & (~(and_4616_cse |
      PECore_RunBias_if_for_and_34_rgt | PECore_DecodeAxiRead_switch_lp_and_2_cse));
  assign operator_4_false_and_cse = PECoreRun_wen & is_start_sva & (fsm_output[2]);
  assign and_5345_cse = start_PopNB_mioi_idat_mxwt & start_PopNB_mioi_ivld_mxwt &
      pe_config_is_valid_sva;
  assign operator_32_true_and_6_rgt = (~ or_dcpl_364) & (fsm_output[2]);
  assign adpfloat_tmp_is_zero_aelse_and_cse = PECoreRun_wen & (~((or_dcpl_364 & (fsm_output[2]))
      | or_tmp_2557));
  assign PECore_RunBias_if_for_and_50_rgt = is_start_sva & PECore_RunBias_if_for_or_m1c_5;
  assign PECore_RunBias_if_for_and_47_cse = (~ is_start_sva) & or_3399_cse;
  assign PECore_RunBias_if_for_and_48_cse = (~ is_start_sva) & PECore_RunBias_if_for_or_m1c_5;
  assign operator_32_true_and_12_cse = PECoreRun_wen & (~ or_dcpl_365) & (fsm_output[2]);
  assign weight_port_read_out_data_and_216_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_16U_16U_for_land_11_lpi_1_dfm
      & (fsm_output[2]);
  assign weight_port_read_out_data_and_232_cse = PECoreRun_wen & while_and_46_tmp_1
      & (fsm_output[2]);
  assign operator_32_true_and_2_rgt = (~ or_dcpl_369) & (fsm_output[2]);
  assign adpfloat_tmp_is_zero_aelse_and_4_cse = PECoreRun_wen & (~((or_dcpl_369 &
      (fsm_output[2])) | or_tmp_2557));
  assign accum_vector_data_and_15_cse = PECoreRun_wen & (PECore_UpdateFSM_switch_lp_equal_tmp_1
      | while_and_29_itm_1) & while_stage_0_2 & (fsm_output[2]);
  assign adpfloat_tmp_is_zero_aelse_and_6_cse = PECoreRun_wen & pe_config_is_bias_sva
      & is_start_sva & (fsm_output[2]);
  assign PECore_UpdateFSM_switch_lp_not_50_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_1;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_1_cse
      = MUX_v_32_2_2(32'b00000000000000000000000000000000, z_out_28, PECore_UpdateFSM_switch_lp_not_50_nl);
  assign or_500_cse = (~ state_2_0_sva_1) | state_2_0_sva_2;
  assign PECore_RunMac_if_nand_56_rgt = ~((fsm_output[2]) & is_start_sva);
  assign PECore_RunMac_if_and_674_rgt = and_dcpl_704 & (fsm_output[2]);
  assign PECore_RunMac_if_and_675_rgt = (~ crossbar_spec_PE_Weight_WordType_16U_16U_for_land_11_lpi_1_dfm)
      & and_dcpl_705 & (fsm_output[2]);
  assign PECore_RunMac_if_and_676_rgt = crossbar_spec_PE_Weight_WordType_16U_16U_for_land_11_lpi_1_dfm
      & and_dcpl_705 & (fsm_output[2]);
  assign PECore_RunMac_if_and_685_cse = PECoreRun_wen & (PECore_RunMac_if_and_674_rgt
      | PECore_RunMac_if_and_675_rgt | PECore_RunMac_if_and_676_rgt);
  assign PECore_RunMac_if_and_627_rgt = (~ while_and_46_tmp_1) & and_dcpl_705 & (fsm_output[2]);
  assign PECore_RunMac_if_and_628_rgt = while_and_46_tmp_1 & and_dcpl_705 & (fsm_output[2]);
  assign PECore_RunMac_if_and_701_cse = PECoreRun_wen & (PECore_RunMac_if_and_674_rgt
      | PECore_RunMac_if_and_627_rgt | PECore_RunMac_if_and_628_rgt);
  assign PECore_RunMac_if_and_580_rgt = and_dcpl_705 & (fsm_output[2]);
  assign PECore_RunMac_if_and_717_cse = PECoreRun_wen & (PECore_RunMac_if_and_674_rgt
      | PECore_RunMac_if_and_580_rgt);
  assign PECore_RunMac_if_and_572_cse = (~(is_start_sva | state_2_0_sva_0)) & (fsm_output[2]);
  assign PECore_RunMac_if_and_569_rgt = and_dcpl_707 & (fsm_output[2]);
  assign PECore_RunMac_if_and_570_rgt = and_dcpl_709 & (fsm_output[2]);
  assign PECore_RunMac_if_and_571_rgt = state_2_0_sva_0 & (fsm_output[2]);
  assign PECore_RunMac_if_and_721_ssc = PECoreRun_wen & (~(((~ state_2_0_sva_0) &
      PECore_RunMac_if_or_5_m1c) | PECore_RunMac_if_and_572_cse));
  assign PECore_RunMac_if_or_145_m1c = (state_2_0_sva_0 & PECore_RunMac_if_or_5_m1c)
      | PECore_RunMac_if_and_571_rgt;
  assign PECore_RunMac_if_and_834_rgt = PECore_RunBias_if_for_and_45_rgt & PECore_RunMac_if_or_145_m1c;
  assign PECore_RunMac_if_and_867_cse = PECore_RunMac_if_and_721_ssc & (~((~ PECore_RunBias_if_for_and_45_rgt)
      & PECore_RunMac_if_or_145_m1c));
  assign PECore_RunMac_if_and_723_ssc = PECoreRun_wen & (~((fsm_output[4]) | (fsm_output[1])
      | PECore_RunMac_if_and_572_cse | ((~ state_2_0_sva_0) & (fsm_output[3]))));
  assign PECore_RunMac_if_or_143_m1c = PECore_RunMac_if_and_571_rgt | (state_2_0_sva_0
      & (fsm_output[3]));
  assign PECore_RunMac_if_and_726_cse = PECoreRun_wen & (PECore_RunMac_if_and_569_rgt
      | PECore_RunMac_if_and_570_rgt | PECore_RunMac_if_and_571_rgt);
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse = PECoreRun_wen & (~ (fsm_output[2]));
  assign PECore_RunBias_if_for_and_45_rgt = is_start_sva & (fsm_output[2]);
  assign PECore_RunBias_if_for_and_42_cse = (~ is_start_sva) & (fsm_output[2]);
  assign PECore_RunBias_if_for_and_34_rgt = is_start_sva & (fsm_output[1]);
  assign PECore_RunBias_if_for_and_cse = (~ is_start_sva) & (fsm_output[1]);
  assign act_port_reg_data_and_24_cse = PECoreRun_wen & (~ state_2_0_sva_0) & (fsm_output[2]);
  assign act_port_reg_data_and_enex5 = act_port_reg_data_and_24_cse & reg_act_port_reg_data_14_enexo;
  assign act_port_reg_data_and_28_enex5 = act_port_reg_data_and_24_cse & reg_act_port_reg_data_13_enexo;
  assign act_port_reg_data_and_29_enex5 = act_port_reg_data_and_24_cse & reg_act_port_reg_data_12_enexo;
  assign act_port_reg_data_and_30_enex5 = act_port_reg_data_and_24_cse & reg_act_port_reg_data_15_enexo;
  assign rva_out_reg_data_and_87_rgt = PECore_PushAxiRsp_if_asn_68 & (~ is_start_sva)
      & (fsm_output[2]);
  assign rva_out_reg_data_and_88_rgt = crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm
      & (~ is_start_sva) & (fsm_output[2]);
  assign rva_out_reg_data_and_91_cse = PECoreRun_wen & ((~ (fsm_output[2])) | rva_out_reg_data_and_87_rgt
      | rva_out_reg_data_and_88_rgt | PECore_RunMac_if_and_674_rgt | PECore_RunMac_if_and_580_rgt);
  assign pe_config_UpdateInputCounter_if_and_cse = PECoreRun_wen & (~ and_4616_cse);
  assign PECore_RunMac_if_and_820_rgt = state_2_0_sva_0 & is_start_sva & (fsm_output[2]);
  assign PECore_RunMac_if_and_872_cse = PECoreRun_wen & (~ (fsm_output[3]));
  assign PECore_RunMac_if_and_434_cse = pe_config_is_cluster_sva & (fsm_output[2]);
  assign PECore_RunMac_if_and_433_cse = (~ pe_config_is_cluster_sva) & (fsm_output[2]);
  assign PECore_RunMac_if_and_430_cse = (~ crossbar_spec_PE_Weight_WordType_16U_16U_for_land_9_lpi_1_dfm)
      & PECore_RunMac_if_and_433_cse;
  assign PECore_RunMac_if_and_431_cse = crossbar_spec_PE_Weight_WordType_16U_16U_for_land_9_lpi_1_dfm
      & PECore_RunMac_if_and_433_cse;
  assign PECore_RunMac_if_and_12_cse = (~ crossbar_spec_PE_Weight_WordType_16U_16U_for_land_9_lpi_1_dfm)
      & and_dcpl_705;
  assign PECore_RunMac_if_and_13_cse = crossbar_spec_PE_Weight_WordType_16U_16U_for_land_9_lpi_1_dfm
      & and_dcpl_705;
  assign PECore_RunMac_if_and_10_cse = (~ crossbar_spec_PE_Weight_WordType_16U_16U_for_land_9_lpi_1_dfm)
      & and_dcpl_709;
  assign PECore_RunMac_if_and_11_cse = crossbar_spec_PE_Weight_WordType_16U_16U_for_land_9_lpi_1_dfm
      & and_dcpl_709;
  assign PECore_RunMac_if_and_cse = PECoreRun_wen & and_dcpl_135 & (~ state_2_0_sva_0)
      & is_start_sva;
  assign PECore_RunMac_if_and_346_rgt = pe_config_is_cluster_sva & (~ (fsm_output[3]));
  assign or_796_cse = (~ input_read_req_valid_lpi_1_dfm_5) | input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_banks_write_if_for_if_mux_cse = MUX_v_128_2_2(input_mem_banks_bank_array_impl_data0_rsci_q_d,
      input_mem_banks_read_read_data_lpi_1, or_796_cse);
  assign and_5335_cse = reg_PECore_RunMac_asn_15_itm_1_ftd_1 & while_asn_41_itm_1;
  assign and_2979_cse = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]) & (fsm_output[1]);
  assign and_2983_cse = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14]) & (fsm_output[1]);
  assign and_2987_cse = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13]) & (fsm_output[1]);
  assign and_2991_cse = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12]) & (fsm_output[1]);
  assign and_2995_cse = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11]) & (fsm_output[1]);
  assign and_2999_cse = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[10]) & (fsm_output[1]);
  assign and_3003_cse = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[9]) & (fsm_output[1]);
  assign and_3007_cse = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8]) & (fsm_output[1]);
  assign and_3011_cse = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]) & (fsm_output[1]);
  assign and_3015_cse = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]) & (fsm_output[1]);
  assign and_3019_cse = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]) & (fsm_output[1]);
  assign and_3023_cse = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]) & (fsm_output[1]);
  assign and_3027_cse = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]) & (fsm_output[1]);
  assign and_3031_cse = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]) & (fsm_output[1]);
  assign and_3035_cse = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]) & (fsm_output[1]);
  assign and_3039_cse = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]) & (fsm_output[1]);
  assign or_1405_cse = weight_mem_read_arbxbar_xbar_for_3_1_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0])) & (fsm_output[1]);
  assign or_1409_cse = weight_mem_read_arbxbar_xbar_for_3_2_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1])) & (fsm_output[1]);
  assign or_1413_cse = weight_mem_read_arbxbar_xbar_for_3_3_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2])) & (fsm_output[1]);
  assign or_1417_cse = weight_mem_read_arbxbar_xbar_for_3_4_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3])) & (fsm_output[1]);
  assign or_1421_cse = weight_mem_read_arbxbar_xbar_for_3_5_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4])) & (fsm_output[1]);
  assign or_1425_cse = weight_mem_read_arbxbar_xbar_for_3_6_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5])) & (fsm_output[1]);
  assign or_1429_cse = weight_mem_read_arbxbar_xbar_for_3_7_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6])) & (fsm_output[1]);
  assign or_1433_cse = weight_mem_read_arbxbar_xbar_for_3_8_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7])) & (fsm_output[1]);
  assign or_1437_cse = weight_mem_read_arbxbar_xbar_for_3_9_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8])) & (fsm_output[1]);
  assign or_1441_cse = weight_mem_read_arbxbar_xbar_for_3_10_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[9])) & (fsm_output[1]);
  assign or_1445_cse = weight_mem_read_arbxbar_xbar_for_3_11_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[10])) & (fsm_output[1]);
  assign or_1449_cse = weight_mem_read_arbxbar_xbar_for_3_12_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11])) & (fsm_output[1]);
  assign or_1453_cse = weight_mem_read_arbxbar_xbar_for_3_13_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12])) & (fsm_output[1]);
  assign or_1457_cse = weight_mem_read_arbxbar_xbar_for_3_14_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13])) & (fsm_output[1]);
  assign or_1461_cse = weight_mem_read_arbxbar_xbar_for_3_15_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14])) & (fsm_output[1]);
  assign or_1465_cse = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[15])) & weight_mem_read_arbxbar_xbar_for_3_16_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      & (fsm_output[1]);
  assign nand_198_nl = ~(or_55_cse & or_1584_cse);
  assign nor_475_nl = ~(state_2_0_sva_2 | state_2_0_sva_1 | (~ input_port_PopNB_mioi_ivld_mxwt)
      | state_2_0_sva_0);
  assign mux_22_nl = MUX_s_1_2_2(nand_198_nl, nor_475_nl, is_start_sva);
  assign or_1183_cse = mux_22_nl & (fsm_output[1]);
  assign PECore_RunBias_if_accum_vector_out_data_6_lpi_1_dfm_mx2 = MUX_v_32_2_2(PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_4_sva,
      z_out_31, PECore_DecodeAxiRead_case_4_switch_lp_and_2_itm);
  assign PECore_RunBias_if_accum_vector_out_data_7_lpi_1_dfm_mx2 = MUX_v_32_2_2(PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_5_sva,
      z_out_32, PECore_DecodeAxiRead_case_4_switch_lp_and_2_itm);
  assign PECore_RunBias_if_accum_vector_out_data_10_lpi_1_dfm_mx2 = MUX_v_32_2_2(PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_1_sva,
      z_out_29, PECore_DecodeAxiRead_case_4_switch_lp_and_2_itm);
  assign PECore_RunBias_if_accum_vector_out_data_11_lpi_1_dfm_mx2 = MUX_v_32_2_2(PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_11_sva,
      z_out_30, PECore_DecodeAxiRead_case_4_switch_lp_and_2_itm);
  assign PECore_RunBias_if_for_11_operator_32_true_slc_operator_32_true_acc_13_svs_mx0
      = MUX_s_1_2_2(z_out_10_13, adpfloat_tmp_is_zero_land_10_lpi_1_dfm_st, or_dcpl_295);
  assign PECore_RunBias_if_for_10_operator_32_true_slc_operator_32_true_acc_13_svs_mx0
      = MUX_s_1_2_2(z_out_11_13, adpfloat_tmp_is_zero_land_10_lpi_1_dfm, or_dcpl_295);
  assign PECore_RunBias_if_for_7_operator_32_true_slc_operator_32_true_acc_13_svs_mx0
      = MUX_s_1_2_2(z_out_12_13, adpfloat_tmp_is_zero_land_11_lpi_1_dfm_st, or_dcpl_295);
  assign PECore_RunBias_if_for_6_operator_32_true_slc_operator_32_true_acc_13_svs_mx0
      = MUX_s_1_2_2(z_out_13_13, adpfloat_tmp_is_zero_land_11_lpi_1_dfm, or_dcpl_295);
  assign while_and_48_tmp_1 = PECore_RunFSM_switch_lp_equal_tmp_2 & is_start_sva;
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_15_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_15_lpi_1_dfm_3,
      PECore_RunMac_if_mux_136_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_1_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_0_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_0_lpi_1_dfm_3,
      PECore_RunMac_if_mux_136_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_14_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_14_lpi_1_dfm_3,
      PECore_RunMac_if_mux_136_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_2_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_1_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_1_lpi_1_dfm_3,
      PECore_RunMac_if_mux_136_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_13_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_13_lpi_1_dfm_3,
      PECore_RunMac_if_mux_136_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_3_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_2_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_2_lpi_1_dfm_3,
      PECore_RunMac_if_mux_136_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_13_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_12_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_12_lpi_1_dfm_3,
      PECore_RunMac_if_mux_136_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_4_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_3_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_3_lpi_1_dfm_3,
      PECore_RunMac_if_mux_136_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_12_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_11_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_11_lpi_1_dfm_3,
      PECore_RunMac_if_mux_136_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_5_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_4_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_4_lpi_1_dfm_3,
      PECore_RunMac_if_mux_136_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_11_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_10_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_10_lpi_1_dfm_3,
      PECore_RunMac_if_mux_136_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_6_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_5_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_5_lpi_1_dfm_3,
      PECore_RunMac_if_mux_136_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_10_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_9_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_9_lpi_1_dfm_3,
      PECore_RunMac_if_mux_136_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_7_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_6_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_6_lpi_1_dfm_3,
      PECore_RunMac_if_mux_136_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_9_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_8_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_8_lpi_1_dfm_3,
      PECore_RunMac_if_mux_136_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_8_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_7_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_7_lpi_1_dfm_3,
      PECore_RunMac_if_mux_136_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_15_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_15_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_126_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_1_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_0_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_0_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_126_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_14_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_14_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_126_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_2_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_1_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_1_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_126_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_13_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_13_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_126_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_3_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_2_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_2_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_126_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_13_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_12_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_12_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_126_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_4_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_3_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_3_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_126_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_12_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_11_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_11_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_126_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_5_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_4_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_4_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_126_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_11_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_10_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_10_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_126_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_6_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_5_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_5_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_126_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_10_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_9_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_9_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_126_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_7_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_6_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_6_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_126_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_9_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_8_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_8_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_126_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_8_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_7_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_7_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_126_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_15_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_15_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_125_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_14_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_14_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_125_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_15_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_15_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_124_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_15_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_15_lpi_1_dfm_3,
      PECore_RunMac_if_mux_134_itm[3:0]);
  assign weight_port_read_out_data_7_15_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_7_15_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm);
  assign weight_port_read_out_data_7_8_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_7_8_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm);
  assign weight_port_read_out_data_7_14_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_7_14_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm);
  assign weight_port_read_out_data_7_9_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_7_9_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm);
  assign weight_port_read_out_data_7_13_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_7_13_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm);
  assign weight_port_read_out_data_7_10_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_7_10_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm);
  assign weight_port_read_out_data_7_12_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_7_12_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm);
  assign weight_port_read_out_data_7_11_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_7_11_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm);
  assign weight_port_read_out_data_7_7_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_7_7_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm);
  assign weight_port_read_out_data_7_0_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_7_0_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm);
  assign weight_port_read_out_data_7_6_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_7_6_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm);
  assign weight_port_read_out_data_7_1_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_7_1_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm);
  assign weight_port_read_out_data_7_5_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_7_5_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm);
  assign weight_port_read_out_data_7_2_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_7_2_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm);
  assign weight_port_read_out_data_7_4_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_7_4_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm);
  assign weight_port_read_out_data_7_3_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_7_3_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm);
  assign weight_port_read_out_data_6_7_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_6_7_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm);
  assign weight_port_read_out_data_6_0_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_6_0_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm);
  assign weight_port_read_out_data_6_6_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_6_6_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm);
  assign weight_port_read_out_data_6_1_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_6_1_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm);
  assign weight_port_read_out_data_6_5_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_6_5_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm);
  assign weight_port_read_out_data_6_2_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_6_2_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm);
  assign weight_port_read_out_data_6_4_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_6_4_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm);
  assign weight_port_read_out_data_6_3_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_6_3_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm);
  assign weight_port_read_out_data_6_15_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_6_15_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm);
  assign weight_port_read_out_data_6_8_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_6_8_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm);
  assign weight_port_read_out_data_6_14_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_6_14_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm);
  assign weight_port_read_out_data_6_9_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_6_9_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm);
  assign weight_port_read_out_data_6_13_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_6_13_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm);
  assign weight_port_read_out_data_6_10_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_6_10_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm);
  assign weight_port_read_out_data_6_12_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_6_12_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm);
  assign weight_port_read_out_data_6_11_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_6_11_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm);
  assign weight_port_read_out_data_5_8_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_5_8_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm);
  assign weight_port_read_out_data_5_9_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_5_9_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm);
  assign weight_port_read_out_data_5_10_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_5_10_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm);
  assign weight_port_read_out_data_5_11_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_5_11_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm);
  assign weight_port_read_out_data_5_12_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_5_12_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm);
  assign weight_port_read_out_data_5_13_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_5_13_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm);
  assign weight_port_read_out_data_5_14_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_5_14_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_15_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_15_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_129_ftd_1);
  assign weight_port_read_out_data_5_15_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_5_15_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm);
  assign weight_port_read_out_data_4_0_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_4_0_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm);
  assign weight_port_read_out_data_4_1_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_4_1_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm);
  assign weight_port_read_out_data_4_2_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_4_2_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm);
  assign weight_port_read_out_data_4_3_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_4_3_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm);
  assign weight_port_read_out_data_4_4_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_4_4_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm);
  assign weight_port_read_out_data_4_5_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_4_5_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm);
  assign weight_port_read_out_data_4_6_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_4_6_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm);
  assign weight_port_read_out_data_4_7_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_4_7_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm);
  assign weight_port_read_out_data_4_8_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_4_8_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm);
  assign weight_port_read_out_data_4_9_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_4_9_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm);
  assign weight_port_read_out_data_4_10_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_4_10_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm);
  assign weight_port_read_out_data_4_11_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_4_11_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm);
  assign weight_port_read_out_data_4_12_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_4_12_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm);
  assign weight_port_read_out_data_4_13_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_4_13_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm);
  assign weight_port_read_out_data_4_14_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_4_14_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm);
  assign weight_port_read_out_data_4_15_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_4_15_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm);
  assign weight_port_read_out_data_3_8_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_3_8_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm);
  assign weight_port_read_out_data_3_9_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_3_9_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm);
  assign weight_port_read_out_data_3_10_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_3_10_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm);
  assign weight_port_read_out_data_3_11_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_3_11_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm);
  assign weight_port_read_out_data_3_12_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_3_12_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm);
  assign weight_port_read_out_data_3_13_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_3_13_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm);
  assign weight_port_read_out_data_3_14_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_3_14_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_15_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_15_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_128_ftd_1);
  assign weight_port_read_out_data_3_15_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_3_15_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm);
  assign weight_port_read_out_data_3_0_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_3_0_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm);
  assign weight_port_read_out_data_3_1_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_3_1_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm);
  assign weight_port_read_out_data_3_2_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_3_2_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm);
  assign weight_port_read_out_data_3_3_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_3_3_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm);
  assign weight_port_read_out_data_3_4_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_3_4_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm);
  assign weight_port_read_out_data_3_5_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_3_5_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm);
  assign weight_port_read_out_data_3_6_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_3_6_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm);
  assign weight_port_read_out_data_3_7_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_3_7_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm);
  assign weight_port_read_out_data_2_0_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_2_0_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm);
  assign weight_port_read_out_data_2_1_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_2_1_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm);
  assign weight_port_read_out_data_2_2_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_2_2_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm);
  assign weight_port_read_out_data_2_3_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_2_3_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm);
  assign weight_port_read_out_data_2_4_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_2_4_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm);
  assign weight_port_read_out_data_2_5_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_2_5_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm);
  assign weight_port_read_out_data_2_6_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_2_6_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm);
  assign weight_port_read_out_data_2_7_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_2_7_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm);
  assign weight_port_read_out_data_2_8_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_2_8_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm);
  assign weight_port_read_out_data_2_9_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_2_9_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm);
  assign weight_port_read_out_data_2_10_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_2_10_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm);
  assign weight_port_read_out_data_2_11_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_2_11_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm);
  assign weight_port_read_out_data_2_12_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_2_12_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm);
  assign weight_port_read_out_data_2_13_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_2_13_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm);
  assign weight_port_read_out_data_2_14_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_2_14_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm);
  assign weight_port_read_out_data_2_15_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_2_15_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm);
  assign weight_port_read_out_data_1_8_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_1_8_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm);
  assign weight_port_read_out_data_1_9_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_1_9_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm);
  assign weight_port_read_out_data_1_10_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_1_10_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm);
  assign weight_port_read_out_data_1_11_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_1_11_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm);
  assign weight_port_read_out_data_1_12_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_1_12_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm);
  assign weight_port_read_out_data_1_13_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_1_13_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm);
  assign weight_port_read_out_data_1_14_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_1_14_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_15_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_15_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_127_ftd_1);
  assign weight_port_read_out_data_1_15_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_1_15_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm);
  assign weight_port_read_out_data_1_0_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_1_0_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm);
  assign weight_port_read_out_data_1_1_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_1_1_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm);
  assign weight_port_read_out_data_1_2_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_1_2_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm);
  assign weight_port_read_out_data_1_3_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_1_3_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm);
  assign weight_port_read_out_data_1_4_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_1_4_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm);
  assign weight_port_read_out_data_1_5_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_1_5_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm);
  assign weight_port_read_out_data_1_6_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_1_6_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm);
  assign weight_port_read_out_data_1_7_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_1_7_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm);
  assign weight_port_read_out_data_0_8_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_0_8_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm);
  assign weight_port_read_out_data_0_9_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_0_9_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm);
  assign weight_port_read_out_data_0_10_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_0_10_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm);
  assign weight_port_read_out_data_0_11_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_0_11_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm);
  assign weight_port_read_out_data_0_12_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_0_12_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm);
  assign weight_port_read_out_data_0_13_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_0_13_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm);
  assign weight_port_read_out_data_0_14_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_0_14_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm);
  assign weight_port_read_out_data_0_15_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_0_15_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_2,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_1_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_0_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_0_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_123_ftd_1);
  assign weight_port_read_out_data_0_0_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_0_0_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_1_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm);
  assign weight_port_read_out_data_0_1_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_0_1_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_13_mx1w2,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm);
  assign weight_port_read_out_data_0_2_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_0_2_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_12_mx1w2,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm);
  assign weight_port_read_out_data_0_3_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_0_3_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_11_mx1w2,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm);
  assign weight_port_read_out_data_0_4_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_0_4_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm);
  assign weight_port_read_out_data_0_5_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_0_5_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm);
  assign weight_port_read_out_data_0_6_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_0_6_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm);
  assign weight_port_read_out_data_0_7_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_0_7_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm);
  assign rva_in_PopNB_mio_mrgout_dat_sva_1 = MUX_v_169_2_2(rva_in_PopNB_mioi_idat_mxwt,
      rva_in_PopNB_mio_mrgout_dat_sva, is_start_sva);
  assign PECore_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_mx1
      = MUX_s_1_2_2(rva_in_PopNB_mioi_ivld_mxwt, PECore_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva,
      is_start_sva);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm_mx1 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm,
      weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_sva_1, weight_mem_read_arbxbar_xbar_for_3_1_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm_mx1 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm,
      weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_sva_1, weight_mem_read_arbxbar_xbar_for_3_2_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm_mx1 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm,
      weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_sva_1, weight_mem_read_arbxbar_xbar_for_3_3_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm_mx1 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm,
      weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_sva_1, weight_mem_read_arbxbar_xbar_for_3_4_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm_mx1 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm,
      weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_sva_1, weight_mem_read_arbxbar_xbar_for_3_5_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm_mx1 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm,
      weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_sva_1, weight_mem_read_arbxbar_xbar_for_3_6_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm_mx1 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm,
      weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_sva_1, weight_mem_read_arbxbar_xbar_for_3_7_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm_mx1 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm,
      weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_sva_1, weight_mem_read_arbxbar_xbar_for_3_8_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm_mx1 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm,
      weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_sva_1, weight_mem_read_arbxbar_xbar_for_3_9_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm_mx1 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm,
      weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_sva_1, weight_mem_read_arbxbar_xbar_for_3_10_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm_mx1 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm,
      weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_sva_1, weight_mem_read_arbxbar_xbar_for_3_11_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm_mx1 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm,
      weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_sva_1, weight_mem_read_arbxbar_xbar_for_3_12_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm_mx1 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm,
      weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_sva_1, weight_mem_read_arbxbar_xbar_for_3_13_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm_mx1 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm,
      weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_sva_1, weight_mem_read_arbxbar_xbar_for_3_14_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm_mx1 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm,
      weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_sva_1, weight_mem_read_arbxbar_xbar_for_3_15_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_14
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_14,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_14,
      weight_mem_read_arbxbar_xbar_for_3_1_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_13
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_13,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_13,
      weight_mem_read_arbxbar_xbar_for_3_1_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_12
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_12,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_12,
      weight_mem_read_arbxbar_xbar_for_3_1_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_11
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_11,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_11,
      weight_mem_read_arbxbar_xbar_for_3_1_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_10
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_10,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_10,
      weight_mem_read_arbxbar_xbar_for_3_1_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_9
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_9,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_9,
      weight_mem_read_arbxbar_xbar_for_3_1_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_8
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_8,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_8,
      weight_mem_read_arbxbar_xbar_for_3_1_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_6
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_6,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_6,
      weight_mem_read_arbxbar_xbar_for_3_1_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_5
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_5,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_5,
      weight_mem_read_arbxbar_xbar_for_3_1_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_4
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_4,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_4,
      weight_mem_read_arbxbar_xbar_for_3_1_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_2
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_2,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_2,
      weight_mem_read_arbxbar_xbar_for_3_1_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_14
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_14,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_14,
      weight_mem_read_arbxbar_xbar_for_3_2_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_13
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_13,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_13,
      weight_mem_read_arbxbar_xbar_for_3_2_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_12
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_12,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_12,
      weight_mem_read_arbxbar_xbar_for_3_2_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_11
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_11,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_11,
      weight_mem_read_arbxbar_xbar_for_3_2_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_10
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_10,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_10,
      weight_mem_read_arbxbar_xbar_for_3_2_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_9
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_9,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_9,
      weight_mem_read_arbxbar_xbar_for_3_2_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_8
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_8,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_8,
      weight_mem_read_arbxbar_xbar_for_3_2_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_6
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_6,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_6,
      weight_mem_read_arbxbar_xbar_for_3_2_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_5
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_5,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_5,
      weight_mem_read_arbxbar_xbar_for_3_2_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_4
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_4,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_4,
      weight_mem_read_arbxbar_xbar_for_3_2_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_2
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_2,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_2,
      weight_mem_read_arbxbar_xbar_for_3_2_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_14
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_14,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_14,
      weight_mem_read_arbxbar_xbar_for_3_3_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_13
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_13,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_13,
      weight_mem_read_arbxbar_xbar_for_3_3_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_12
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_12,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_12,
      weight_mem_read_arbxbar_xbar_for_3_3_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_11
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_11,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_11,
      weight_mem_read_arbxbar_xbar_for_3_3_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_10
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_10,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_10,
      weight_mem_read_arbxbar_xbar_for_3_3_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_9
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_9,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_9,
      weight_mem_read_arbxbar_xbar_for_3_3_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_8
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_8,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_8,
      weight_mem_read_arbxbar_xbar_for_3_3_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_6
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_6,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_6,
      weight_mem_read_arbxbar_xbar_for_3_3_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_5
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_5,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_5,
      weight_mem_read_arbxbar_xbar_for_3_3_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_4
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_4,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_4,
      weight_mem_read_arbxbar_xbar_for_3_3_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_2
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_2,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_2,
      weight_mem_read_arbxbar_xbar_for_3_3_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_14
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_14,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_14,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_3_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_13
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_13,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_13,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_3_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_12
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_12,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_12,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_3_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_11
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_11,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_11,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_3_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_10
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_10,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_10,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_3_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_9
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_9,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_9,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_3_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_8
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_8,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_8,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_3_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_6
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_6,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_6,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_3_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_5
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_5,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_5,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_3_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_4
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_4,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_4,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_3_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_2
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_2,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_2,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_3_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_14
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_14,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_14,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_4_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_13
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_13,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_13,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_4_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_12
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_12,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_12,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_4_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_11
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_11,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_11,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_4_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_10
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_10,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_10,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_4_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_9
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_9,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_9,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_4_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_8
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_8,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_8,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_4_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_6
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_6,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_6,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_4_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_5
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_5,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_5,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_4_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_4
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_4,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_4,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_4_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_2
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_2,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_2,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_4_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_14
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_14,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_14,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_5_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_13
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_13,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_13,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_5_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_12
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_12,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_12,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_5_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_11
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_11,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_11,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_5_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_10
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_10,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_10,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_5_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_9
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_9,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_9,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_5_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_8
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_8,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_8,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_5_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_6
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_6,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_6,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_5_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_5
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_5,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_5,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_5_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_4
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_4,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_4,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_5_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_2
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_2,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_2,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_5_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_14
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_14,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_14,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_6_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_13
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_13,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_13,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_6_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_12
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_12,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_12,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_6_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_11
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_11,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_11,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_6_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_10
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_10,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_10,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_6_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_9
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_9,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_9,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_6_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_8
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_8,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_8,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_6_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_6
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_6,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_6,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_6_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_5
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_5,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_5,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_6_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_4
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_4,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_4,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_6_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_2
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_2,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_2,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_6_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_14
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_14,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_14,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_7_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_13
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_13,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_13,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_7_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_12
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_12,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_12,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_7_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_11
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_11,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_11,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_7_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_10
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_10,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_10,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_7_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_9
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_9,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_9,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_7_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_8
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_8,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_8,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_7_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_6
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_6,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_6,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_7_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_5
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_5,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_5,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_7_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_4
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_4,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_4,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_7_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_2
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_2,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_2,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_7_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_14
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_14,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_14,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_8_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_13
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_13,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_13,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_8_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_12
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_12,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_12,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_8_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_11
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_11,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_11,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_8_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_10
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_10,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_10,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_8_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_9
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_9,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_9,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_8_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_8
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_8,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_8,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_8_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_6
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_6,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_6,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_8_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_5
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_5,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_5,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_8_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_4
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_4,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_4,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_8_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_2
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_2,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_2,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_8_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_14
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_14,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_14,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_9_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_13
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_13,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_13,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_9_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_12
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_12,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_12,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_9_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_11
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_11,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_11,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_9_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_10
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_10,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_10,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_9_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_9
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_9,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_9,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_9_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_8
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_8,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_8,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_9_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_6
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_6,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_6,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_9_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_5
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_5,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_5,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_9_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_4
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_4,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_4,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_9_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_2
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_2,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_2,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_9_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_14
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_14,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_14,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_10_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_13
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_13,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_13,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_10_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_12
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_12,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_12,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_10_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_11
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_11,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_11,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_10_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_10
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_10,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_10,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_10_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_9
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_9,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_9,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_10_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_8
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_8,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_8,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_10_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_6
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_6,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_6,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_10_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_5
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_5,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_5,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_10_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_4
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_4,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_4,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_10_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_2
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_2,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_2,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_10_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_14
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_14,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_14,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_11_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_13
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_13,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_13,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_11_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_12
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_12,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_12,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_11_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_11
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_11,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_11,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_11_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_10
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_10,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_10,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_11_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_9
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_9,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_9,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_11_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_8
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_8,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_8,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_11_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_6
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_6,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_6,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_11_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_5
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_5,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_5,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_11_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_4
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_4,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_4,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_11_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_2
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_2,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_2,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_11_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_14
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_14,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_14,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_12_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_13
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_13,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_13,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_12_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_12
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_12,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_12,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_12_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_11
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_11,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_11,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_12_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_10
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_10,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_10,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_12_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_9
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_9,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_9,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_12_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_8
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_8,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_8,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_12_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_6
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_6,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_6,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_12_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_5
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_5,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_5,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_12_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_4
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_4,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_4,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_12_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_2
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_2,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_2,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_12_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_14
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_14,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_14,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_13_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_13
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_13,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_13,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_13_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_12
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_12,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_12,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_13_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_11
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_11,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_11,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_13_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_10
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_10,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_10,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_13_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_9
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_9,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_9,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_13_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_8
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_8,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_8,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_13_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_6
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_6,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_6,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_13_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_5
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_5,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_5,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_13_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_4
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_4,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_4,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_13_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_2
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_2,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_2,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_13_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_14
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_14,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_14,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_14_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_13
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_13,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_13,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_14_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_12
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_12,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_12,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_14_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_11
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_11,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_11,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_14_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_10
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_10,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_10,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_14_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_9
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_9,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_9,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_14_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_8
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_8,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_8,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_14_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_6
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_6,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_6,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_14_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_5
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_5,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_5,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_14_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_4
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_4,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_4,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_14_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_2
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_2,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_2,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_14_tmp);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_14
      = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_13
      = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_1,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_1_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_12
      = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_2,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_2_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_11
      = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_3,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_3_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_10
      = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_4,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_4_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_9
      = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_5,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_5_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_8
      = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_6,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_6_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_6
      = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_8,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_8_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_5
      = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_9,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_9_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_4
      = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_10,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_10_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_2
      = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_12,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_12_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0 = (rva_in_PopNB_mioi_idat_mxwt[151:148]==4'b0110);
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0 = (rva_in_PopNB_mioi_idat_mxwt[151:148]==4'b0101);
  assign adpfloat_tmp_is_zero_land_11_lpi_1_dfm_mx1w0 = ~((input_mem_banks_write_if_for_if_mux_cse[86:80]!=7'b0000000));
  assign adpfloat_tmp_is_zero_land_10_lpi_1_dfm_mx1w0 = ~((input_mem_banks_write_if_for_if_mux_cse[78:72]!=7'b0000000));
  assign adpfloat_tmp_is_zero_land_7_lpi_1_dfm_mx1w0 = ~((input_mem_banks_write_if_for_if_mux_cse[54:48]!=7'b0000000));
  assign adpfloat_tmp_is_zero_land_6_lpi_1_dfm_mx1w0 = ~((input_mem_banks_write_if_for_if_mux_cse[46:40]!=7'b0000000));
  assign PECore_RunBias_if_for_16_operator_32_true_slc_operator_32_true_acc_13_svs_mx1
      = MUX_s_1_2_2(z_out_10_13, PECore_RunBias_if_for_16_operator_32_true_slc_operator_32_true_acc_13_svs,
      or_dcpl_365);
  assign PECore_RunBias_if_for_15_operator_32_true_slc_operator_32_true_acc_13_svs_mx1
      = MUX_s_1_2_2(z_out_11_13, PECore_RunBias_if_for_15_operator_32_true_slc_operator_32_true_acc_13_svs,
      or_dcpl_365);
  assign PECore_RunBias_if_for_14_operator_32_true_slc_operator_32_true_acc_13_svs_mx1
      = MUX_s_1_2_2(z_out_12_13, PECore_RunBias_if_for_14_operator_32_true_slc_operator_32_true_acc_13_svs,
      or_dcpl_365);
  assign PECore_RunBias_if_for_13_operator_32_true_slc_operator_32_true_acc_13_svs_mx1
      = MUX_s_1_2_2(z_out_13_13, PECore_RunBias_if_for_13_operator_32_true_slc_operator_32_true_acc_13_svs,
      or_dcpl_365);
  assign PECore_RunBias_if_for_12_operator_32_true_slc_operator_32_true_acc_13_svs_mx2
      = MUX_s_1_2_2(z_out_11_13, PECore_RunBias_if_for_12_operator_32_true_slc_operator_32_true_acc_13_svs,
      or_dcpl_365);
  assign PECore_RunBias_if_for_1_operator_32_true_slc_operator_32_true_acc_13_svs_mx2
      = MUX_s_1_2_2(z_out_10_13, PECore_RunBias_if_for_1_operator_32_true_slc_operator_32_true_acc_13_svs,
      or_dcpl_365);
  assign PECore_RunBias_if_for_2_operator_32_true_slc_operator_32_true_acc_13_svs_mx2
      = MUX_s_1_2_2(z_out_10_13, PECore_RunBias_if_for_2_operator_32_true_slc_operator_32_true_acc_13_svs,
      or_dcpl_365);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_15_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_15_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_11_ftd_1);
  assign weight_port_read_out_data_5_0_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_5_0_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm);
  assign weight_port_read_out_data_5_1_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_5_1_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm);
  assign weight_port_read_out_data_5_2_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_5_2_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm);
  assign weight_port_read_out_data_5_3_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_5_3_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm);
  assign weight_port_read_out_data_5_4_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_5_4_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm);
  assign weight_port_read_out_data_5_5_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_5_5_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm);
  assign weight_port_read_out_data_5_6_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_5_6_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm);
  assign weight_port_read_out_data_5_7_sva_dfm_mx1 = MUX_v_8_2_2(weight_port_read_out_data_5_7_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm);
  assign PECore_RunMac_PECore_RunMac_and_2_cse = state_2_0_sva_2 & PECore_UpdateFSM_switch_lp_nor_6_cse;
  assign while_and_32_cse_1 = (~(PECore_RunFSM_switch_lp_equal_tmp_2 | PECore_RunMac_PECore_RunMac_and_2_cse
      | PECore_RunMac_nor_tmp)) & is_start_sva;
  assign PECore_RunBias_if_accum_vector_out_data_mux_5_cse = MUX_v_32_2_2(PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_1_sva,
      z_out_29, pe_config_is_bias_sva);
  assign PECore_RunBias_if_accum_vector_out_data_mux_7_cse = MUX_v_32_2_2(PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_11_sva,
      z_out_30, pe_config_is_bias_sva);
  assign PECore_RunBias_if_accum_vector_out_data_mux_9_cse = MUX_v_32_2_2(PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_4_sva,
      z_out_31, pe_config_is_bias_sva);
  assign PECore_RunBias_if_accum_vector_out_data_mux_11_cse = MUX_v_32_2_2(PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_5_sva,
      z_out_32, pe_config_is_bias_sva);
  assign input_mem_banks_load_store_for_else_and_cse_1 = input_read_req_valid_lpi_1_dfm_5
      & (~ input_write_req_valid_lpi_1_dfm_5);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm_1 = (weight_read_addrs_8_2_0_lpi_1_dfm_1[0])
      & PECore_RunFSM_switch_lp_equal_tmp_5 & weight_read_ack_10_lpi_1_dfm_15_mx0;
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm_1 = (weight_read_addrs_4_1_0_lpi_1_dfm_1[0])
      & weight_read_ack_2_lpi_1_dfm_15_mx0;
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm_1 = (weight_read_addrs_4_1_0_lpi_1_dfm_1[0])
      & weight_read_ack_6_lpi_1_dfm_15_mx0;
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm_1 = (weight_read_addrs_8_15_3_lpi_1_dfm_3[0])
      & weight_read_ack_8_lpi_1_dfm_15_mx0;
  assign PECore_RunFSM_switch_lp_equal_tmp_3 = ~(state_2_0_sva_2 | state_2_0_sva_1
      | state_2_0_sva_0);
  assign while_and_127_cse_1 = PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0 &
      (rva_in_PopNB_mio_mrgout_dat_sva_1[168]) & PECore_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_mx1
      & (~ is_start_sva);
  assign PECore_RunFSM_switch_lp_equal_tmp_4 = state_2_0_sva_1 & state_2_0_sva_0
      & (~ state_2_0_sva_2);
  assign PECore_RunFSM_switch_lp_nor_3_cse_1 = PECore_RunFSM_switch_lp_equal_tmp_5
      | PECore_RunFSM_switch_lp_equal_tmp_4;
  assign input_read_req_valid_lpi_1_dfm_6 = (pe_config_is_bias_sva & PECore_RunFSM_switch_lp_nor_3_cse_1)
      | PECore_RunFSM_switch_lp_equal_tmp_5;
  assign PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5 = (rva_in_PopNB_mioi_idat_mxwt[134])
      & (rva_in_PopNB_mioi_idat_mxwt[132]) & PECore_DecodeAxiWrite_case_4_switch_lp_nor_9_tmp;
  assign PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6 = (rva_in_PopNB_mioi_idat_mxwt[133])
      & PECore_DecodeAxiWrite_case_4_switch_lp_nor_15_tmp;
  assign PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7 = (rva_in_PopNB_mioi_idat_mxwt[133:132]==2'b11)
      & PECore_DecodeAxiWrite_case_4_switch_lp_nor_13_tmp;
  assign PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8 = (rva_in_PopNB_mioi_idat_mxwt[134])
      & PECore_DecodeAxiWrite_case_4_switch_lp_nor_11_tmp;
  assign PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_5 = (rva_in_PopNB_mioi_idat_mxwt[132])
      & PECore_DecodeAxiWrite_case_4_switch_lp_nor_7_tmp;
  assign PECore_DecodeAxiWrite_case_4_switch_lp_nor_tmp_1 = ~(PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_5
      | PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6 | PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7
      | PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8 | PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5);
  assign PECore_DecodeAxiRead_switch_lp_nor_tmp_mx0w0 = ~(PECore_DecodeAxiRead_switch_lp_equal_tmp_4
      | PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_31 | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0);
  assign PECore_DecodeAxiRead_switch_lp_nor_2_itm_mx0w0 = ~((rva_in_PopNB_mioi_idat_mxwt[151])
      | (rva_in_PopNB_mioi_idat_mxwt[149]) | (rva_in_PopNB_mioi_idat_mxwt[148]));
  assign PECore_RunFSM_switch_lp_equal_tmp_5 = state_2_0_sva_1 & (~(state_2_0_sva_2
      | state_2_0_sva_0));
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_13_cse_1 = ~(PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_5
      | PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6 | PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8
      | PECore_DecodeAxiWrite_case_4_switch_lp_nor_tmp_1);
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_12_cse_1 = ~(PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_5
      | PECore_DecodeAxiWrite_case_4_switch_lp_nor_tmp_1);
  assign PECore_DecodeAxiRead_switch_lp_nor_14_cse_1 = ~(PECore_DecodeAxiRead_switch_lp_equal_tmp_4
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0
      | PECore_DecodeAxiRead_switch_lp_nor_tmp_mx0w0);
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_4 = (rva_in_PopNB_mioi_idat_mxwt[151:148]==4'b0011);
  assign nl_PEManager_16U_GetWeightAddr_if_acc_2_psp_sva_1 = PEManager_16U_GetWeightAddr_if_acc_4_cmp_z
      + (PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx1[15:3]);
  assign PEManager_16U_GetWeightAddr_if_acc_2_psp_sva_1 = nl_PEManager_16U_GetWeightAddr_if_acc_2_psp_sva_1[12:0];
  assign PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx0_3_0
      = MUX_v_4_2_2((pe_manager_base_weight_0_sva[3:0]), (pe_manager_base_weight_1_sva[3:0]),
      pe_config_manager_counter_sva[0]);
  assign PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx1
      = MUX_v_16_2_2(pe_manager_base_weight_0_sva, pe_manager_base_weight_1_sva,
      pe_config_manager_counter_sva[0]);
  assign nl_PEManager_16U_GetWeightAddr_1_else_acc_2_psp_sva_1 = (PEManager_16U_GetWeightAddr_if_acc_4_cmp_z[11:0])
      + (PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx1[15:4]);
  assign PEManager_16U_GetWeightAddr_1_else_acc_2_psp_sva_1 = nl_PEManager_16U_GetWeightAddr_1_else_acc_2_psp_sva_1[11:0];
  assign pe_config_is_cluster_not_39_nl = ~ pe_config_is_cluster_sva;
  assign weight_read_addrs_8_2_0_lpi_1_dfm_1 = MUX_v_3_2_2(3'b000, (PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx0_3_0[2:0]),
      pe_config_is_cluster_not_39_nl);
  assign while_asn_294_mx0w0 = MUX_v_4_2_2(4'b0000, pe_config_manager_counter_sva,
      PECore_DecodeAxiWrite_case_4_switch_lp_or_6_cse_1);
  assign pe_config_manager_counter_sva_dfm_4_mx0_0 = MUX_s_1_2_2((while_asn_294_mx0w0[0]),
      (pe_config_manager_counter_sva[0]), or_dcpl_375);
  assign pe_config_manager_counter_sva_dfm_4_mx1 = MUX_v_4_2_2(while_asn_294_mx0w0,
      pe_config_manager_counter_sva, or_dcpl_375);
  assign pe_config_input_counter_sva_dfm_4_mx0 = MUX_v_8_2_2(({{7{PECore_DecodeAxiWrite_case_4_switch_lp_or_6_cse_1}},
      PECore_DecodeAxiWrite_case_4_switch_lp_or_6_cse_1}), pe_config_input_counter_sva,
      or_dcpl_724);
  assign pe_config_output_counter_sva_dfm_4_mx0 = MUX_v_8_2_2(({{7{PECore_DecodeAxiWrite_case_4_switch_lp_or_6_cse_1}},
      PECore_DecodeAxiWrite_case_4_switch_lp_or_6_cse_1}), pe_config_output_counter_sva,
      or_dcpl_724);
  assign PECore_DecodeAxiWrite_case_4_switch_lp_or_6_cse_1 = PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6
      | PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7 | PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8
      | PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5 | PECore_DecodeAxiWrite_case_4_switch_lp_nor_tmp_1;
  assign PECore_RunFSM_switch_lp_mux_28_nl = MUX_v_12_2_2(PEManager_16U_GetWeightAddr_1_else_acc_2_psp_sva_1,
      (PEManager_16U_GetWeightAddr_if_acc_2_psp_sva_1[12:1]), pe_config_is_cluster_sva);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_40_nl
      = MUX_v_12_2_2(12'b000000000000, PECore_RunFSM_switch_lp_mux_28_nl, PECore_RunFSM_switch_lp_equal_tmp_5);
  assign weight_read_addrs_0_15_4_lpi_1_dfm_5_mx0 = MUX_v_12_2_2((rva_in_PopNB_mio_mrgout_dat_sva_1[147:136]),
      PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_40_nl,
      or_dcpl_378);
  assign weight_read_addrs_4_1_0_lpi_1_dfm_1 = MUX_v_2_2_2(2'b00, (PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx1[1:0]),
      PECore_RunFSM_switch_lp_equal_tmp_5);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_43_nl
      = (PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx0_3_0[2])
      & PECore_RunFSM_switch_lp_equal_tmp_5;
  assign weight_read_addrs_0_2_0_lpi_1_dfm_4_2_mx0 = MUX_s_1_2_2((rva_in_PopNB_mio_mrgout_dat_sva_1[134]),
      PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_43_nl,
      or_dcpl_378);
  assign weight_read_addrs_0_2_0_lpi_1_dfm_4_1_mx0 = MUX_s_1_2_2((rva_in_PopNB_mio_mrgout_dat_sva_1[133]),
      (weight_read_addrs_4_1_0_lpi_1_dfm_1[1]), or_dcpl_378);
  assign weight_read_addrs_0_2_0_lpi_1_dfm_4_0_mx0 = MUX_s_1_2_2((rva_in_PopNB_mio_mrgout_dat_sva_1[132]),
      (weight_read_addrs_4_1_0_lpi_1_dfm_1[0]), or_dcpl_378);
  assign PECore_RunFSM_switch_lp_mux_29_nl = MUX_s_1_2_2((PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx0_3_0[3]),
      (PEManager_16U_GetWeightAddr_if_acc_2_psp_sva_1[0]), pe_config_is_cluster_sva);
  assign weight_read_addrs_0_3_lpi_1_dfm_6 = PECore_RunFSM_switch_lp_mux_29_nl &
      PECore_RunFSM_switch_lp_equal_tmp_5;
  assign Arbiter_16U_Roundrobin_pick_mux_3212_nl = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_7,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_7_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_2_3_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3212_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_14;
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1_3 = weight_read_addrs_0_3_lpi_1_dfm_5_mx0
      & weight_read_ack_0_lpi_1_dfm_15_mx0;
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1_2 = weight_read_addrs_0_2_0_lpi_1_dfm_4_2_mx0
      & weight_read_ack_0_lpi_1_dfm_15_mx0;
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1_1 = weight_read_addrs_0_2_0_lpi_1_dfm_4_1_mx0
      & weight_read_ack_0_lpi_1_dfm_15_mx0;
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1_0 = weight_read_addrs_0_2_0_lpi_1_dfm_4_0_mx0
      & weight_read_ack_0_lpi_1_dfm_15_mx0;
  assign weight_mem_run_1_if_for_if_and_stg_2_0_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_3_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_0_1_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_1_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_4_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_0_2_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_2_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_5_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_0_3_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_3_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_6_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_0_4_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_4_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_7_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_0_5_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_5_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_8_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_0_6_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_6_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_9_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_0_7_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_7_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_10_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_0_8_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_8_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_11_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_0_9_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_9_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_12_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_0_10_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_10_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_13_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_0_11_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_11_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_14_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_0_12_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_12_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_15_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_0_13_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_13_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_16_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_0_14_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_14_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_17_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_702_nl = weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_224_tmp
      & (~(weight_mem_run_1_if_for_if_and_stg_2_0_15_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_2_3_sva_1)));
  assign weight_read_ack_0_lpi_1_dfm_15_mx0 = MUX_s_1_2_2(weight_mem_run_1_if_for_if_and_702_nl,
      weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_224_tmp, or_dcpl_34);
  assign weight_mem_run_1_if_for_if_and_stg_2_0_15_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_15_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_2_2_sva_1);
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_224_tmp = weight_read_req_valid_0_lpi_1_dfm_4_mx0
      & (Arbiter_16U_Roundrobin_pick_return_0_1_lpi_1_dfm_2 | Arbiter_16U_Roundrobin_pick_return_0_2_lpi_1_dfm_2
      | Arbiter_16U_Roundrobin_pick_return_0_3_lpi_1_dfm_2 | Arbiter_16U_Roundrobin_pick_return_0_4_lpi_1_dfm_2
      | Arbiter_16U_Roundrobin_pick_return_0_5_lpi_1_dfm_2 | Arbiter_16U_Roundrobin_pick_return_0_6_lpi_1_dfm_2
      | Arbiter_16U_Roundrobin_pick_return_0_7_lpi_1_dfm_2 | Arbiter_16U_Roundrobin_pick_return_0_8_lpi_1_dfm_2
      | Arbiter_16U_Roundrobin_pick_return_0_9_lpi_1_dfm_2 | Arbiter_16U_Roundrobin_pick_return_0_10_lpi_1_dfm_2
      | Arbiter_16U_Roundrobin_pick_return_0_11_lpi_1_dfm_2 | Arbiter_16U_Roundrobin_pick_return_0_12_lpi_1_dfm_2
      | Arbiter_16U_Roundrobin_pick_return_0_13_lpi_1_dfm_2 | Arbiter_16U_Roundrobin_pick_return_0_14_lpi_1_dfm_2
      | Arbiter_16U_Roundrobin_pick_return_0_15_lpi_1_dfm_2 | Arbiter_16U_Roundrobin_pick_return_0_lpi_1_dfm_2)
      & (~(weight_mem_run_1_if_for_if_and_stg_2_0_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_1_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_0_1_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_2_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_0_2_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_3_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_0_3_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_4_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_0_4_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_5_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_0_5_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_6_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_0_6_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_7_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_0_7_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_8_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_0_8_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_9_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_0_9_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_10_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_0_10_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_11_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_0_11_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_12_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_0_12_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_13_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_0_13_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_14_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_0_14_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_15_lpi_1_dfm_1));
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_tmp = MUX_s_1_16_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[9]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[10]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]), {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1_3
      , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1_2 , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1_1
      , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1_0});
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_mux_5_nl =
      MUX_s_1_2_2(weight_read_addrs_0_3_lpi_1_dfm_6, (rva_in_PopNB_mioi_idat_mxwt[135]),
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0);
  assign PECore_DecodeAxi_if_mux_122_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_mux_5_nl,
      weight_read_addrs_0_3_lpi_1_dfm_6, rva_in_PopNB_mioi_idat_mxwt[168]);
  assign PECore_DecodeAxi_mux_134_nl = MUX_s_1_2_2(weight_read_addrs_0_3_lpi_1_dfm_6,
      PECore_DecodeAxi_if_mux_122_nl, rva_in_PopNB_mioi_ivld_mxwt);
  assign weight_read_addrs_0_3_lpi_1_dfm_5_mx0 = MUX_s_1_2_2(PECore_DecodeAxi_mux_134_nl,
      weight_read_addrs_0_3_lpi_1_dfm_6, is_start_sva);
  assign weight_mem_run_1_if_for_land_1_lpi_1_dfm_1 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0])
      & weight_mem_read_arbxbar_xbar_for_3_1_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  assign weight_mem_run_1_if_for_land_2_lpi_1_dfm_1 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1])
      & weight_mem_read_arbxbar_xbar_for_3_2_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  assign weight_mem_run_1_if_for_land_3_lpi_1_dfm_1 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2])
      & weight_mem_read_arbxbar_xbar_for_3_3_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  assign weight_mem_run_1_if_for_land_4_lpi_1_dfm_1 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3])
      & weight_mem_read_arbxbar_xbar_for_3_4_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  assign weight_mem_run_1_if_for_land_5_lpi_1_dfm_1 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4])
      & weight_mem_read_arbxbar_xbar_for_3_5_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  assign weight_mem_run_1_if_for_land_6_lpi_1_dfm_1 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5])
      & weight_mem_read_arbxbar_xbar_for_3_6_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  assign weight_mem_run_1_if_for_land_7_lpi_1_dfm_1 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6])
      & weight_mem_read_arbxbar_xbar_for_3_7_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  assign weight_mem_run_1_if_for_land_8_lpi_1_dfm_1 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7])
      & weight_mem_read_arbxbar_xbar_for_3_8_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  assign weight_mem_run_1_if_for_land_9_lpi_1_dfm_1 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8])
      & weight_mem_read_arbxbar_xbar_for_3_9_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  assign weight_mem_run_1_if_for_land_10_lpi_1_dfm_1 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[9])
      & weight_mem_read_arbxbar_xbar_for_3_10_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  assign weight_mem_run_1_if_for_land_11_lpi_1_dfm_1 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[10])
      & weight_mem_read_arbxbar_xbar_for_3_11_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  assign weight_mem_run_1_if_for_land_12_lpi_1_dfm_1 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11])
      & weight_mem_read_arbxbar_xbar_for_3_12_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  assign weight_mem_run_1_if_for_land_13_lpi_1_dfm_1 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12])
      & weight_mem_read_arbxbar_xbar_for_3_13_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  assign weight_mem_run_1_if_for_land_14_lpi_1_dfm_1 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13])
      & weight_mem_read_arbxbar_xbar_for_3_14_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  assign weight_mem_run_1_if_for_land_15_lpi_1_dfm_1 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14])
      & weight_mem_read_arbxbar_xbar_for_3_15_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_or_nl
      = PECore_RunFSM_switch_lp_equal_tmp_5 | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
  assign PECore_DecodeAxi_if_mux_123_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_or_nl,
      PECore_RunFSM_switch_lp_equal_tmp_5, rva_in_PopNB_mioi_idat_mxwt[168]);
  assign PECore_DecodeAxi_mux_135_nl = MUX_s_1_2_2(PECore_RunFSM_switch_lp_equal_tmp_5,
      PECore_DecodeAxi_if_mux_123_nl, rva_in_PopNB_mioi_ivld_mxwt);
  assign weight_read_req_valid_0_lpi_1_dfm_4_mx0 = MUX_s_1_2_2(PECore_DecodeAxi_mux_135_nl,
      PECore_RunFSM_switch_lp_equal_tmp_5, is_start_sva);
  assign Arbiter_16U_Roundrobin_pick_return_0_1_lpi_1_dfm_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_1_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_return_0_2_lpi_1_dfm_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_1
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_2_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_return_0_3_lpi_1_dfm_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_2
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_return_0_4_lpi_1_dfm_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_3
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_4_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_return_0_5_lpi_1_dfm_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_4
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_5_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_return_0_6_lpi_1_dfm_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_5
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_6_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_return_0_7_lpi_1_dfm_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_6
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_7_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_return_0_8_lpi_1_dfm_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_7
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_8_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_return_0_9_lpi_1_dfm_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_8
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_9_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_return_0_10_lpi_1_dfm_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_9
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_10_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_return_0_11_lpi_1_dfm_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_10
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_11_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_return_0_12_lpi_1_dfm_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_11
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_12_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_return_0_13_lpi_1_dfm_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_12
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_13_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_return_0_14_lpi_1_dfm_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_13
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_14_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_return_0_15_lpi_1_dfm_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_14
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_15_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_return_0_lpi_1_dfm_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_15
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_lpi_1_dfm_mx0;
  assign or_1624_nl = or_dcpl | state_2_0_sva_2;
  assign PECore_RunFSM_case_0_if_mux_1_nl = MUX_s_1_2_2(input_port_PopNB_mioi_ivld_mxwt,
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva,
      or_1624_nl);
  assign input_write_req_valid_lpi_1_dfm_6 = PECore_RunFSM_case_0_if_mux_1_nl & PECore_RunFSM_switch_lp_equal_tmp_3;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_14
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14 & weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14 & (~ weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_13
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13 & weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13 & (~ weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_12
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12 & weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12 & (~ weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_11
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11 & weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11 & (~ weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_10
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10 & weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10 & (~ weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_9
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9 & weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9 & (~ weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_8
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8 & weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8 & (~ weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_7
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7 & weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7 & (~ weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_6
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6 & weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6 & (~ weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_5
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5 & weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5 & (~ weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_4
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4 & weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4 & (~ weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_3
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3 & weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3 & (~ weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_2
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2 & weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2 & (~ weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_1
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1 & weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1 & (~ weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_0
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0 & weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0 & (~ weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_nl
      = Arbiter_16U_Roundrobin_pick_priority_29_1_sva_1 & (~ Arbiter_16U_Roundrobin_pick_priority_30_1_sva_1);
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_465_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_1_sva_1) & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_450_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_466_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_1_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_450_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_468_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_1_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_452_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_469_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_1_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_452_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_470_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_1_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_453_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_471_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_1_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_453_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_472_nl
      = (~ operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_454_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_473_nl
      = operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_454_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_474_nl
      = (~ operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_455_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_475_nl
      = operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_455_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_476_nl
      = (~ operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_1_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_456_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_477_nl
      = operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_1_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_456_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_478_nl
      = (~ operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_457_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_479_nl
      = operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_457_cse;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_15_2(Arbiter_16U_Roundrobin_pick_priority_25_1_sva_1, Arbiter_16U_Roundrobin_pick_priority_27_1_sva_1,
      nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_nl,
      Arbiter_16U_Roundrobin_pick_priority_17_1_sva_1, Arbiter_16U_Roundrobin_pick_priority_19_1_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_21_1_sva_1, Arbiter_16U_Roundrobin_pick_priority_23_1_sva_1,
      (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[0]), (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[0]),
      (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[0]), (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]),
      (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[0]), (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[0]),
      (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[0]), (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[0]),
      {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_465_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_466_nl
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_1_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_468_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_469_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_470_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_471_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_472_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_473_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_474_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_475_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_476_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_477_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_478_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_479_nl});
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_450_cse
      = (~ operator_3_false_operator_3_false_operator_3_false_or_mdf_1_sva_1) & weight_mem_read_arbxbar_xbar_for_3_1_operator_7_false_operator_7_false_operator_7_false_or_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_452_cse
      = (~ operator_4_false_operator_4_false_operator_4_false_or_mdf_1_sva_1) & and_dcpl_725;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_453_cse
      = operator_4_false_operator_4_false_operator_4_false_or_mdf_1_sva_1 & and_dcpl_725;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_454_cse
      = (~ operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_1_sva_1)
      & and_dcpl_726;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_455_cse
      = operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_1_sva_1 &
      and_dcpl_726;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_456_cse
      = (~ operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_1_sva_1)
      & and_dcpl_733;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_457_cse
      = operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_1_sva_1 &
      and_dcpl_733;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_8_2(operator_2_false_operator_2_false_operator_2_false_or_mdf_1_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_30_1_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_1_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_1_sva_1, operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1,
      operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1, operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_1_sva_1,
      operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1, {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_450_cse
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_1_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_452_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_453_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_454_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_455_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_456_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_457_cse});
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(operator_3_false_operator_3_false_operator_3_false_or_mdf_1_sva_1,
      operator_4_false_operator_4_false_operator_4_false_or_mdf_1_sva_1, operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_1_sva_1,
      operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_1_sva_1, {weight_mem_read_arbxbar_xbar_for_3_1_operator_7_false_operator_7_false_operator_7_false_or_cse
      , and_dcpl_725 , and_dcpl_726 , and_dcpl_733});
  assign weight_mem_read_arbxbar_xbar_for_3_1_operator_7_false_operator_7_false_operator_7_false_or_cse
      = Arbiter_16U_Roundrobin_pick_priority_30_1_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_1_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_1_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_1_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_1_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_1_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_1_sva_1;
  assign weight_mem_read_arbxbar_xbar_for_3_1_operator_8_false_operator_8_false_operator_8_false_or_nl
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[0]);
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_1_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_1_operator_8_false_operator_8_false_operator_8_false_or_nl,
      weight_mem_read_arbxbar_xbar_for_3_1_operator_7_false_operator_7_false_operator_7_false_or_cse,
      weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign Arbiter_16U_Roundrobin_pick_priority_25_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_10_sva
      & (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[0]);
  assign Arbiter_16U_Roundrobin_pick_priority_27_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_12_sva
      & (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[0]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_1_sva_1 = Arbiter_16U_Roundrobin_pick_priority_27_1_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_1_sva_1;
  assign operator_3_false_operator_3_false_operator_3_false_or_mdf_1_sva_1 = Arbiter_16U_Roundrobin_pick_priority_30_1_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_29_1_sva_1 | Arbiter_16U_Roundrobin_pick_priority_28_1_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_29_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_14_sva
      & (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[0]);
  assign Arbiter_16U_Roundrobin_pick_priority_30_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_15_sva
      & (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[0]);
  assign Arbiter_16U_Roundrobin_pick_priority_26_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_11_sva
      & (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[0]);
  assign Arbiter_16U_Roundrobin_pick_priority_28_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_13_sva
      & (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[0]);
  assign Arbiter_16U_Roundrobin_pick_priority_21_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_6_sva
      & (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[0]);
  assign Arbiter_16U_Roundrobin_pick_priority_23_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_8_sva
      & (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[0]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_1_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_23_1_sva_1 | Arbiter_16U_Roundrobin_pick_priority_22_1_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_17_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_2_sva
      & (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[0]);
  assign Arbiter_16U_Roundrobin_pick_priority_19_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_4_sva
      & (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[0]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_1_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_19_1_sva_1 | Arbiter_16U_Roundrobin_pick_priority_18_1_sva_1;
  assign operator_4_false_operator_4_false_operator_4_false_or_mdf_1_sva_1 = Arbiter_16U_Roundrobin_pick_priority_23_1_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_1_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_1_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_1_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_22_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_7_sva
      & (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[0]);
  assign Arbiter_16U_Roundrobin_pick_priority_18_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_3_sva
      & (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[0]);
  assign Arbiter_16U_Roundrobin_pick_priority_20_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_5_sva
      & (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[0]);
  assign Arbiter_16U_Roundrobin_pick_priority_24_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_9_sva
      & (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[0]);
  assign operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[0]);
  assign operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1
      = (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[0]);
  assign operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_1_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[0]);
  assign operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[0]);
  assign operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_1_sva_1
      = (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[0]);
  assign operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_1_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[0]);
  assign weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp
      = Arbiter_16U_Roundrobin_pick_priority_30_1_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_1_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_1_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_1_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_1_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_1_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_1_sva_1 | Arbiter_16U_Roundrobin_pick_priority_23_1_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_1_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_1_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_1_sva_1 | Arbiter_16U_Roundrobin_pick_priority_19_1_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_18_1_sva_1 | Arbiter_16U_Roundrobin_pick_priority_17_1_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_0_1_sva & (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[0]));
  assign Arbiter_16U_Roundrobin_pick_mux_2995_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_0,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_0,
      weight_mem_read_arbxbar_xbar_for_3_1_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_3_0_sva_1 = Arbiter_16U_Roundrobin_pick_mux_2995_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_2994_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_1,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_1,
      weight_mem_read_arbxbar_xbar_for_3_1_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_3_1_sva_1 = Arbiter_16U_Roundrobin_pick_mux_2994_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_2992_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_3,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_3,
      weight_mem_read_arbxbar_xbar_for_3_1_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_3_2_sva_1 = Arbiter_16U_Roundrobin_pick_mux_2992_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_2988_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_7,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_7,
      weight_mem_read_arbxbar_xbar_for_3_1_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_sva_1 = Arbiter_16U_Roundrobin_pick_mux_2988_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_14;
  assign nl_operator_16_false_1_acc_12_nl = operator_16_false_1_mux_16_cse + 16'b0000000000000001;
  assign operator_16_false_1_acc_12_nl = nl_operator_16_false_1_acc_12_nl[15:0];
  assign weight_read_addrs_1_lpi_1_dfm_2 = MUX_v_16_2_2(16'b0000000000000000, operator_16_false_1_acc_12_nl,
      PECore_RunFSM_switch_lp_equal_tmp_5);
  assign nl_operator_16_false_1_acc_nl = ({operator_16_false_1_mux_10_cse , operator_16_false_1_mux_14_cse
      , (PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx1[2:1])})
      + 15'b000000000000001;
  assign operator_16_false_1_acc_nl = nl_operator_16_false_1_acc_nl[14:0];
  assign weight_read_addrs_2_15_1_lpi_1_dfm_2 = MUX_v_15_2_2(15'b000000000000000,
      operator_16_false_1_acc_nl, PECore_RunFSM_switch_lp_equal_tmp_5);
  assign nl_operator_16_false_1_acc_11_nl = operator_16_false_1_mux_16_cse + 16'b0000000000000011;
  assign operator_16_false_1_acc_11_nl = nl_operator_16_false_1_acc_11_nl[15:0];
  assign weight_read_addrs_3_lpi_1_dfm_2 = MUX_v_16_2_2(16'b0000000000000000, operator_16_false_1_acc_11_nl,
      PECore_RunFSM_switch_lp_equal_tmp_5);
  assign operator_16_false_1_mux_20_nl = MUX_v_14_2_2(({PEManager_16U_GetWeightAddr_1_else_acc_2_psp_sva_1
      , (PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx1[3:2])}),
      ({PEManager_16U_GetWeightAddr_if_acc_2_psp_sva_1 , (PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx0_3_0[2])}),
      and_5541_cse);
  assign nl_operator_16_false_1_acc_8_nl = operator_16_false_1_mux_20_nl + 14'b00000000000001;
  assign operator_16_false_1_acc_8_nl = nl_operator_16_false_1_acc_8_nl[13:0];
  assign weight_read_addrs_4_15_2_lpi_1_dfm_2 = MUX_v_14_2_2(14'b00000000000000,
      operator_16_false_1_acc_8_nl, PECore_RunFSM_switch_lp_equal_tmp_5);
  assign nl_operator_16_false_1_acc_10_nl = operator_16_false_1_mux_16_cse + 16'b0000000000000101;
  assign operator_16_false_1_acc_10_nl = nl_operator_16_false_1_acc_10_nl[15:0];
  assign weight_read_addrs_5_lpi_1_dfm_2 = MUX_v_16_2_2(16'b0000000000000000, operator_16_false_1_acc_10_nl,
      PECore_RunFSM_switch_lp_equal_tmp_5);
  assign nl_operator_16_false_1_acc_7_nl = ({operator_16_false_1_mux_10_cse , operator_16_false_1_mux_14_cse
      , (PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx1[2:1])})
      + 15'b000000000000011;
  assign operator_16_false_1_acc_7_nl = nl_operator_16_false_1_acc_7_nl[14:0];
  assign weight_read_addrs_6_15_1_lpi_1_dfm_2 = MUX_v_15_2_2(15'b000000000000000,
      operator_16_false_1_acc_7_nl, PECore_RunFSM_switch_lp_equal_tmp_5);
  assign nl_operator_16_false_1_acc_9_nl = operator_16_false_1_mux_16_cse + 16'b0000000000000111;
  assign operator_16_false_1_acc_9_nl = nl_operator_16_false_1_acc_9_nl[15:0];
  assign weight_read_addrs_7_lpi_1_dfm_2 = MUX_v_16_2_2(16'b0000000000000000, operator_16_false_1_acc_9_nl,
      PECore_RunFSM_switch_lp_equal_tmp_5);
  assign nl_operator_16_false_1_acc_3_nl = ({PEManager_16U_GetWeightAddr_1_else_acc_2_psp_sva_1
      , (PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx0_3_0[3])})
      + 13'b0000000000001;
  assign operator_16_false_1_acc_3_nl = nl_operator_16_false_1_acc_3_nl[12:0];
  assign weight_read_addrs_8_15_3_lpi_1_dfm_3 = operator_16_false_1_acc_3_nl & (signext_13_1(~
      pe_config_is_cluster_sva)) & ({{12{PECore_RunFSM_switch_lp_equal_tmp_5}}, PECore_RunFSM_switch_lp_equal_tmp_5});
  assign nl_PECore_RunFSM_case_2_else_for_10_operator_16_false_1_acc_nl = ({PEManager_16U_GetWeightAddr_1_else_acc_2_psp_sva_1
      , (PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx1[3:0])})
      + 16'b0000000000001001;
  assign PECore_RunFSM_case_2_else_for_10_operator_16_false_1_acc_nl = nl_PECore_RunFSM_case_2_else_for_10_operator_16_false_1_acc_nl[15:0];
  assign weight_read_addrs_9_lpi_1_dfm_3 = PECore_RunFSM_case_2_else_for_10_operator_16_false_1_acc_nl
      & (signext_16_1(~ pe_config_is_cluster_sva)) & ({{15{PECore_RunFSM_switch_lp_equal_tmp_5}},
      PECore_RunFSM_switch_lp_equal_tmp_5});
  assign nl_operator_16_false_1_acc_4_nl = ({PEManager_16U_GetWeightAddr_1_else_acc_2_psp_sva_1
      , (PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx1[3:1])})
      + 15'b000000000000101;
  assign operator_16_false_1_acc_4_nl = nl_operator_16_false_1_acc_4_nl[14:0];
  assign weight_read_addrs_10_15_1_lpi_1_dfm_3 = operator_16_false_1_acc_4_nl & (signext_15_1(~
      pe_config_is_cluster_sva)) & ({{14{PECore_RunFSM_switch_lp_equal_tmp_5}}, PECore_RunFSM_switch_lp_equal_tmp_5});
  assign nl_PECore_RunFSM_case_2_else_for_12_operator_16_false_1_acc_nl = ({PEManager_16U_GetWeightAddr_1_else_acc_2_psp_sva_1
      , (PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx1[3:0])})
      + 16'b0000000000001011;
  assign PECore_RunFSM_case_2_else_for_12_operator_16_false_1_acc_nl = nl_PECore_RunFSM_case_2_else_for_12_operator_16_false_1_acc_nl[15:0];
  assign weight_read_addrs_11_lpi_1_dfm_3 = PECore_RunFSM_case_2_else_for_12_operator_16_false_1_acc_nl
      & (signext_16_1(~ pe_config_is_cluster_sva)) & ({{15{PECore_RunFSM_switch_lp_equal_tmp_5}},
      PECore_RunFSM_switch_lp_equal_tmp_5});
  assign nl_operator_16_false_1_acc_5_nl = ({PEManager_16U_GetWeightAddr_1_else_acc_2_psp_sva_1
      , (PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx1[3:2])})
      + 14'b00000000000011;
  assign operator_16_false_1_acc_5_nl = nl_operator_16_false_1_acc_5_nl[13:0];
  assign weight_read_addrs_12_15_2_lpi_1_dfm_3 = operator_16_false_1_acc_5_nl & (signext_14_1(~
      pe_config_is_cluster_sva)) & ({{13{PECore_RunFSM_switch_lp_equal_tmp_5}}, PECore_RunFSM_switch_lp_equal_tmp_5});
  assign nl_PECore_RunFSM_case_2_else_for_14_operator_16_false_1_acc_nl = ({PEManager_16U_GetWeightAddr_1_else_acc_2_psp_sva_1
      , (PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx1[3:0])})
      + 16'b0000000000001101;
  assign PECore_RunFSM_case_2_else_for_14_operator_16_false_1_acc_nl = nl_PECore_RunFSM_case_2_else_for_14_operator_16_false_1_acc_nl[15:0];
  assign weight_read_addrs_13_lpi_1_dfm_3 = PECore_RunFSM_case_2_else_for_14_operator_16_false_1_acc_nl
      & (signext_16_1(~ pe_config_is_cluster_sva)) & ({{15{PECore_RunFSM_switch_lp_equal_tmp_5}},
      PECore_RunFSM_switch_lp_equal_tmp_5});
  assign nl_operator_16_false_1_acc_6_nl = ({PEManager_16U_GetWeightAddr_1_else_acc_2_psp_sva_1
      , (PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx1[3:1])})
      + 15'b000000000000111;
  assign operator_16_false_1_acc_6_nl = nl_operator_16_false_1_acc_6_nl[14:0];
  assign weight_read_addrs_14_15_1_lpi_1_dfm_3 = operator_16_false_1_acc_6_nl & (signext_15_1(~
      pe_config_is_cluster_sva)) & ({{14{PECore_RunFSM_switch_lp_equal_tmp_5}}, PECore_RunFSM_switch_lp_equal_tmp_5});
  assign nl_PECore_RunFSM_case_2_else_for_16_operator_16_false_1_acc_nl = ({PEManager_16U_GetWeightAddr_1_else_acc_2_psp_sva_1
      , (PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx1[3:0])})
      + 16'b0000000000001111;
  assign PECore_RunFSM_case_2_else_for_16_operator_16_false_1_acc_nl = nl_PECore_RunFSM_case_2_else_for_16_operator_16_false_1_acc_nl[15:0];
  assign weight_read_addrs_15_lpi_1_dfm_3 = PECore_RunFSM_case_2_else_for_16_operator_16_false_1_acc_nl
      & (signext_16_1(~ pe_config_is_cluster_sva)) & ({{15{PECore_RunFSM_switch_lp_equal_tmp_5}},
      PECore_RunFSM_switch_lp_equal_tmp_5});
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_14
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_1 & weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_1 & (~ weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_13
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_1 & weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_1 & (~ weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_12
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_1 & weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_1 & (~ weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_11
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_1 & weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_1 & (~ weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_10
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_1 & weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_1 & (~ weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_9
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_1 & weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_1 & (~ weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_8
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_1 & weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_1 & (~ weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_7
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_1 & weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_1 & (~ weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_6
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_1 & weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_1 & (~ weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_5
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_1 & weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_1 & (~ weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_4
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_1 & weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_1 & (~ weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_3
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_1 & weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_1 & (~ weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_2
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_1 & weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_1 & (~ weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_1
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_1 & weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_1 & (~ weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_0
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_1 & weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_1 & (~ weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_1_nl
      = Arbiter_16U_Roundrobin_pick_priority_29_2_sva_1 & (~ Arbiter_16U_Roundrobin_pick_priority_30_2_sva_1);
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_435_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_2_sva_1) & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_420_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_436_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_2_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_420_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_438_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_2_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_422_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_439_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_2_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_422_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_440_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_2_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_423_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_441_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_2_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_423_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_442_nl
      = (~ operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_424_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_443_nl
      = operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_424_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_444_nl
      = (~ operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_425_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_445_nl
      = operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_425_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_446_nl
      = (~ operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_2_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_426_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_447_nl
      = operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_2_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_426_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_448_nl
      = (~ operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_427_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_449_nl
      = operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_427_cse;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_2_lpi_1_dfm_mx0
      = MUX1HOT_s_1_15_2(Arbiter_16U_Roundrobin_pick_priority_25_2_sva_1, Arbiter_16U_Roundrobin_pick_priority_27_2_sva_1,
      nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_1_nl,
      Arbiter_16U_Roundrobin_pick_priority_17_2_sva_1, Arbiter_16U_Roundrobin_pick_priority_19_2_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_21_2_sva_1, Arbiter_16U_Roundrobin_pick_priority_23_2_sva_1,
      (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[1]), (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[1]),
      (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[1]), (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]),
      (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[1]), (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[1]),
      (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[1]), (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[1]),
      {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_435_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_436_nl
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_2_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_438_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_439_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_440_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_441_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_442_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_443_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_444_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_445_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_446_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_447_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_448_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_449_nl});
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_420_cse
      = (~ operator_3_false_operator_3_false_operator_3_false_or_mdf_2_sva_1) & weight_mem_read_arbxbar_xbar_for_3_2_operator_7_false_operator_7_false_operator_7_false_or_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_422_cse
      = (~ operator_4_false_operator_4_false_operator_4_false_or_mdf_2_sva_1) & and_dcpl_748;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_423_cse
      = operator_4_false_operator_4_false_operator_4_false_or_mdf_2_sva_1 & and_dcpl_748;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_424_cse
      = (~ operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_2_sva_1)
      & and_dcpl_749;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_425_cse
      = operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_2_sva_1 &
      and_dcpl_749;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_426_cse
      = (~ operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_2_sva_1)
      & and_dcpl_756;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_427_cse
      = operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_2_sva_1 &
      and_dcpl_756;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_2_lpi_1_dfm_mx0
      = MUX1HOT_s_1_8_2(operator_2_false_operator_2_false_operator_2_false_or_mdf_2_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_30_2_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_2_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_2_sva_1, operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1,
      operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1, operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_2_sva_1,
      operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1, {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_420_cse
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_2_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_422_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_423_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_424_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_425_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_426_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_427_cse});
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_2_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(operator_3_false_operator_3_false_operator_3_false_or_mdf_2_sva_1,
      operator_4_false_operator_4_false_operator_4_false_or_mdf_2_sva_1, operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_2_sva_1,
      operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_2_sva_1, {weight_mem_read_arbxbar_xbar_for_3_2_operator_7_false_operator_7_false_operator_7_false_or_cse
      , and_dcpl_748 , and_dcpl_749 , and_dcpl_756});
  assign weight_mem_read_arbxbar_xbar_for_3_2_operator_7_false_operator_7_false_operator_7_false_or_cse
      = Arbiter_16U_Roundrobin_pick_priority_30_2_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_2_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_2_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_2_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_2_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_2_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_2_sva_1;
  assign weight_mem_read_arbxbar_xbar_for_3_2_operator_8_false_operator_8_false_operator_8_false_or_nl
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[1]);
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_2_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_2_operator_8_false_operator_8_false_operator_8_false_or_nl,
      weight_mem_read_arbxbar_xbar_for_3_2_operator_7_false_operator_7_false_operator_7_false_or_cse,
      weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign Arbiter_16U_Roundrobin_pick_priority_25_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_10_sva
      & (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[1]);
  assign Arbiter_16U_Roundrobin_pick_priority_27_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_12_sva
      & (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[1]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_2_sva_1 = Arbiter_16U_Roundrobin_pick_priority_27_2_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_2_sva_1;
  assign operator_3_false_operator_3_false_operator_3_false_or_mdf_2_sva_1 = Arbiter_16U_Roundrobin_pick_priority_30_2_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_29_2_sva_1 | Arbiter_16U_Roundrobin_pick_priority_28_2_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_29_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_14_sva
      & (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[1]);
  assign Arbiter_16U_Roundrobin_pick_priority_30_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_15_sva
      & (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[1]);
  assign Arbiter_16U_Roundrobin_pick_priority_26_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_11_sva
      & (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[1]);
  assign Arbiter_16U_Roundrobin_pick_priority_28_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_13_sva
      & (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[1]);
  assign Arbiter_16U_Roundrobin_pick_priority_21_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_6_sva
      & (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[1]);
  assign Arbiter_16U_Roundrobin_pick_priority_23_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_8_sva
      & (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[1]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_2_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_23_2_sva_1 | Arbiter_16U_Roundrobin_pick_priority_22_2_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_17_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_2_sva
      & (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[1]);
  assign Arbiter_16U_Roundrobin_pick_priority_19_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_4_sva
      & (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[1]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_2_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_19_2_sva_1 | Arbiter_16U_Roundrobin_pick_priority_18_2_sva_1;
  assign operator_4_false_operator_4_false_operator_4_false_or_mdf_2_sva_1 = Arbiter_16U_Roundrobin_pick_priority_23_2_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_2_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_2_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_2_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_22_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_7_sva
      & (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[1]);
  assign Arbiter_16U_Roundrobin_pick_priority_18_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_3_sva
      & (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[1]);
  assign Arbiter_16U_Roundrobin_pick_priority_20_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_5_sva
      & (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[1]);
  assign Arbiter_16U_Roundrobin_pick_priority_24_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_9_sva
      & (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[1]);
  assign operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[1]);
  assign operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1
      = (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[1]);
  assign operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_2_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[1]);
  assign operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[1]);
  assign operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_2_sva_1
      = (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[1]);
  assign operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_2_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[1]);
  assign weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp
      = Arbiter_16U_Roundrobin_pick_priority_30_2_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_2_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_2_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_2_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_2_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_2_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_2_sva_1 | Arbiter_16U_Roundrobin_pick_priority_23_2_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_2_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_2_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_2_sva_1 | Arbiter_16U_Roundrobin_pick_priority_19_2_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_18_2_sva_1 | Arbiter_16U_Roundrobin_pick_priority_17_2_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_1_1_sva & (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[1]));
  assign Arbiter_16U_Roundrobin_pick_mux_3009_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_0,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_0,
      weight_mem_read_arbxbar_xbar_for_3_2_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_4_0_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3009_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3008_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_1,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_1,
      weight_mem_read_arbxbar_xbar_for_3_2_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_4_1_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3008_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3006_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_3,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_3,
      weight_mem_read_arbxbar_xbar_for_3_2_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_4_2_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3006_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3002_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_7,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_7,
      weight_mem_read_arbxbar_xbar_for_3_2_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3002_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_14;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_14
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_2 & weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_2 & (~ weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_13
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_2 & weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_2 & (~ weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_12
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_2 & weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_2 & (~ weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_11
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_2 & weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_2 & (~ weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_10
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_2 & weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_2 & (~ weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_9
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_2 & weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_2 & (~ weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_8
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_2 & weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_2 & (~ weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_7
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_2 & weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_2 & (~ weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_6
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_2 & weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_2 & (~ weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_5
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_2 & weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_2 & (~ weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_4
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_2 & weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_2 & (~ weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_3
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_2 & weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_2 & (~ weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_2
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_2 & weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_2 & (~ weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_1
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_2 & weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_2 & (~ weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_0
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_2 & weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_2 & (~ weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_2_nl
      = Arbiter_16U_Roundrobin_pick_priority_29_3_sva_1 & (~ Arbiter_16U_Roundrobin_pick_priority_30_3_sva_1);
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_405_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_3_sva_1) & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_390_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_406_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_3_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_390_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_408_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_3_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_392_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_409_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_3_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_392_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_410_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_3_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_393_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_411_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_3_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_393_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_412_nl
      = (~ operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_394_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_413_nl
      = operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_394_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_414_nl
      = (~ operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_395_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_415_nl
      = operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_395_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_416_nl
      = (~ operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_3_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_396_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_417_nl
      = operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_3_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_396_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_418_nl
      = (~ operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_397_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_419_nl
      = operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_397_cse;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_3_lpi_1_dfm_mx0
      = MUX1HOT_s_1_15_2(Arbiter_16U_Roundrobin_pick_priority_25_3_sva_1, Arbiter_16U_Roundrobin_pick_priority_27_3_sva_1,
      nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_2_nl,
      Arbiter_16U_Roundrobin_pick_priority_17_3_sva_1, Arbiter_16U_Roundrobin_pick_priority_19_3_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_21_3_sva_1, Arbiter_16U_Roundrobin_pick_priority_23_3_sva_1,
      (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[2]), (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[2]),
      (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[2]), (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]),
      (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[2]), (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[2]),
      (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[2]), (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[2]),
      {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_405_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_406_nl
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_3_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_408_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_409_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_410_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_411_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_412_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_413_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_414_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_415_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_416_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_417_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_418_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_419_nl});
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_390_cse
      = (~ operator_3_false_operator_3_false_operator_3_false_or_mdf_3_sva_1) & weight_mem_read_arbxbar_xbar_for_3_3_operator_7_false_operator_7_false_operator_7_false_or_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_392_cse
      = (~ operator_4_false_operator_4_false_operator_4_false_or_mdf_3_sva_1) & and_dcpl_771;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_393_cse
      = operator_4_false_operator_4_false_operator_4_false_or_mdf_3_sva_1 & and_dcpl_771;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_394_cse
      = (~ operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_3_sva_1)
      & and_dcpl_772;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_395_cse
      = operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_3_sva_1 &
      and_dcpl_772;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_396_cse
      = (~ operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_3_sva_1)
      & and_dcpl_779;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_397_cse
      = operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_3_sva_1 &
      and_dcpl_779;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_3_lpi_1_dfm_mx0
      = MUX1HOT_s_1_8_2(operator_2_false_operator_2_false_operator_2_false_or_mdf_3_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_30_3_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_3_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_3_sva_1, operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1,
      operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1, operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_3_sva_1,
      operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1, {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_390_cse
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_3_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_392_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_393_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_394_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_395_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_396_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_397_cse});
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_3_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(operator_3_false_operator_3_false_operator_3_false_or_mdf_3_sva_1,
      operator_4_false_operator_4_false_operator_4_false_or_mdf_3_sva_1, operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_3_sva_1,
      operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_3_sva_1, {weight_mem_read_arbxbar_xbar_for_3_3_operator_7_false_operator_7_false_operator_7_false_or_cse
      , and_dcpl_771 , and_dcpl_772 , and_dcpl_779});
  assign weight_mem_read_arbxbar_xbar_for_3_3_operator_7_false_operator_7_false_operator_7_false_or_cse
      = Arbiter_16U_Roundrobin_pick_priority_30_3_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_3_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_3_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_3_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_3_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_3_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_3_sva_1;
  assign weight_mem_read_arbxbar_xbar_for_3_3_operator_8_false_operator_8_false_operator_8_false_or_nl
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[2]);
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_3_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_3_operator_8_false_operator_8_false_operator_8_false_or_nl,
      weight_mem_read_arbxbar_xbar_for_3_3_operator_7_false_operator_7_false_operator_7_false_or_cse,
      weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign Arbiter_16U_Roundrobin_pick_priority_25_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_10_sva
      & (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[2]);
  assign Arbiter_16U_Roundrobin_pick_priority_27_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_12_sva
      & (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[2]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_3_sva_1 = Arbiter_16U_Roundrobin_pick_priority_27_3_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_3_sva_1;
  assign operator_3_false_operator_3_false_operator_3_false_or_mdf_3_sva_1 = Arbiter_16U_Roundrobin_pick_priority_30_3_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_29_3_sva_1 | Arbiter_16U_Roundrobin_pick_priority_28_3_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_29_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_14_sva
      & (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[2]);
  assign Arbiter_16U_Roundrobin_pick_priority_30_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_15_sva
      & (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[2]);
  assign Arbiter_16U_Roundrobin_pick_priority_26_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_11_sva
      & (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[2]);
  assign Arbiter_16U_Roundrobin_pick_priority_28_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_13_sva
      & (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[2]);
  assign Arbiter_16U_Roundrobin_pick_priority_21_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_6_sva
      & (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[2]);
  assign Arbiter_16U_Roundrobin_pick_priority_23_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_8_sva
      & (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[2]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_3_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_23_3_sva_1 | Arbiter_16U_Roundrobin_pick_priority_22_3_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_17_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_2_sva
      & (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[2]);
  assign Arbiter_16U_Roundrobin_pick_priority_19_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_4_sva
      & (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[2]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_3_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_19_3_sva_1 | Arbiter_16U_Roundrobin_pick_priority_18_3_sva_1;
  assign operator_4_false_operator_4_false_operator_4_false_or_mdf_3_sva_1 = Arbiter_16U_Roundrobin_pick_priority_23_3_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_3_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_3_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_3_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_22_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_7_sva
      & (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[2]);
  assign Arbiter_16U_Roundrobin_pick_priority_18_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_3_sva
      & (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[2]);
  assign Arbiter_16U_Roundrobin_pick_priority_20_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_5_sva
      & (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[2]);
  assign Arbiter_16U_Roundrobin_pick_priority_24_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_9_sva
      & (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[2]);
  assign operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[2]);
  assign operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1
      = (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[2]);
  assign operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_3_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[2]);
  assign operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[2]);
  assign operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_3_sva_1
      = (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[2]);
  assign operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_3_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[2]);
  assign weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp
      = Arbiter_16U_Roundrobin_pick_priority_30_3_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_3_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_3_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_3_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_3_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_3_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_3_sva_1 | Arbiter_16U_Roundrobin_pick_priority_23_3_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_3_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_3_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_3_sva_1 | Arbiter_16U_Roundrobin_pick_priority_19_3_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_18_3_sva_1 | Arbiter_16U_Roundrobin_pick_priority_17_3_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_2_1_sva & (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[2]));
  assign Arbiter_16U_Roundrobin_pick_mux_3023_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_0,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_0,
      weight_mem_read_arbxbar_xbar_for_3_3_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_5_0_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3023_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3022_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_1,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_1,
      weight_mem_read_arbxbar_xbar_for_3_3_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_5_1_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3022_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3020_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_3,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_3,
      weight_mem_read_arbxbar_xbar_for_3_3_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_5_2_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3020_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3016_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_7,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_7,
      weight_mem_read_arbxbar_xbar_for_3_3_operator_31_false_operator_31_false_operator_31_false_or_seb);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3016_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_14;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_14
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_3 & weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_3 & (~ weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_13
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_3 & weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_3 & (~ weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_12
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_3 & weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_3 & (~ weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_11
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_3 & weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_3 & (~ weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_10
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_3 & weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_3 & (~ weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_9
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_3 & weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_3 & (~ weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_8
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_3 & weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_3 & (~ weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_7
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_3 & weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_3 & (~ weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_6
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_3 & weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_3 & (~ weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_5
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_3 & weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_3 & (~ weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_4
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_3 & weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_3 & (~ weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_3
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_3 & weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_3 & (~ weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_2
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_3 & weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_3 & (~ weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_1
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_3 & weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_3 & (~ weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_0
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_3 & weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_3 & (~ weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_3_nl
      = Arbiter_16U_Roundrobin_pick_priority_29_4_sva_1 & (~ Arbiter_16U_Roundrobin_pick_priority_30_4_sva_1);
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_375_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_4_sva_1) & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_360_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_376_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_4_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_360_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_378_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_4_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_362_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_379_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_4_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_362_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_380_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_4_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_363_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_381_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_4_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_363_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_382_nl
      = (~ operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_364_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_383_nl
      = operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_364_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_384_nl
      = (~ operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_365_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_385_nl
      = operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_365_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_386_nl
      = (~ operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_4_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_366_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_387_nl
      = operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_4_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_366_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_388_nl
      = (~ operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_367_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_389_nl
      = operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_367_cse;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_4_lpi_1_dfm_mx0
      = MUX1HOT_s_1_15_2(Arbiter_16U_Roundrobin_pick_priority_25_4_sva_1, Arbiter_16U_Roundrobin_pick_priority_27_4_sva_1,
      nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_3_nl,
      Arbiter_16U_Roundrobin_pick_priority_17_4_sva_1, Arbiter_16U_Roundrobin_pick_priority_19_4_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_21_4_sva_1, Arbiter_16U_Roundrobin_pick_priority_23_4_sva_1,
      (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[3]), (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[3]),
      (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[3]), (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]),
      (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[3]), (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[3]),
      (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[3]), (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[3]),
      {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_375_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_376_nl
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_4_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_378_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_379_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_380_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_381_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_382_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_383_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_384_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_385_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_386_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_387_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_388_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_389_nl});
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_360_cse
      = (~ operator_3_false_operator_3_false_operator_3_false_or_mdf_4_sva_1) & weight_mem_read_arbxbar_xbar_for_3_4_operator_7_false_operator_7_false_operator_7_false_or_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_362_cse
      = (~ operator_4_false_operator_4_false_operator_4_false_or_mdf_4_sva_1) & and_dcpl_794;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_363_cse
      = operator_4_false_operator_4_false_operator_4_false_or_mdf_4_sva_1 & and_dcpl_794;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_364_cse
      = (~ operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_4_sva_1)
      & and_dcpl_795;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_365_cse
      = operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_4_sva_1 &
      and_dcpl_795;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_366_cse
      = (~ operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_4_sva_1)
      & and_dcpl_802;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_367_cse
      = operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_4_sva_1 &
      and_dcpl_802;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_4_lpi_1_dfm_mx0
      = MUX1HOT_s_1_8_2(operator_2_false_operator_2_false_operator_2_false_or_mdf_4_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_30_4_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_4_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_4_sva_1, operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1,
      operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1, operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_4_sva_1,
      operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1, {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_360_cse
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_4_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_362_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_363_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_364_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_365_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_366_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_367_cse});
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_4_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(operator_3_false_operator_3_false_operator_3_false_or_mdf_4_sva_1,
      operator_4_false_operator_4_false_operator_4_false_or_mdf_4_sva_1, operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_4_sva_1,
      operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_4_sva_1, {weight_mem_read_arbxbar_xbar_for_3_4_operator_7_false_operator_7_false_operator_7_false_or_cse
      , and_dcpl_794 , and_dcpl_795 , and_dcpl_802});
  assign weight_mem_read_arbxbar_xbar_for_3_4_operator_7_false_operator_7_false_operator_7_false_or_cse
      = Arbiter_16U_Roundrobin_pick_priority_30_4_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_4_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_4_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_4_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_4_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_4_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_4_sva_1;
  assign weight_mem_read_arbxbar_xbar_for_3_4_operator_8_false_operator_8_false_operator_8_false_or_nl
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[3]);
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_4_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_4_operator_8_false_operator_8_false_operator_8_false_or_nl,
      weight_mem_read_arbxbar_xbar_for_3_4_operator_7_false_operator_7_false_operator_7_false_or_cse,
      weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign Arbiter_16U_Roundrobin_pick_priority_25_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_10_sva
      & (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[3]);
  assign Arbiter_16U_Roundrobin_pick_priority_27_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_12_sva
      & (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[3]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_4_sva_1 = Arbiter_16U_Roundrobin_pick_priority_27_4_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_4_sva_1;
  assign operator_3_false_operator_3_false_operator_3_false_or_mdf_4_sva_1 = Arbiter_16U_Roundrobin_pick_priority_30_4_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_29_4_sva_1 | Arbiter_16U_Roundrobin_pick_priority_28_4_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_29_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_14_sva
      & (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[3]);
  assign Arbiter_16U_Roundrobin_pick_priority_30_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_15_sva
      & (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[3]);
  assign Arbiter_16U_Roundrobin_pick_priority_26_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_11_sva
      & (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[3]);
  assign Arbiter_16U_Roundrobin_pick_priority_28_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_13_sva
      & (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[3]);
  assign Arbiter_16U_Roundrobin_pick_priority_21_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_6_sva
      & (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[3]);
  assign Arbiter_16U_Roundrobin_pick_priority_23_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_8_sva
      & (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[3]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_4_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_23_4_sva_1 | Arbiter_16U_Roundrobin_pick_priority_22_4_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_17_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_2_sva
      & (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[3]);
  assign Arbiter_16U_Roundrobin_pick_priority_19_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_4_sva
      & (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[3]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_4_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_19_4_sva_1 | Arbiter_16U_Roundrobin_pick_priority_18_4_sva_1;
  assign operator_4_false_operator_4_false_operator_4_false_or_mdf_4_sva_1 = Arbiter_16U_Roundrobin_pick_priority_23_4_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_4_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_4_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_4_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_22_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_7_sva
      & (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[3]);
  assign Arbiter_16U_Roundrobin_pick_priority_18_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_3_sva
      & (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[3]);
  assign Arbiter_16U_Roundrobin_pick_priority_20_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_5_sva
      & (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[3]);
  assign Arbiter_16U_Roundrobin_pick_priority_24_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_9_sva
      & (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[3]);
  assign operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[3]);
  assign operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1
      = (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[3]);
  assign operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_4_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[3]);
  assign operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[3]);
  assign operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_4_sva_1
      = (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[3]);
  assign operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_4_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[3]);
  assign weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp
      = Arbiter_16U_Roundrobin_pick_priority_30_4_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_4_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_4_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_4_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_4_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_4_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_4_sva_1 | Arbiter_16U_Roundrobin_pick_priority_23_4_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_4_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_4_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_4_sva_1 | Arbiter_16U_Roundrobin_pick_priority_19_4_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_18_4_sva_1 | Arbiter_16U_Roundrobin_pick_priority_17_4_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_3_1_sva & (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[3]));
  assign Arbiter_16U_Roundrobin_pick_mux_3037_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_0,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_0,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_3_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_6_0_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3037_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3036_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_1,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_1,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_3_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_6_1_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3036_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3034_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_3,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_3,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_3_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_6_2_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3034_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3030_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_7,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_7,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_3_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3030_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_14;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_14
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_4 & weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_4 & (~ weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_13
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_4 & weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_4 & (~ weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_12
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_4 & weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_4 & (~ weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_11
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_4 & weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_4 & (~ weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_10
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_4 & weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_4 & (~ weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_9
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_4 & weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_4 & (~ weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_8
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_4 & weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_4 & (~ weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_7
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_4 & weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_4 & (~ weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_6
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_4 & weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_4 & (~ weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_5
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_4 & weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_4 & (~ weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_4
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_4 & weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_4 & (~ weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_3
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_4 & weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_4 & (~ weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_2
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_4 & weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_4 & (~ weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_1
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_4 & weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_4 & (~ weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_0
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_4 & weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_4 & (~ weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_4_nl
      = Arbiter_16U_Roundrobin_pick_priority_29_5_sva_1 & (~ Arbiter_16U_Roundrobin_pick_priority_30_5_sva_1);
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_345_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_5_sva_1) & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_330_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_346_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_5_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_330_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_348_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_5_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_332_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_349_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_5_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_332_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_350_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_5_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_333_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_351_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_5_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_333_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_352_nl
      = (~ operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_334_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_353_nl
      = operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_334_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_354_nl
      = (~ operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_335_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_355_nl
      = operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_335_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_356_nl
      = (~ operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_5_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_336_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_357_nl
      = operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_5_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_336_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_358_nl
      = (~ operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_337_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_359_nl
      = operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_337_cse;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_5_lpi_1_dfm_mx0
      = MUX1HOT_s_1_15_2(Arbiter_16U_Roundrobin_pick_priority_25_5_sva_1, Arbiter_16U_Roundrobin_pick_priority_27_5_sva_1,
      nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_4_nl,
      Arbiter_16U_Roundrobin_pick_priority_17_5_sva_1, Arbiter_16U_Roundrobin_pick_priority_19_5_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_21_5_sva_1, Arbiter_16U_Roundrobin_pick_priority_23_5_sva_1,
      (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[4]), (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[4]),
      (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[4]), (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]),
      (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[4]), (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[4]),
      (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[4]), (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[4]),
      {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_345_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_346_nl
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_5_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_348_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_349_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_350_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_351_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_352_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_353_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_354_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_355_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_356_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_357_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_358_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_359_nl});
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_330_cse
      = (~ operator_3_false_operator_3_false_operator_3_false_or_mdf_5_sva_1) & weight_mem_read_arbxbar_xbar_for_3_5_operator_7_false_operator_7_false_operator_7_false_or_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_332_cse
      = (~ operator_4_false_operator_4_false_operator_4_false_or_mdf_5_sva_1) & and_dcpl_817;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_333_cse
      = operator_4_false_operator_4_false_operator_4_false_or_mdf_5_sva_1 & and_dcpl_817;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_334_cse
      = (~ operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_5_sva_1)
      & and_dcpl_818;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_335_cse
      = operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_5_sva_1 &
      and_dcpl_818;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_336_cse
      = (~ operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_5_sva_1)
      & and_dcpl_825;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_337_cse
      = operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_5_sva_1 &
      and_dcpl_825;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_5_lpi_1_dfm_mx0
      = MUX1HOT_s_1_8_2(operator_2_false_operator_2_false_operator_2_false_or_mdf_5_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_30_5_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_5_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_5_sva_1, operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1,
      operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1, operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_5_sva_1,
      operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1, {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_330_cse
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_5_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_332_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_333_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_334_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_335_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_336_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_337_cse});
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_5_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(operator_3_false_operator_3_false_operator_3_false_or_mdf_5_sva_1,
      operator_4_false_operator_4_false_operator_4_false_or_mdf_5_sva_1, operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_5_sva_1,
      operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_5_sva_1, {weight_mem_read_arbxbar_xbar_for_3_5_operator_7_false_operator_7_false_operator_7_false_or_cse
      , and_dcpl_817 , and_dcpl_818 , and_dcpl_825});
  assign weight_mem_read_arbxbar_xbar_for_3_5_operator_7_false_operator_7_false_operator_7_false_or_cse
      = Arbiter_16U_Roundrobin_pick_priority_30_5_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_5_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_5_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_5_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_5_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_5_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_5_sva_1;
  assign weight_mem_read_arbxbar_xbar_for_3_5_operator_8_false_operator_8_false_operator_8_false_or_nl
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[4]);
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_5_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_5_operator_8_false_operator_8_false_operator_8_false_or_nl,
      weight_mem_read_arbxbar_xbar_for_3_5_operator_7_false_operator_7_false_operator_7_false_or_cse,
      weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign Arbiter_16U_Roundrobin_pick_priority_25_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_10_sva
      & (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[4]);
  assign Arbiter_16U_Roundrobin_pick_priority_27_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_12_sva
      & (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[4]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_5_sva_1 = Arbiter_16U_Roundrobin_pick_priority_27_5_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_5_sva_1;
  assign operator_3_false_operator_3_false_operator_3_false_or_mdf_5_sva_1 = Arbiter_16U_Roundrobin_pick_priority_30_5_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_29_5_sva_1 | Arbiter_16U_Roundrobin_pick_priority_28_5_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_29_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_14_sva
      & (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[4]);
  assign Arbiter_16U_Roundrobin_pick_priority_30_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_15_sva
      & (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[4]);
  assign Arbiter_16U_Roundrobin_pick_priority_26_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_11_sva
      & (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[4]);
  assign Arbiter_16U_Roundrobin_pick_priority_28_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_13_sva
      & (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[4]);
  assign Arbiter_16U_Roundrobin_pick_priority_21_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_6_sva
      & (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[4]);
  assign Arbiter_16U_Roundrobin_pick_priority_23_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_8_sva
      & (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[4]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_5_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_23_5_sva_1 | Arbiter_16U_Roundrobin_pick_priority_22_5_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_17_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_2_sva
      & (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[4]);
  assign Arbiter_16U_Roundrobin_pick_priority_19_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_4_sva
      & (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[4]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_5_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_19_5_sva_1 | Arbiter_16U_Roundrobin_pick_priority_18_5_sva_1;
  assign operator_4_false_operator_4_false_operator_4_false_or_mdf_5_sva_1 = Arbiter_16U_Roundrobin_pick_priority_23_5_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_5_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_5_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_5_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_22_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_7_sva
      & (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[4]);
  assign Arbiter_16U_Roundrobin_pick_priority_18_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_3_sva
      & (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[4]);
  assign Arbiter_16U_Roundrobin_pick_priority_20_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_5_sva
      & (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[4]);
  assign Arbiter_16U_Roundrobin_pick_priority_24_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_9_sva
      & (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[4]);
  assign operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[4]);
  assign operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1
      = (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[4]);
  assign operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_5_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[4]);
  assign operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[4]);
  assign operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_5_sva_1
      = (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[4]);
  assign operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_5_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[4]);
  assign weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp
      = Arbiter_16U_Roundrobin_pick_priority_30_5_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_5_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_5_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_5_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_5_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_5_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_5_sva_1 | Arbiter_16U_Roundrobin_pick_priority_23_5_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_5_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_5_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_5_sva_1 | Arbiter_16U_Roundrobin_pick_priority_19_5_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_18_5_sva_1 | Arbiter_16U_Roundrobin_pick_priority_17_5_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_4_1_sva & (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[4]));
  assign Arbiter_16U_Roundrobin_pick_mux_3051_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_0,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_0,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_4_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_7_0_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3051_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3050_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_1,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_1,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_4_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_7_1_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3050_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3048_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_3,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_3,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_4_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_7_2_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3048_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3044_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_7,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_7,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_4_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3044_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_14;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_14
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_5 & weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_5 & (~ weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_13
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_5 & weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_5 & (~ weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_12
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_5 & weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_5 & (~ weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_11
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_5 & weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_5 & (~ weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_10
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_5 & weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_5 & (~ weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_9
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_5 & weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_5 & (~ weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_8
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_5 & weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_5 & (~ weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_7
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_5 & weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_5 & (~ weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_6
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_5 & weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_5 & (~ weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_5
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_5 & weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_5 & (~ weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_4
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_5 & weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_5 & (~ weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_3
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_5 & weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_5 & (~ weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_2
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_5 & weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_5 & (~ weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_1
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_5 & weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_5 & (~ weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_0
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_5 & weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_5 & (~ weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_5_nl
      = Arbiter_16U_Roundrobin_pick_priority_29_6_sva_1 & (~ Arbiter_16U_Roundrobin_pick_priority_30_6_sva_1);
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_315_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_6_sva_1) & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_300_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_316_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_6_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_300_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_318_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_6_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_302_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_319_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_6_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_302_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_320_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_6_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_303_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_321_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_6_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_303_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_322_nl
      = (~ operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_304_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_323_nl
      = operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_304_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_324_nl
      = (~ operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_305_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_325_nl
      = operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_305_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_326_nl
      = (~ operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_6_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_306_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_327_nl
      = operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_6_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_306_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_328_nl
      = (~ operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_307_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_329_nl
      = operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_307_cse;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_6_lpi_1_dfm_mx0
      = MUX1HOT_s_1_15_2(Arbiter_16U_Roundrobin_pick_priority_25_6_sva_1, Arbiter_16U_Roundrobin_pick_priority_27_6_sva_1,
      nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_5_nl,
      Arbiter_16U_Roundrobin_pick_priority_17_6_sva_1, Arbiter_16U_Roundrobin_pick_priority_19_6_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_21_6_sva_1, Arbiter_16U_Roundrobin_pick_priority_23_6_sva_1,
      (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[5]), (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[5]),
      (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[5]), (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]),
      (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[5]), (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[5]),
      (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[5]), (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[5]),
      {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_315_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_316_nl
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_6_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_318_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_319_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_320_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_321_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_322_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_323_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_324_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_325_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_326_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_327_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_328_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_329_nl});
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_300_cse
      = (~ operator_3_false_operator_3_false_operator_3_false_or_mdf_6_sva_1) & weight_mem_read_arbxbar_xbar_for_3_6_operator_7_false_operator_7_false_operator_7_false_or_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_302_cse
      = (~ operator_4_false_operator_4_false_operator_4_false_or_mdf_6_sva_1) & and_dcpl_840;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_303_cse
      = operator_4_false_operator_4_false_operator_4_false_or_mdf_6_sva_1 & and_dcpl_840;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_304_cse
      = (~ operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_6_sva_1)
      & and_dcpl_841;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_305_cse
      = operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_6_sva_1 &
      and_dcpl_841;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_306_cse
      = (~ operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_6_sva_1)
      & and_dcpl_848;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_307_cse
      = operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_6_sva_1 &
      and_dcpl_848;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_6_lpi_1_dfm_mx0
      = MUX1HOT_s_1_8_2(operator_2_false_operator_2_false_operator_2_false_or_mdf_6_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_30_6_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_6_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_6_sva_1, operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1,
      operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1, operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_6_sva_1,
      operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1, {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_300_cse
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_6_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_302_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_303_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_304_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_305_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_306_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_307_cse});
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_6_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(operator_3_false_operator_3_false_operator_3_false_or_mdf_6_sva_1,
      operator_4_false_operator_4_false_operator_4_false_or_mdf_6_sva_1, operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_6_sva_1,
      operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_6_sva_1, {weight_mem_read_arbxbar_xbar_for_3_6_operator_7_false_operator_7_false_operator_7_false_or_cse
      , and_dcpl_840 , and_dcpl_841 , and_dcpl_848});
  assign weight_mem_read_arbxbar_xbar_for_3_6_operator_7_false_operator_7_false_operator_7_false_or_cse
      = Arbiter_16U_Roundrobin_pick_priority_30_6_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_6_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_6_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_6_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_6_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_6_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_6_sva_1;
  assign weight_mem_read_arbxbar_xbar_for_3_6_operator_8_false_operator_8_false_operator_8_false_or_nl
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[5]);
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_6_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_6_operator_8_false_operator_8_false_operator_8_false_or_nl,
      weight_mem_read_arbxbar_xbar_for_3_6_operator_7_false_operator_7_false_operator_7_false_or_cse,
      weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign Arbiter_16U_Roundrobin_pick_priority_25_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_10_sva
      & (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[5]);
  assign Arbiter_16U_Roundrobin_pick_priority_27_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_12_sva
      & (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[5]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_6_sva_1 = Arbiter_16U_Roundrobin_pick_priority_27_6_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_6_sva_1;
  assign operator_3_false_operator_3_false_operator_3_false_or_mdf_6_sva_1 = Arbiter_16U_Roundrobin_pick_priority_30_6_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_29_6_sva_1 | Arbiter_16U_Roundrobin_pick_priority_28_6_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_29_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_14_sva
      & (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[5]);
  assign Arbiter_16U_Roundrobin_pick_priority_30_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_15_sva
      & (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[5]);
  assign Arbiter_16U_Roundrobin_pick_priority_26_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_11_sva
      & (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[5]);
  assign Arbiter_16U_Roundrobin_pick_priority_28_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_13_sva
      & (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[5]);
  assign Arbiter_16U_Roundrobin_pick_priority_21_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_6_sva
      & (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[5]);
  assign Arbiter_16U_Roundrobin_pick_priority_23_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_8_sva
      & (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[5]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_6_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_23_6_sva_1 | Arbiter_16U_Roundrobin_pick_priority_22_6_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_17_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_2_sva
      & (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[5]);
  assign Arbiter_16U_Roundrobin_pick_priority_19_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_4_sva
      & (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[5]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_6_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_19_6_sva_1 | Arbiter_16U_Roundrobin_pick_priority_18_6_sva_1;
  assign operator_4_false_operator_4_false_operator_4_false_or_mdf_6_sva_1 = Arbiter_16U_Roundrobin_pick_priority_23_6_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_6_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_6_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_6_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_22_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_7_sva
      & (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[5]);
  assign Arbiter_16U_Roundrobin_pick_priority_18_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_3_sva
      & (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[5]);
  assign Arbiter_16U_Roundrobin_pick_priority_20_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_5_sva
      & (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[5]);
  assign Arbiter_16U_Roundrobin_pick_priority_24_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_9_sva
      & (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[5]);
  assign operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[5]);
  assign operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1
      = (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[5]);
  assign operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_6_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[5]);
  assign operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[5]);
  assign operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_6_sva_1
      = (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[5]);
  assign operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_6_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[5]);
  assign weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp
      = Arbiter_16U_Roundrobin_pick_priority_30_6_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_6_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_6_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_6_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_6_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_6_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_6_sva_1 | Arbiter_16U_Roundrobin_pick_priority_23_6_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_6_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_6_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_6_sva_1 | Arbiter_16U_Roundrobin_pick_priority_19_6_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_18_6_sva_1 | Arbiter_16U_Roundrobin_pick_priority_17_6_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_5_1_sva & (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[5]));
  assign Arbiter_16U_Roundrobin_pick_mux_3065_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_0,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_0,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_5_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_8_0_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3065_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3064_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_1,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_1,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_5_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_8_1_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3064_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3062_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_3,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_3,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_5_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_8_2_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3062_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3058_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_7,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_7,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_5_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3058_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_14;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_14
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_6 & weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_6 & (~ weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_13
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_6 & weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_6 & (~ weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_12
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_6 & weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_6 & (~ weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_11
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_6 & weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_6 & (~ weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_10
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_6 & weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_6 & (~ weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_9
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_6 & weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_6 & (~ weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_8
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_6 & weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_6 & (~ weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_7
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_6 & weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_6 & (~ weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_6
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_6 & weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_6 & (~ weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_5
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_6 & weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_6 & (~ weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_4
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_6 & weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_6 & (~ weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_3
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_6 & weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_6 & (~ weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_2
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_6 & weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_6 & (~ weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_1
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_6 & weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_6 & (~ weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_0
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_6 & weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_6 & (~ weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_6_nl
      = Arbiter_16U_Roundrobin_pick_priority_29_7_sva_1 & (~ Arbiter_16U_Roundrobin_pick_priority_30_7_sva_1);
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_285_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_7_sva_1) & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_270_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_286_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_7_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_270_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_288_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_7_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_272_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_289_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_7_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_272_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_290_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_7_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_273_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_291_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_7_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_273_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_292_nl
      = (~ operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_274_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_293_nl
      = operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_274_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_294_nl
      = (~ operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_275_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_295_nl
      = operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_275_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_296_nl
      = (~ operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_7_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_276_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_297_nl
      = operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_7_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_276_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_298_nl
      = (~ operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_277_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_299_nl
      = operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_277_cse;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_7_lpi_1_dfm_mx0
      = MUX1HOT_s_1_15_2(Arbiter_16U_Roundrobin_pick_priority_25_7_sva_1, Arbiter_16U_Roundrobin_pick_priority_27_7_sva_1,
      nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_6_nl,
      Arbiter_16U_Roundrobin_pick_priority_17_7_sva_1, Arbiter_16U_Roundrobin_pick_priority_19_7_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_21_7_sva_1, Arbiter_16U_Roundrobin_pick_priority_23_7_sva_1,
      (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[6]), (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[6]),
      (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[6]), (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]),
      (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[6]), (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[6]),
      (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[6]), (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[6]),
      {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_285_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_286_nl
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_7_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_288_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_289_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_290_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_291_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_292_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_293_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_294_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_295_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_296_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_297_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_298_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_299_nl});
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_270_cse
      = (~ operator_3_false_operator_3_false_operator_3_false_or_mdf_7_sva_1) & weight_mem_read_arbxbar_xbar_for_3_7_operator_7_false_operator_7_false_operator_7_false_or_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_272_cse
      = (~ operator_4_false_operator_4_false_operator_4_false_or_mdf_7_sva_1) & and_dcpl_863;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_273_cse
      = operator_4_false_operator_4_false_operator_4_false_or_mdf_7_sva_1 & and_dcpl_863;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_274_cse
      = (~ operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_7_sva_1)
      & and_dcpl_864;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_275_cse
      = operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_7_sva_1 &
      and_dcpl_864;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_276_cse
      = (~ operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_7_sva_1)
      & and_dcpl_871;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_277_cse
      = operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_7_sva_1 &
      and_dcpl_871;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_7_lpi_1_dfm_mx0
      = MUX1HOT_s_1_8_2(operator_2_false_operator_2_false_operator_2_false_or_mdf_7_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_30_7_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_7_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_7_sva_1, operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1,
      operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1, operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_7_sva_1,
      operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1, {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_270_cse
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_7_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_272_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_273_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_274_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_275_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_276_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_277_cse});
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_7_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(operator_3_false_operator_3_false_operator_3_false_or_mdf_7_sva_1,
      operator_4_false_operator_4_false_operator_4_false_or_mdf_7_sva_1, operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_7_sva_1,
      operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_7_sva_1, {weight_mem_read_arbxbar_xbar_for_3_7_operator_7_false_operator_7_false_operator_7_false_or_cse
      , and_dcpl_863 , and_dcpl_864 , and_dcpl_871});
  assign weight_mem_read_arbxbar_xbar_for_3_7_operator_7_false_operator_7_false_operator_7_false_or_cse
      = Arbiter_16U_Roundrobin_pick_priority_30_7_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_7_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_7_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_7_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_7_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_7_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_7_sva_1;
  assign weight_mem_read_arbxbar_xbar_for_3_7_operator_8_false_operator_8_false_operator_8_false_or_nl
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[6]);
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_7_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_7_operator_8_false_operator_8_false_operator_8_false_or_nl,
      weight_mem_read_arbxbar_xbar_for_3_7_operator_7_false_operator_7_false_operator_7_false_or_cse,
      weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign Arbiter_16U_Roundrobin_pick_priority_25_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_10_sva
      & (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[6]);
  assign Arbiter_16U_Roundrobin_pick_priority_27_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_12_sva
      & (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[6]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_7_sva_1 = Arbiter_16U_Roundrobin_pick_priority_27_7_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_7_sva_1;
  assign operator_3_false_operator_3_false_operator_3_false_or_mdf_7_sva_1 = Arbiter_16U_Roundrobin_pick_priority_30_7_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_29_7_sva_1 | Arbiter_16U_Roundrobin_pick_priority_28_7_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_29_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_14_sva
      & (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[6]);
  assign Arbiter_16U_Roundrobin_pick_priority_30_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_15_sva
      & (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[6]);
  assign Arbiter_16U_Roundrobin_pick_priority_26_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_11_sva
      & (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[6]);
  assign Arbiter_16U_Roundrobin_pick_priority_28_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_13_sva
      & (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[6]);
  assign Arbiter_16U_Roundrobin_pick_priority_21_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_6_sva
      & (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[6]);
  assign Arbiter_16U_Roundrobin_pick_priority_23_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_8_sva
      & (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[6]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_7_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_23_7_sva_1 | Arbiter_16U_Roundrobin_pick_priority_22_7_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_17_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_2_sva
      & (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[6]);
  assign Arbiter_16U_Roundrobin_pick_priority_19_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_4_sva
      & (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[6]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_7_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_19_7_sva_1 | Arbiter_16U_Roundrobin_pick_priority_18_7_sva_1;
  assign operator_4_false_operator_4_false_operator_4_false_or_mdf_7_sva_1 = Arbiter_16U_Roundrobin_pick_priority_23_7_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_7_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_7_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_7_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_22_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_7_sva
      & (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[6]);
  assign Arbiter_16U_Roundrobin_pick_priority_18_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_3_sva
      & (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[6]);
  assign Arbiter_16U_Roundrobin_pick_priority_20_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_5_sva
      & (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[6]);
  assign Arbiter_16U_Roundrobin_pick_priority_24_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_9_sva
      & (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[6]);
  assign operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[6]);
  assign operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1
      = (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[6]);
  assign operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_7_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[6]);
  assign operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[6]);
  assign operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_7_sva_1
      = (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[6]);
  assign operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_7_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[6]);
  assign weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp
      = Arbiter_16U_Roundrobin_pick_priority_30_7_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_7_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_7_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_7_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_7_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_7_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_7_sva_1 | Arbiter_16U_Roundrobin_pick_priority_23_7_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_7_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_7_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_7_sva_1 | Arbiter_16U_Roundrobin_pick_priority_19_7_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_18_7_sva_1 | Arbiter_16U_Roundrobin_pick_priority_17_7_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_6_1_sva & (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[6]));
  assign Arbiter_16U_Roundrobin_pick_mux_3079_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_0,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_0,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_6_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_9_0_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3079_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3078_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_1,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_1,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_6_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_9_1_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3078_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3076_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_3,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_3,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_6_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_9_2_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3076_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3072_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_7,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_7,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_6_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3072_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_14;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_14
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_7 & weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_7 & (~ weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_13
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_7 & weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_7 & (~ weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_12
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_7 & weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_7 & (~ weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_11
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_7 & weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_7 & (~ weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_10
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_7 & weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_7 & (~ weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_9
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_7 & weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_7 & (~ weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_8
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_7 & weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_7 & (~ weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_7
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_7 & weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_7 & (~ weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_6
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_7 & weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_7 & (~ weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_5
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_7 & weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_7 & (~ weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_4
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_7 & weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_7 & (~ weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_3
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_7 & weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_7 & (~ weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_2
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_7 & weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_7 & (~ weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_1
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_7 & weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_7 & (~ weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_0
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_7 & weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_7 & (~ weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_7_nl
      = Arbiter_16U_Roundrobin_pick_priority_29_8_sva_1 & (~ Arbiter_16U_Roundrobin_pick_priority_30_8_sva_1);
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_255_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_8_sva_1) & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_240_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_256_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_8_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_240_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_258_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_8_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_242_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_259_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_8_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_242_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_260_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_8_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_243_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_261_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_8_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_243_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_262_nl
      = (~ operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_8_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_244_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_263_nl
      = operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_8_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_244_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_264_nl
      = (~ operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_8_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_245_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_265_nl
      = operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_8_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_245_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_266_nl
      = (~ operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_8_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_246_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_267_nl
      = operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_8_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_246_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_268_nl
      = (~ operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_8_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_247_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_269_nl
      = operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_8_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_247_cse;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_8_lpi_1_dfm_mx0
      = MUX1HOT_s_1_15_2(Arbiter_16U_Roundrobin_pick_priority_25_8_sva_1, Arbiter_16U_Roundrobin_pick_priority_27_8_sva_1,
      nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_7_nl,
      Arbiter_16U_Roundrobin_pick_priority_17_8_sva_1, Arbiter_16U_Roundrobin_pick_priority_19_8_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_21_8_sva_1, Arbiter_16U_Roundrobin_pick_priority_23_8_sva_1,
      (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[7]), (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[7]),
      (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[7]), (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]),
      (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[7]), (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[7]),
      (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[7]), (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[7]),
      {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_255_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_256_nl
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_8_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_258_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_259_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_260_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_261_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_262_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_263_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_264_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_265_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_266_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_267_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_268_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_269_nl});
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_240_cse
      = (~ operator_3_false_operator_3_false_operator_3_false_or_mdf_8_sva_1) & weight_mem_read_arbxbar_xbar_for_3_8_operator_7_false_operator_7_false_operator_7_false_or_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_242_cse
      = (~ operator_4_false_operator_4_false_operator_4_false_or_mdf_8_sva_1) & and_dcpl_886;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_243_cse
      = operator_4_false_operator_4_false_operator_4_false_or_mdf_8_sva_1 & and_dcpl_886;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_244_cse
      = (~ operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_8_sva_1)
      & and_dcpl_887;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_245_cse
      = operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_8_sva_1 &
      and_dcpl_887;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_246_cse
      = (~ operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_8_sva_1)
      & and_dcpl_894;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_247_cse
      = operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_8_sva_1 &
      and_dcpl_894;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_8_lpi_1_dfm_mx0
      = MUX1HOT_s_1_8_2(operator_2_false_operator_2_false_operator_2_false_or_mdf_8_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_30_8_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_8_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_8_sva_1, operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_8_sva_1,
      operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_8_sva_1, operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_8_sva_1,
      operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_8_sva_1, {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_240_cse
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_8_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_242_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_243_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_244_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_245_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_246_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_247_cse});
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_8_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(operator_3_false_operator_3_false_operator_3_false_or_mdf_8_sva_1,
      operator_4_false_operator_4_false_operator_4_false_or_mdf_8_sva_1, operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_8_sva_1,
      operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_8_sva_1, {weight_mem_read_arbxbar_xbar_for_3_8_operator_7_false_operator_7_false_operator_7_false_or_cse
      , and_dcpl_886 , and_dcpl_887 , and_dcpl_894});
  assign weight_mem_read_arbxbar_xbar_for_3_8_operator_7_false_operator_7_false_operator_7_false_or_cse
      = Arbiter_16U_Roundrobin_pick_priority_30_8_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_8_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_8_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_8_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_8_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_8_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_8_sva_1;
  assign weight_mem_read_arbxbar_xbar_for_3_8_operator_8_false_operator_8_false_operator_8_false_or_nl
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[7]);
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_8_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_8_operator_8_false_operator_8_false_operator_8_false_or_nl,
      weight_mem_read_arbxbar_xbar_for_3_8_operator_7_false_operator_7_false_operator_7_false_or_cse,
      weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign Arbiter_16U_Roundrobin_pick_priority_25_8_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_10_sva
      & (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[7]);
  assign Arbiter_16U_Roundrobin_pick_priority_27_8_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_12_sva
      & (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[7]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_8_sva_1 = Arbiter_16U_Roundrobin_pick_priority_27_8_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_8_sva_1;
  assign operator_3_false_operator_3_false_operator_3_false_or_mdf_8_sva_1 = Arbiter_16U_Roundrobin_pick_priority_30_8_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_29_8_sva_1 | Arbiter_16U_Roundrobin_pick_priority_28_8_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_29_8_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_14_sva
      & (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[7]);
  assign Arbiter_16U_Roundrobin_pick_priority_30_8_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_15_sva
      & (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[7]);
  assign Arbiter_16U_Roundrobin_pick_priority_26_8_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_11_sva
      & (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[7]);
  assign Arbiter_16U_Roundrobin_pick_priority_28_8_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_13_sva
      & (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[7]);
  assign Arbiter_16U_Roundrobin_pick_priority_21_8_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_6_sva
      & (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[7]);
  assign Arbiter_16U_Roundrobin_pick_priority_23_8_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_8_sva
      & (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[7]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_8_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_23_8_sva_1 | Arbiter_16U_Roundrobin_pick_priority_22_8_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_17_8_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_2_sva
      & (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[7]);
  assign Arbiter_16U_Roundrobin_pick_priority_19_8_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_4_sva
      & (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[7]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_8_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_19_8_sva_1 | Arbiter_16U_Roundrobin_pick_priority_18_8_sva_1;
  assign operator_4_false_operator_4_false_operator_4_false_or_mdf_8_sva_1 = Arbiter_16U_Roundrobin_pick_priority_23_8_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_8_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_8_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_8_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_22_8_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_7_sva
      & (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[7]);
  assign Arbiter_16U_Roundrobin_pick_priority_18_8_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_3_sva
      & (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[7]);
  assign Arbiter_16U_Roundrobin_pick_priority_20_8_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_5_sva
      & (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[7]);
  assign Arbiter_16U_Roundrobin_pick_priority_24_8_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_9_sva
      & (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[7]);
  assign operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_8_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[7]);
  assign operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_8_sva_1
      = (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[7]);
  assign operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_8_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[7]);
  assign operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_8_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[7]);
  assign operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_8_sva_1
      = (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[7]);
  assign operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_8_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[7]);
  assign weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp
      = Arbiter_16U_Roundrobin_pick_priority_30_8_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_8_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_8_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_8_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_8_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_8_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_8_sva_1 | Arbiter_16U_Roundrobin_pick_priority_23_8_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_8_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_8_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_8_sva_1 | Arbiter_16U_Roundrobin_pick_priority_19_8_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_18_8_sva_1 | Arbiter_16U_Roundrobin_pick_priority_17_8_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_7_1_sva & (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[7]));
  assign Arbiter_16U_Roundrobin_pick_mux_3093_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_0,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_0,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_7_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_10_0_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3093_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3092_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_1,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_1,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_7_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_10_1_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3092_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3090_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_3,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_3,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_7_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_10_2_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3090_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3086_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_7,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_7,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_7_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3086_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_14;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_14
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_8 & weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_8 & (~ weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_13
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_8 & weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_8 & (~ weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_12
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_8 & weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_8 & (~ weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_11
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_8 & weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_8 & (~ weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_10
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_8 & weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_8 & (~ weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_9
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_8 & weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_8 & (~ weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_8
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_8 & weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_8 & (~ weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_7
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_8 & weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_8 & (~ weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_6
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_8 & weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_8 & (~ weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_5
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_8 & weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_8 & (~ weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_4
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_8 & weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_8 & (~ weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_3
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_8 & weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_8 & (~ weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_2
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_8 & weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_8 & (~ weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_1
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_8 & weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_8 & (~ weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_0
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_8 & weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_8 & (~ weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_8_nl
      = Arbiter_16U_Roundrobin_pick_priority_29_9_sva_1 & (~ Arbiter_16U_Roundrobin_pick_priority_30_9_sva_1);
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_225_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_9_sva_1) & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_210_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_226_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_9_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_210_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_228_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_9_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_212_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_229_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_9_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_212_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_230_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_9_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_213_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_231_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_9_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_213_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_232_nl
      = (~ operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_9_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_214_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_233_nl
      = operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_9_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_214_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_234_nl
      = (~ operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_9_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_215_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_235_nl
      = operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_9_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_215_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_236_nl
      = (~ operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_9_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_216_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_237_nl
      = operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_9_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_216_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_238_nl
      = (~ operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_9_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_217_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_239_nl
      = operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_9_sva_1 &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_217_cse;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_9_lpi_1_dfm_mx0
      = MUX1HOT_s_1_15_2(Arbiter_16U_Roundrobin_pick_priority_25_9_sva_1, Arbiter_16U_Roundrobin_pick_priority_27_9_sva_1,
      nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_8_nl,
      Arbiter_16U_Roundrobin_pick_priority_17_9_sva_1, Arbiter_16U_Roundrobin_pick_priority_19_9_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_21_9_sva_1, Arbiter_16U_Roundrobin_pick_priority_23_9_sva_1,
      (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[8]), (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[8]),
      (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[8]), (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[8]),
      (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[8]), (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[8]),
      (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[8]), (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[8]),
      {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_225_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_226_nl
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_9_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_228_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_229_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_230_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_231_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_232_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_233_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_234_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_235_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_236_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_237_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_238_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_239_nl});
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_210_cse
      = (~ operator_3_false_operator_3_false_operator_3_false_or_mdf_9_sva_1) & weight_mem_read_arbxbar_xbar_for_3_9_operator_7_false_operator_7_false_operator_7_false_or_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_212_cse
      = (~ operator_4_false_operator_4_false_operator_4_false_or_mdf_9_sva_1) & and_dcpl_909;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_213_cse
      = operator_4_false_operator_4_false_operator_4_false_or_mdf_9_sva_1 & and_dcpl_909;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_214_cse
      = (~ operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_9_sva_1)
      & and_dcpl_910;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_215_cse
      = operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_9_sva_1 &
      and_dcpl_910;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_216_cse
      = (~ operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_9_sva_1)
      & and_dcpl_917;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_217_cse
      = operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_9_sva_1 &
      and_dcpl_917;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_9_lpi_1_dfm_mx0
      = MUX1HOT_s_1_8_2(operator_2_false_operator_2_false_operator_2_false_or_mdf_9_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_30_9_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_9_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_9_sva_1, operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_9_sva_1,
      operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_9_sva_1, operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_9_sva_1,
      operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_9_sva_1, {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_210_cse
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_9_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_212_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_213_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_214_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_215_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_216_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_217_cse});
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_9_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(operator_3_false_operator_3_false_operator_3_false_or_mdf_9_sva_1,
      operator_4_false_operator_4_false_operator_4_false_or_mdf_9_sva_1, operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_9_sva_1,
      operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_9_sva_1, {weight_mem_read_arbxbar_xbar_for_3_9_operator_7_false_operator_7_false_operator_7_false_or_cse
      , and_dcpl_909 , and_dcpl_910 , and_dcpl_917});
  assign weight_mem_read_arbxbar_xbar_for_3_9_operator_7_false_operator_7_false_operator_7_false_or_cse
      = Arbiter_16U_Roundrobin_pick_priority_30_9_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_9_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_9_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_9_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_9_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_9_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_9_sva_1;
  assign weight_mem_read_arbxbar_xbar_for_3_9_operator_8_false_operator_8_false_operator_8_false_or_nl
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[8])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[8])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[8])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[8]);
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_9_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_9_operator_8_false_operator_8_false_operator_8_false_or_nl,
      weight_mem_read_arbxbar_xbar_for_3_9_operator_7_false_operator_7_false_operator_7_false_or_cse,
      weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign Arbiter_16U_Roundrobin_pick_priority_25_9_sva_1 = weight_mem_read_arbxbar_arbiters_next_8_10_sva
      & (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[8]);
  assign Arbiter_16U_Roundrobin_pick_priority_27_9_sva_1 = weight_mem_read_arbxbar_arbiters_next_8_12_sva
      & (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[8]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_9_sva_1 = Arbiter_16U_Roundrobin_pick_priority_27_9_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_9_sva_1;
  assign operator_3_false_operator_3_false_operator_3_false_or_mdf_9_sva_1 = Arbiter_16U_Roundrobin_pick_priority_30_9_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_29_9_sva_1 | Arbiter_16U_Roundrobin_pick_priority_28_9_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_29_9_sva_1 = weight_mem_read_arbxbar_arbiters_next_8_14_sva
      & (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[8]);
  assign Arbiter_16U_Roundrobin_pick_priority_30_9_sva_1 = weight_mem_read_arbxbar_arbiters_next_8_15_sva
      & (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[8]);
  assign Arbiter_16U_Roundrobin_pick_priority_26_9_sva_1 = weight_mem_read_arbxbar_arbiters_next_8_11_sva
      & (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[8]);
  assign Arbiter_16U_Roundrobin_pick_priority_28_9_sva_1 = weight_mem_read_arbxbar_arbiters_next_8_13_sva
      & (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[8]);
  assign Arbiter_16U_Roundrobin_pick_priority_21_9_sva_1 = weight_mem_read_arbxbar_arbiters_next_8_6_sva
      & (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[8]);
  assign Arbiter_16U_Roundrobin_pick_priority_23_9_sva_1 = weight_mem_read_arbxbar_arbiters_next_8_8_sva
      & (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[8]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_9_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_23_9_sva_1 | Arbiter_16U_Roundrobin_pick_priority_22_9_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_17_9_sva_1 = weight_mem_read_arbxbar_arbiters_next_8_2_sva
      & (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[8]);
  assign Arbiter_16U_Roundrobin_pick_priority_19_9_sva_1 = weight_mem_read_arbxbar_arbiters_next_8_4_sva
      & (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[8]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_9_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_19_9_sva_1 | Arbiter_16U_Roundrobin_pick_priority_18_9_sva_1;
  assign operator_4_false_operator_4_false_operator_4_false_or_mdf_9_sva_1 = Arbiter_16U_Roundrobin_pick_priority_23_9_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_9_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_9_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_9_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_22_9_sva_1 = weight_mem_read_arbxbar_arbiters_next_8_7_sva
      & (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[8]);
  assign Arbiter_16U_Roundrobin_pick_priority_18_9_sva_1 = weight_mem_read_arbxbar_arbiters_next_8_3_sva
      & (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[8]);
  assign Arbiter_16U_Roundrobin_pick_priority_20_9_sva_1 = weight_mem_read_arbxbar_arbiters_next_8_5_sva
      & (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[8]);
  assign Arbiter_16U_Roundrobin_pick_priority_24_9_sva_1 = weight_mem_read_arbxbar_arbiters_next_8_9_sva
      & (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[8]);
  assign operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_9_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[8]);
  assign operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_9_sva_1
      = (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[8]);
  assign operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_9_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[8])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[8]);
  assign operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_9_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[8]);
  assign operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_9_sva_1
      = (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[8]);
  assign operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_9_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[8])
      | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[8]);
  assign weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp
      = Arbiter_16U_Roundrobin_pick_priority_30_9_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_9_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_9_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_9_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_9_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_9_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_9_sva_1 | Arbiter_16U_Roundrobin_pick_priority_23_9_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_9_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_9_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_9_sva_1 | Arbiter_16U_Roundrobin_pick_priority_19_9_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_18_9_sva_1 | Arbiter_16U_Roundrobin_pick_priority_17_9_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_8_1_sva & (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[8]));
  assign Arbiter_16U_Roundrobin_pick_mux_3107_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_0,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_0,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_8_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_11_0_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3107_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3106_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_1,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_1,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_8_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_11_1_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3106_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3104_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_3,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_3,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_8_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_11_2_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3104_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3100_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_7,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_7,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_8_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3100_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_14;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_14
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_9 & weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_9 & (~ weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_13
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_9 & weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_9 & (~ weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_12
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_9 & weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_9 & (~ weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_11
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_9 & weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_9 & (~ weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_10
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_9 & weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_9 & (~ weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_9
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_9 & weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_9 & (~ weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_8
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_9 & weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_9 & (~ weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_7
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_9 & weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_9 & (~ weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_6
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_9 & weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_9 & (~ weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_5
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_9 & weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_9 & (~ weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_4
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_9 & weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_9 & (~ weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_3
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_9 & weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_9 & (~ weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_2
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_9 & weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_9 & (~ weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_1
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_9 & weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_9 & (~ weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_0
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_9 & weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_9 & (~ weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_9_nl
      = Arbiter_16U_Roundrobin_pick_priority_29_10_sva_1 & (~ Arbiter_16U_Roundrobin_pick_priority_30_10_sva_1);
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_195_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_10_sva_1) &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_180_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_196_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_10_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_180_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_198_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_10_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_182_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_199_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_10_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_182_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_200_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_10_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_183_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_201_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_10_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_183_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_202_nl
      = (~ operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_10_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_184_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_203_nl
      = operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_10_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_184_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_204_nl
      = (~ operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_10_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_185_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_205_nl
      = operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_10_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_185_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_206_nl
      = (~ operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_10_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_186_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_207_nl
      = operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_10_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_186_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_208_nl
      = (~ operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_10_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_187_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_209_nl
      = operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_10_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_187_cse;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_10_lpi_1_dfm_mx0
      = MUX1HOT_s_1_15_2(Arbiter_16U_Roundrobin_pick_priority_25_10_sva_1, Arbiter_16U_Roundrobin_pick_priority_27_10_sva_1,
      nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_9_nl,
      Arbiter_16U_Roundrobin_pick_priority_17_10_sva_1, Arbiter_16U_Roundrobin_pick_priority_19_10_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_21_10_sva_1, Arbiter_16U_Roundrobin_pick_priority_23_10_sva_1,
      (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[9]), (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[9]),
      (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[9]), (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[9]),
      (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[9]), (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[9]),
      (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[9]), (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[9]),
      {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_195_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_196_nl
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_10_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_198_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_199_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_200_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_201_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_202_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_203_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_204_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_205_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_206_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_207_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_208_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_209_nl});
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_180_cse
      = (~ operator_3_false_operator_3_false_operator_3_false_or_mdf_10_sva_1) &
      weight_mem_read_arbxbar_xbar_for_3_10_operator_7_false_operator_7_false_operator_7_false_or_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_182_cse
      = (~ operator_4_false_operator_4_false_operator_4_false_or_mdf_10_sva_1) &
      and_dcpl_932;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_183_cse
      = operator_4_false_operator_4_false_operator_4_false_or_mdf_10_sva_1 & and_dcpl_932;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_184_cse
      = (~ operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_10_sva_1)
      & and_dcpl_933;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_185_cse
      = operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_10_sva_1
      & and_dcpl_933;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_186_cse
      = (~ operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_10_sva_1)
      & and_dcpl_939;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_187_cse
      = operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_10_sva_1
      & and_dcpl_939;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_10_lpi_1_dfm_mx0
      = MUX1HOT_s_1_8_2(operator_2_false_operator_2_false_operator_2_false_or_mdf_10_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_30_10_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_10_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_10_sva_1, operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_10_sva_1,
      operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_10_sva_1, operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_10_sva_1,
      operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_10_sva_1, {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_180_cse
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_10_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_182_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_183_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_184_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_185_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_186_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_187_cse});
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_10_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(operator_3_false_operator_3_false_operator_3_false_or_mdf_10_sva_1,
      operator_4_false_operator_4_false_operator_4_false_or_mdf_10_sva_1, operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_10_sva_1,
      operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_10_sva_1, {weight_mem_read_arbxbar_xbar_for_3_10_operator_7_false_operator_7_false_operator_7_false_or_cse
      , and_dcpl_932 , and_dcpl_933 , and_dcpl_939});
  assign weight_mem_read_arbxbar_xbar_for_3_10_operator_7_false_operator_7_false_operator_7_false_or_cse
      = Arbiter_16U_Roundrobin_pick_priority_30_10_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_10_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_10_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_10_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_10_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_10_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_10_sva_1;
  assign weight_mem_read_arbxbar_xbar_for_3_10_operator_8_false_operator_8_false_operator_8_false_or_nl
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[9])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[9])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[9])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[9]);
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_10_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_10_operator_8_false_operator_8_false_operator_8_false_or_nl,
      weight_mem_read_arbxbar_xbar_for_3_10_operator_7_false_operator_7_false_operator_7_false_or_cse,
      weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign Arbiter_16U_Roundrobin_pick_priority_25_10_sva_1 = weight_mem_read_arbxbar_arbiters_next_9_10_sva
      & (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[9]);
  assign Arbiter_16U_Roundrobin_pick_priority_27_10_sva_1 = weight_mem_read_arbxbar_arbiters_next_9_12_sva
      & (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[9]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_10_sva_1 = Arbiter_16U_Roundrobin_pick_priority_27_10_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_10_sva_1;
  assign operator_3_false_operator_3_false_operator_3_false_or_mdf_10_sva_1 = Arbiter_16U_Roundrobin_pick_priority_30_10_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_29_10_sva_1 | Arbiter_16U_Roundrobin_pick_priority_28_10_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_29_10_sva_1 = weight_mem_read_arbxbar_arbiters_next_9_14_sva
      & (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[9]);
  assign Arbiter_16U_Roundrobin_pick_priority_30_10_sva_1 = weight_mem_read_arbxbar_arbiters_next_9_15_sva
      & (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[9]);
  assign Arbiter_16U_Roundrobin_pick_priority_26_10_sva_1 = weight_mem_read_arbxbar_arbiters_next_9_11_sva
      & (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[9]);
  assign Arbiter_16U_Roundrobin_pick_priority_28_10_sva_1 = weight_mem_read_arbxbar_arbiters_next_9_13_sva
      & (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[9]);
  assign Arbiter_16U_Roundrobin_pick_priority_21_10_sva_1 = weight_mem_read_arbxbar_arbiters_next_9_6_sva
      & (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[9]);
  assign Arbiter_16U_Roundrobin_pick_priority_23_10_sva_1 = weight_mem_read_arbxbar_arbiters_next_9_8_sva
      & (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[9]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_10_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_23_10_sva_1 | Arbiter_16U_Roundrobin_pick_priority_22_10_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_17_10_sva_1 = weight_mem_read_arbxbar_arbiters_next_9_2_sva
      & (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[9]);
  assign Arbiter_16U_Roundrobin_pick_priority_19_10_sva_1 = weight_mem_read_arbxbar_arbiters_next_9_4_sva
      & (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[9]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_10_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_19_10_sva_1 | Arbiter_16U_Roundrobin_pick_priority_18_10_sva_1;
  assign operator_4_false_operator_4_false_operator_4_false_or_mdf_10_sva_1 = Arbiter_16U_Roundrobin_pick_priority_23_10_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_10_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_10_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_10_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_22_10_sva_1 = weight_mem_read_arbxbar_arbiters_next_9_7_sva
      & (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[9]);
  assign Arbiter_16U_Roundrobin_pick_priority_18_10_sva_1 = weight_mem_read_arbxbar_arbiters_next_9_3_sva
      & (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[9]);
  assign Arbiter_16U_Roundrobin_pick_priority_20_10_sva_1 = weight_mem_read_arbxbar_arbiters_next_9_5_sva
      & (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[9]);
  assign Arbiter_16U_Roundrobin_pick_priority_24_10_sva_1 = weight_mem_read_arbxbar_arbiters_next_9_9_sva
      & (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[9]);
  assign operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_10_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[9]);
  assign operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_10_sva_1
      = (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[9]);
  assign operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_10_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[9])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[9]);
  assign operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_10_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[9]);
  assign operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_10_sva_1
      = (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[9]);
  assign operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_10_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[9])
      | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[9]);
  assign weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp
      = Arbiter_16U_Roundrobin_pick_priority_30_10_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_10_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_10_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_10_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_10_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_10_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_10_sva_1 | Arbiter_16U_Roundrobin_pick_priority_23_10_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_10_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_10_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_10_sva_1 | Arbiter_16U_Roundrobin_pick_priority_19_10_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_18_10_sva_1 | Arbiter_16U_Roundrobin_pick_priority_17_10_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_9_1_sva & (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[9]));
  assign Arbiter_16U_Roundrobin_pick_mux_3121_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_0,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_0,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_9_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_12_0_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3121_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3120_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_1,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_1,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_9_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_12_1_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3120_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3118_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_3,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_3,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_9_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_12_2_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3118_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3114_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_7,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_7,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_9_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3114_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_14;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_14
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_10 & weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_10 & (~ weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_13
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_10 & weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_10 & (~ weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_12
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_10 & weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_10 & (~ weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_11
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_10 & weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_10 & (~ weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_10
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_10 & weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_10 & (~ weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_9
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_10 & weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_10 & (~ weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_8
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_10 & weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_10 & (~ weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_7
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_10 & weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_10 & (~ weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_6
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_10 & weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_10 & (~ weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_5
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_10 & weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_10 & (~ weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_4
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_10 & weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_10 & (~ weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_3
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_10 & weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_10 & (~ weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_2
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_10 & weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_10 & (~ weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_1
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_10 & weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_10 & (~ weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_0
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_10 & weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_10 & (~ weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_10_nl
      = Arbiter_16U_Roundrobin_pick_priority_29_11_sva_1 & (~ Arbiter_16U_Roundrobin_pick_priority_30_11_sva_1);
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_165_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_11_sva_1) &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_150_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_166_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_11_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_150_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_168_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_11_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_152_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_169_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_11_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_152_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_170_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_11_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_153_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_171_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_11_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_153_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_172_nl
      = (~ operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_11_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_154_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_173_nl
      = operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_11_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_154_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_174_nl
      = (~ operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_11_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_155_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_175_nl
      = operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_11_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_155_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_176_nl
      = (~ operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_11_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_156_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_177_nl
      = operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_11_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_156_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_178_nl
      = (~ operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_11_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_157_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_179_nl
      = operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_11_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_157_cse;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_11_lpi_1_dfm_mx0
      = MUX1HOT_s_1_15_2(Arbiter_16U_Roundrobin_pick_priority_25_11_sva_1, Arbiter_16U_Roundrobin_pick_priority_27_11_sva_1,
      nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_10_nl,
      Arbiter_16U_Roundrobin_pick_priority_17_11_sva_1, Arbiter_16U_Roundrobin_pick_priority_19_11_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_21_11_sva_1, Arbiter_16U_Roundrobin_pick_priority_23_11_sva_1,
      (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[10]), (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[10]),
      (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[10]), (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[10]),
      (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[10]), (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[10]),
      (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[10]), (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[10]),
      {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_165_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_166_nl
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_11_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_168_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_169_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_170_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_171_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_172_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_173_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_174_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_175_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_176_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_177_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_178_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_179_nl});
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_150_cse
      = (~ operator_3_false_operator_3_false_operator_3_false_or_mdf_11_sva_1) &
      weight_mem_read_arbxbar_xbar_for_3_11_operator_7_false_operator_7_false_operator_7_false_or_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_152_cse
      = (~ operator_4_false_operator_4_false_operator_4_false_or_mdf_11_sva_1) &
      and_dcpl_954;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_153_cse
      = operator_4_false_operator_4_false_operator_4_false_or_mdf_11_sva_1 & and_dcpl_954;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_154_cse
      = (~ operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_11_sva_1)
      & and_dcpl_955;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_155_cse
      = operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_11_sva_1
      & and_dcpl_955;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_156_cse
      = (~ operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_11_sva_1)
      & and_dcpl_962;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_157_cse
      = operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_11_sva_1
      & and_dcpl_962;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_11_lpi_1_dfm_mx0
      = MUX1HOT_s_1_8_2(operator_2_false_operator_2_false_operator_2_false_or_mdf_11_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_30_11_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_11_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_11_sva_1, operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_11_sva_1,
      operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_11_sva_1, operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_11_sva_1,
      operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_11_sva_1, {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_150_cse
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_11_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_152_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_153_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_154_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_155_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_156_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_157_cse});
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_11_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(operator_3_false_operator_3_false_operator_3_false_or_mdf_11_sva_1,
      operator_4_false_operator_4_false_operator_4_false_or_mdf_11_sva_1, operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_11_sva_1,
      operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_11_sva_1, {weight_mem_read_arbxbar_xbar_for_3_11_operator_7_false_operator_7_false_operator_7_false_or_cse
      , and_dcpl_954 , and_dcpl_955 , and_dcpl_962});
  assign weight_mem_read_arbxbar_xbar_for_3_11_operator_7_false_operator_7_false_operator_7_false_or_cse
      = Arbiter_16U_Roundrobin_pick_priority_30_11_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_11_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_11_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_11_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_11_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_11_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_11_sva_1;
  assign weight_mem_read_arbxbar_xbar_for_3_11_operator_8_false_operator_8_false_operator_8_false_or_nl
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[10])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[10])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[10])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[10]);
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_11_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_11_operator_8_false_operator_8_false_operator_8_false_or_nl,
      weight_mem_read_arbxbar_xbar_for_3_11_operator_7_false_operator_7_false_operator_7_false_or_cse,
      weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign Arbiter_16U_Roundrobin_pick_priority_25_11_sva_1 = weight_mem_read_arbxbar_arbiters_next_10_10_sva
      & (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[10]);
  assign Arbiter_16U_Roundrobin_pick_priority_27_11_sva_1 = weight_mem_read_arbxbar_arbiters_next_10_12_sva
      & (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[10]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_11_sva_1 = Arbiter_16U_Roundrobin_pick_priority_27_11_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_11_sva_1;
  assign operator_3_false_operator_3_false_operator_3_false_or_mdf_11_sva_1 = Arbiter_16U_Roundrobin_pick_priority_30_11_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_29_11_sva_1 | Arbiter_16U_Roundrobin_pick_priority_28_11_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_29_11_sva_1 = weight_mem_read_arbxbar_arbiters_next_10_14_sva
      & (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[10]);
  assign Arbiter_16U_Roundrobin_pick_priority_30_11_sva_1 = weight_mem_read_arbxbar_arbiters_next_10_15_sva
      & (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[10]);
  assign Arbiter_16U_Roundrobin_pick_priority_26_11_sva_1 = weight_mem_read_arbxbar_arbiters_next_10_11_sva
      & (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[10]);
  assign Arbiter_16U_Roundrobin_pick_priority_28_11_sva_1 = weight_mem_read_arbxbar_arbiters_next_10_13_sva
      & (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[10]);
  assign Arbiter_16U_Roundrobin_pick_priority_21_11_sva_1 = weight_mem_read_arbxbar_arbiters_next_10_6_sva
      & (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[10]);
  assign Arbiter_16U_Roundrobin_pick_priority_23_11_sva_1 = weight_mem_read_arbxbar_arbiters_next_10_8_sva
      & (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[10]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_11_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_23_11_sva_1 | Arbiter_16U_Roundrobin_pick_priority_22_11_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_17_11_sva_1 = weight_mem_read_arbxbar_arbiters_next_10_2_sva
      & (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[10]);
  assign Arbiter_16U_Roundrobin_pick_priority_19_11_sva_1 = weight_mem_read_arbxbar_arbiters_next_10_4_sva
      & (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[10]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_11_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_19_11_sva_1 | Arbiter_16U_Roundrobin_pick_priority_18_11_sva_1;
  assign operator_4_false_operator_4_false_operator_4_false_or_mdf_11_sva_1 = Arbiter_16U_Roundrobin_pick_priority_23_11_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_11_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_11_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_11_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_22_11_sva_1 = weight_mem_read_arbxbar_arbiters_next_10_7_sva
      & (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[10]);
  assign Arbiter_16U_Roundrobin_pick_priority_18_11_sva_1 = weight_mem_read_arbxbar_arbiters_next_10_3_sva
      & (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[10]);
  assign Arbiter_16U_Roundrobin_pick_priority_20_11_sva_1 = weight_mem_read_arbxbar_arbiters_next_10_5_sva
      & (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[10]);
  assign Arbiter_16U_Roundrobin_pick_priority_24_11_sva_1 = weight_mem_read_arbxbar_arbiters_next_10_9_sva
      & (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[10]);
  assign operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_11_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[10]);
  assign operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_11_sva_1
      = (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[10]);
  assign operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_11_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[10])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[10]);
  assign operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_11_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[10]);
  assign operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_11_sva_1
      = (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[10]);
  assign operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_11_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[10])
      | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[10]);
  assign weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp
      = Arbiter_16U_Roundrobin_pick_priority_30_11_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_11_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_11_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_11_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_11_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_11_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_11_sva_1 | Arbiter_16U_Roundrobin_pick_priority_23_11_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_11_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_11_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_11_sva_1 | Arbiter_16U_Roundrobin_pick_priority_19_11_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_18_11_sva_1 | Arbiter_16U_Roundrobin_pick_priority_17_11_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_10_1_sva & (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[10]));
  assign Arbiter_16U_Roundrobin_pick_mux_3135_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_0,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_0,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_10_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_13_0_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3135_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3134_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_1,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_1,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_10_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_13_1_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3134_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3132_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_3,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_3,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_10_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_13_2_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3132_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3128_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_7,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_7,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_10_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3128_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_14;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_14
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_11 & weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_11 & (~ weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_13
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_11 & weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_11 & (~ weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_12
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_11 & weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_11 & (~ weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_11
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_11 & weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_11 & (~ weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_10
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_11 & weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_11 & (~ weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_9
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_11 & weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_11 & (~ weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_8
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_11 & weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_11 & (~ weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_7
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_11 & weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_11 & (~ weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_6
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_11 & weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_11 & (~ weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_5
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_11 & weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_11 & (~ weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_4
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_11 & weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_11 & (~ weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_3
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_11 & weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_11 & (~ weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_2
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_11 & weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_11 & (~ weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_1
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_11 & weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_11 & (~ weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_0
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_11 & weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_11 & (~ weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_11_nl
      = Arbiter_16U_Roundrobin_pick_priority_29_12_sva_1 & (~ Arbiter_16U_Roundrobin_pick_priority_30_12_sva_1);
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_135_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_12_sva_1) &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_120_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_136_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_12_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_120_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_138_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_12_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_122_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_139_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_12_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_122_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_140_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_12_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_123_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_141_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_12_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_123_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_142_nl
      = (~ operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_12_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_124_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_143_nl
      = operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_12_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_124_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_144_nl
      = (~ operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_12_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_125_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_145_nl
      = operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_12_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_125_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_146_nl
      = (~ operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_12_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_126_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_147_nl
      = operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_12_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_126_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_148_nl
      = (~ operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_12_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_127_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_149_nl
      = operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_12_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_127_cse;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_12_lpi_1_dfm_mx0
      = MUX1HOT_s_1_15_2(Arbiter_16U_Roundrobin_pick_priority_25_12_sva_1, Arbiter_16U_Roundrobin_pick_priority_27_12_sva_1,
      nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_11_nl,
      Arbiter_16U_Roundrobin_pick_priority_17_12_sva_1, Arbiter_16U_Roundrobin_pick_priority_19_12_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_21_12_sva_1, Arbiter_16U_Roundrobin_pick_priority_23_12_sva_1,
      (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[11]), (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[11]),
      (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[11]), (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[11]),
      (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[11]), (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[11]),
      (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[11]), (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[11]),
      {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_135_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_136_nl
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_12_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_138_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_139_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_140_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_141_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_142_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_143_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_144_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_145_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_146_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_147_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_148_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_149_nl});
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_120_cse
      = (~ operator_3_false_operator_3_false_operator_3_false_or_mdf_12_sva_1) &
      weight_mem_read_arbxbar_xbar_for_3_12_operator_7_false_operator_7_false_operator_7_false_or_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_122_cse
      = (~ operator_4_false_operator_4_false_operator_4_false_or_mdf_12_sva_1) &
      and_dcpl_977;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_123_cse
      = operator_4_false_operator_4_false_operator_4_false_or_mdf_12_sva_1 & and_dcpl_977;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_124_cse
      = (~ operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_12_sva_1)
      & and_dcpl_978;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_125_cse
      = operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_12_sva_1
      & and_dcpl_978;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_126_cse
      = (~ operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_12_sva_1)
      & and_dcpl_985;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_127_cse
      = operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_12_sva_1
      & and_dcpl_985;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_12_lpi_1_dfm_mx0
      = MUX1HOT_s_1_8_2(operator_2_false_operator_2_false_operator_2_false_or_mdf_12_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_30_12_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_12_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_12_sva_1, operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_12_sva_1,
      operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_12_sva_1, operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_12_sva_1,
      operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_12_sva_1, {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_120_cse
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_12_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_122_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_123_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_124_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_125_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_126_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_127_cse});
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_12_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(operator_3_false_operator_3_false_operator_3_false_or_mdf_12_sva_1,
      operator_4_false_operator_4_false_operator_4_false_or_mdf_12_sva_1, operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_12_sva_1,
      operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_12_sva_1, {weight_mem_read_arbxbar_xbar_for_3_12_operator_7_false_operator_7_false_operator_7_false_or_cse
      , and_dcpl_977 , and_dcpl_978 , and_dcpl_985});
  assign weight_mem_read_arbxbar_xbar_for_3_12_operator_7_false_operator_7_false_operator_7_false_or_cse
      = Arbiter_16U_Roundrobin_pick_priority_30_12_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_12_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_12_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_12_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_12_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_12_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_12_sva_1;
  assign weight_mem_read_arbxbar_xbar_for_3_12_operator_8_false_operator_8_false_operator_8_false_or_nl
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[11])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[11])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[11])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[11]);
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_12_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_12_operator_8_false_operator_8_false_operator_8_false_or_nl,
      weight_mem_read_arbxbar_xbar_for_3_12_operator_7_false_operator_7_false_operator_7_false_or_cse,
      weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign Arbiter_16U_Roundrobin_pick_priority_25_12_sva_1 = weight_mem_read_arbxbar_arbiters_next_11_10_sva
      & (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[11]);
  assign Arbiter_16U_Roundrobin_pick_priority_27_12_sva_1 = weight_mem_read_arbxbar_arbiters_next_11_12_sva
      & (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[11]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_12_sva_1 = Arbiter_16U_Roundrobin_pick_priority_27_12_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_12_sva_1;
  assign operator_3_false_operator_3_false_operator_3_false_or_mdf_12_sva_1 = Arbiter_16U_Roundrobin_pick_priority_30_12_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_29_12_sva_1 | Arbiter_16U_Roundrobin_pick_priority_28_12_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_29_12_sva_1 = weight_mem_read_arbxbar_arbiters_next_11_14_sva
      & (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[11]);
  assign Arbiter_16U_Roundrobin_pick_priority_30_12_sva_1 = weight_mem_read_arbxbar_arbiters_next_11_15_sva
      & (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[11]);
  assign Arbiter_16U_Roundrobin_pick_priority_26_12_sva_1 = weight_mem_read_arbxbar_arbiters_next_11_11_sva
      & (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[11]);
  assign Arbiter_16U_Roundrobin_pick_priority_28_12_sva_1 = weight_mem_read_arbxbar_arbiters_next_11_13_sva
      & (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[11]);
  assign Arbiter_16U_Roundrobin_pick_priority_21_12_sva_1 = weight_mem_read_arbxbar_arbiters_next_11_6_sva
      & (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[11]);
  assign Arbiter_16U_Roundrobin_pick_priority_23_12_sva_1 = weight_mem_read_arbxbar_arbiters_next_11_8_sva
      & (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[11]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_12_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_23_12_sva_1 | Arbiter_16U_Roundrobin_pick_priority_22_12_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_17_12_sva_1 = weight_mem_read_arbxbar_arbiters_next_11_2_sva
      & (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[11]);
  assign Arbiter_16U_Roundrobin_pick_priority_19_12_sva_1 = weight_mem_read_arbxbar_arbiters_next_11_4_sva
      & (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[11]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_12_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_19_12_sva_1 | Arbiter_16U_Roundrobin_pick_priority_18_12_sva_1;
  assign operator_4_false_operator_4_false_operator_4_false_or_mdf_12_sva_1 = Arbiter_16U_Roundrobin_pick_priority_23_12_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_12_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_12_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_12_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_22_12_sva_1 = weight_mem_read_arbxbar_arbiters_next_11_7_sva
      & (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[11]);
  assign Arbiter_16U_Roundrobin_pick_priority_18_12_sva_1 = weight_mem_read_arbxbar_arbiters_next_11_3_sva
      & (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[11]);
  assign Arbiter_16U_Roundrobin_pick_priority_20_12_sva_1 = weight_mem_read_arbxbar_arbiters_next_11_5_sva
      & (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[11]);
  assign Arbiter_16U_Roundrobin_pick_priority_24_12_sva_1 = weight_mem_read_arbxbar_arbiters_next_11_9_sva
      & (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[11]);
  assign operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_12_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[11]);
  assign operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_12_sva_1
      = (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[11]);
  assign operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_12_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[11])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[11]);
  assign operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_12_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[11]);
  assign operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_12_sva_1
      = (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[11]);
  assign operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_12_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[11])
      | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[11]);
  assign weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp
      = Arbiter_16U_Roundrobin_pick_priority_30_12_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_12_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_12_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_12_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_12_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_12_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_12_sva_1 | Arbiter_16U_Roundrobin_pick_priority_23_12_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_12_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_12_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_12_sva_1 | Arbiter_16U_Roundrobin_pick_priority_19_12_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_18_12_sva_1 | Arbiter_16U_Roundrobin_pick_priority_17_12_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_11_1_sva & (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[11]));
  assign Arbiter_16U_Roundrobin_pick_mux_3149_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_0,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_0,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_11_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_14_0_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3149_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3148_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_1,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_1,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_11_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_14_1_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3148_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3146_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_3,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_3,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_11_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_14_2_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3146_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3142_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_7,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_7,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_11_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3142_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_14;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_14
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_12 & weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_12 & (~ weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_13
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_12 & weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_12 & (~ weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_12
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_12 & weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_12 & (~ weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_11
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_12 & weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_12 & (~ weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_10
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_12 & weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_12 & (~ weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_9
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_12 & weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_12 & (~ weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_8
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_12 & weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_12 & (~ weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_7
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_12 & weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_12 & (~ weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_6
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_12 & weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_12 & (~ weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_5
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_12 & weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_12 & (~ weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_4
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_12 & weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_12 & (~ weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_3
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_12 & weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_12 & (~ weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_2
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_12 & weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_12 & (~ weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_1
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_12 & weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_12 & (~ weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_0
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_12 & weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_12 & (~ weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_12_nl
      = Arbiter_16U_Roundrobin_pick_priority_29_13_sva_1 & (~ Arbiter_16U_Roundrobin_pick_priority_30_13_sva_1);
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_105_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_13_sva_1) &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_90_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_106_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_13_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_90_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_108_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_13_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_92_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_109_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_13_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_92_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_110_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_13_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_93_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_111_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_13_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_93_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_112_nl
      = (~ operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_13_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_94_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_113_nl
      = operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_13_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_94_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_114_nl
      = (~ operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_13_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_95_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_115_nl
      = operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_13_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_95_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_116_nl
      = (~ operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_13_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_96_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_117_nl
      = operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_13_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_96_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_118_nl
      = (~ operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_13_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_97_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_119_nl
      = operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_13_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_97_cse;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_13_lpi_1_dfm_mx0
      = MUX1HOT_s_1_15_2(Arbiter_16U_Roundrobin_pick_priority_25_13_sva_1, Arbiter_16U_Roundrobin_pick_priority_27_13_sva_1,
      nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_12_nl,
      Arbiter_16U_Roundrobin_pick_priority_17_13_sva_1, Arbiter_16U_Roundrobin_pick_priority_19_13_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_21_13_sva_1, Arbiter_16U_Roundrobin_pick_priority_23_13_sva_1,
      (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[12]), (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[12]),
      (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[12]), (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[12]),
      (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[12]), (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[12]),
      (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[12]), (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[12]),
      {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_105_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_106_nl
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_13_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_108_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_109_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_110_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_111_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_112_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_113_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_114_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_115_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_116_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_117_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_118_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_119_nl});
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_90_cse
      = (~ operator_3_false_operator_3_false_operator_3_false_or_mdf_13_sva_1) &
      weight_mem_read_arbxbar_xbar_for_3_13_operator_7_false_operator_7_false_operator_7_false_or_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_92_cse
      = (~ operator_4_false_operator_4_false_operator_4_false_or_mdf_13_sva_1) &
      and_dcpl_1000;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_93_cse
      = operator_4_false_operator_4_false_operator_4_false_or_mdf_13_sva_1 & and_dcpl_1000;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_94_cse
      = (~ operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_13_sva_1)
      & and_dcpl_1001;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_95_cse
      = operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_13_sva_1
      & and_dcpl_1001;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_96_cse
      = (~ operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_13_sva_1)
      & and_dcpl_1008;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_97_cse
      = operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_13_sva_1
      & and_dcpl_1008;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_13_lpi_1_dfm_mx0
      = MUX1HOT_s_1_8_2(operator_2_false_operator_2_false_operator_2_false_or_mdf_13_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_30_13_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_13_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_13_sva_1, operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_13_sva_1,
      operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_13_sva_1, operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_13_sva_1,
      operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_13_sva_1, {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_90_cse
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_13_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_92_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_93_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_94_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_95_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_96_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_97_cse});
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_13_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(operator_3_false_operator_3_false_operator_3_false_or_mdf_13_sva_1,
      operator_4_false_operator_4_false_operator_4_false_or_mdf_13_sva_1, operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_13_sva_1,
      operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_13_sva_1, {weight_mem_read_arbxbar_xbar_for_3_13_operator_7_false_operator_7_false_operator_7_false_or_cse
      , and_dcpl_1000 , and_dcpl_1001 , and_dcpl_1008});
  assign weight_mem_read_arbxbar_xbar_for_3_13_operator_7_false_operator_7_false_operator_7_false_or_cse
      = Arbiter_16U_Roundrobin_pick_priority_30_13_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_13_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_13_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_13_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_13_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_13_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_13_sva_1;
  assign weight_mem_read_arbxbar_xbar_for_3_13_operator_8_false_operator_8_false_operator_8_false_or_nl
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[12])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[12])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[12])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[12]);
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_13_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_13_operator_8_false_operator_8_false_operator_8_false_or_nl,
      weight_mem_read_arbxbar_xbar_for_3_13_operator_7_false_operator_7_false_operator_7_false_or_cse,
      weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign Arbiter_16U_Roundrobin_pick_priority_25_13_sva_1 = weight_mem_read_arbxbar_arbiters_next_12_10_sva
      & (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[12]);
  assign Arbiter_16U_Roundrobin_pick_priority_27_13_sva_1 = weight_mem_read_arbxbar_arbiters_next_12_12_sva
      & (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[12]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_13_sva_1 = Arbiter_16U_Roundrobin_pick_priority_27_13_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_13_sva_1;
  assign operator_3_false_operator_3_false_operator_3_false_or_mdf_13_sva_1 = Arbiter_16U_Roundrobin_pick_priority_30_13_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_29_13_sva_1 | Arbiter_16U_Roundrobin_pick_priority_28_13_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_29_13_sva_1 = weight_mem_read_arbxbar_arbiters_next_12_14_sva
      & (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[12]);
  assign Arbiter_16U_Roundrobin_pick_priority_30_13_sva_1 = weight_mem_read_arbxbar_arbiters_next_12_15_sva
      & (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[12]);
  assign Arbiter_16U_Roundrobin_pick_priority_26_13_sva_1 = weight_mem_read_arbxbar_arbiters_next_12_11_sva
      & (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[12]);
  assign Arbiter_16U_Roundrobin_pick_priority_28_13_sva_1 = weight_mem_read_arbxbar_arbiters_next_12_13_sva
      & (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[12]);
  assign Arbiter_16U_Roundrobin_pick_priority_21_13_sva_1 = weight_mem_read_arbxbar_arbiters_next_12_6_sva
      & (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[12]);
  assign Arbiter_16U_Roundrobin_pick_priority_23_13_sva_1 = weight_mem_read_arbxbar_arbiters_next_12_8_sva
      & (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[12]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_13_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_23_13_sva_1 | Arbiter_16U_Roundrobin_pick_priority_22_13_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_17_13_sva_1 = weight_mem_read_arbxbar_arbiters_next_12_2_sva
      & (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[12]);
  assign Arbiter_16U_Roundrobin_pick_priority_19_13_sva_1 = weight_mem_read_arbxbar_arbiters_next_12_4_sva
      & (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[12]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_13_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_19_13_sva_1 | Arbiter_16U_Roundrobin_pick_priority_18_13_sva_1;
  assign operator_4_false_operator_4_false_operator_4_false_or_mdf_13_sva_1 = Arbiter_16U_Roundrobin_pick_priority_23_13_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_13_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_13_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_13_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_22_13_sva_1 = weight_mem_read_arbxbar_arbiters_next_12_7_sva
      & (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[12]);
  assign Arbiter_16U_Roundrobin_pick_priority_18_13_sva_1 = weight_mem_read_arbxbar_arbiters_next_12_3_sva
      & (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[12]);
  assign Arbiter_16U_Roundrobin_pick_priority_20_13_sva_1 = weight_mem_read_arbxbar_arbiters_next_12_5_sva
      & (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[12]);
  assign Arbiter_16U_Roundrobin_pick_priority_24_13_sva_1 = weight_mem_read_arbxbar_arbiters_next_12_9_sva
      & (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[12]);
  assign operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_13_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[12]);
  assign operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_13_sva_1
      = (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[12]);
  assign operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_13_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[12])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[12]);
  assign operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_13_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[12]);
  assign operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_13_sva_1
      = (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[12]);
  assign operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_13_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[12])
      | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[12]);
  assign weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp
      = Arbiter_16U_Roundrobin_pick_priority_30_13_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_13_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_13_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_13_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_13_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_13_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_13_sva_1 | Arbiter_16U_Roundrobin_pick_priority_23_13_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_13_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_13_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_13_sva_1 | Arbiter_16U_Roundrobin_pick_priority_19_13_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_18_13_sva_1 | Arbiter_16U_Roundrobin_pick_priority_17_13_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_12_1_sva & (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[12]));
  assign Arbiter_16U_Roundrobin_pick_mux_3163_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_0,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_0,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_12_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_15_0_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3163_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3162_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_1,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_1,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_12_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_15_1_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3162_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3160_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_3,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_3,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_12_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_15_2_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3160_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3156_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_7,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_7,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_12_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3156_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_14;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_14
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_13 & weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_13 & (~ weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_13
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_13 & weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_13 & (~ weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_12
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_13 & weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_13 & (~ weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_11
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_13 & weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_13 & (~ weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_10
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_13 & weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_13 & (~ weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_9
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_13 & weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_13 & (~ weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_8
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_13 & weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_13 & (~ weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_7
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_13 & weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_13 & (~ weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_6
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_13 & weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_13 & (~ weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_5
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_13 & weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_13 & (~ weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_4
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_13 & weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_13 & (~ weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_3
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_13 & weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_13 & (~ weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_2
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_13 & weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_13 & (~ weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_1
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_13 & weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_13 & (~ weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_0
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_13 & weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_13 & (~ weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_13_nl
      = Arbiter_16U_Roundrobin_pick_priority_29_14_sva_1 & (~ Arbiter_16U_Roundrobin_pick_priority_30_14_sva_1);
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_75_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_14_sva_1) &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_60_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_76_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_14_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_60_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_78_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_14_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_62_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_79_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_14_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_62_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_80_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_14_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_63_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_81_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_14_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_63_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_82_nl
      = (~ operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_14_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_64_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_83_nl
      = operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_14_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_64_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_84_nl
      = (~ operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_14_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_65_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_85_nl
      = operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_14_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_65_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_86_nl
      = (~ operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_14_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_66_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_87_nl
      = operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_14_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_66_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_88_nl
      = (~ operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_14_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_67_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_89_nl
      = operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_14_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_67_cse;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_14_lpi_1_dfm_mx0
      = MUX1HOT_s_1_15_2(Arbiter_16U_Roundrobin_pick_priority_25_14_sva_1, Arbiter_16U_Roundrobin_pick_priority_27_14_sva_1,
      nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_13_nl,
      Arbiter_16U_Roundrobin_pick_priority_17_14_sva_1, Arbiter_16U_Roundrobin_pick_priority_19_14_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_21_14_sva_1, Arbiter_16U_Roundrobin_pick_priority_23_14_sva_1,
      (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[13]), (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[13]),
      (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[13]), (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[13]),
      (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[13]), (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[13]),
      (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[13]), (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[13]),
      {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_75_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_76_nl
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_14_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_78_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_79_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_80_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_81_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_82_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_83_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_84_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_85_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_86_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_87_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_88_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_89_nl});
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_60_cse
      = (~ operator_3_false_operator_3_false_operator_3_false_or_mdf_14_sva_1) &
      weight_mem_read_arbxbar_xbar_for_3_14_operator_7_false_operator_7_false_operator_7_false_or_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_62_cse
      = (~ operator_4_false_operator_4_false_operator_4_false_or_mdf_14_sva_1) &
      and_dcpl_1023;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_63_cse
      = operator_4_false_operator_4_false_operator_4_false_or_mdf_14_sva_1 & and_dcpl_1023;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_64_cse
      = (~ operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_14_sva_1)
      & and_dcpl_1024;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_65_cse
      = operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_14_sva_1
      & and_dcpl_1024;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_66_cse
      = (~ operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_14_sva_1)
      & and_dcpl_1029;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_67_cse
      = operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_14_sva_1
      & and_dcpl_1029;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_14_lpi_1_dfm_mx0
      = MUX1HOT_s_1_8_2(operator_2_false_operator_2_false_operator_2_false_or_mdf_14_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_30_14_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_14_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_14_sva_1, operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_14_sva_1,
      operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_14_sva_1, operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_14_sva_1,
      operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_14_sva_1, {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_60_cse
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_14_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_62_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_63_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_64_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_65_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_66_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_67_cse});
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_14_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(operator_3_false_operator_3_false_operator_3_false_or_mdf_14_sva_1,
      operator_4_false_operator_4_false_operator_4_false_or_mdf_14_sva_1, operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_14_sva_1,
      operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_14_sva_1, {weight_mem_read_arbxbar_xbar_for_3_14_operator_7_false_operator_7_false_operator_7_false_or_cse
      , and_dcpl_1023 , and_dcpl_1024 , and_dcpl_1029});
  assign weight_mem_read_arbxbar_xbar_for_3_14_operator_7_false_operator_7_false_operator_7_false_or_cse
      = Arbiter_16U_Roundrobin_pick_priority_30_14_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_14_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_14_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_14_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_14_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_14_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_14_sva_1;
  assign weight_mem_read_arbxbar_xbar_for_3_14_operator_8_false_operator_8_false_operator_8_false_or_nl
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[13])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[13])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[13])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[13]);
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_14_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_14_operator_8_false_operator_8_false_operator_8_false_or_nl,
      weight_mem_read_arbxbar_xbar_for_3_14_operator_7_false_operator_7_false_operator_7_false_or_cse,
      weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign Arbiter_16U_Roundrobin_pick_priority_25_14_sva_1 = weight_mem_read_arbxbar_arbiters_next_13_10_sva
      & (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[13]);
  assign Arbiter_16U_Roundrobin_pick_priority_27_14_sva_1 = weight_mem_read_arbxbar_arbiters_next_13_12_sva
      & (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[13]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_14_sva_1 = Arbiter_16U_Roundrobin_pick_priority_27_14_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_14_sva_1;
  assign operator_3_false_operator_3_false_operator_3_false_or_mdf_14_sva_1 = Arbiter_16U_Roundrobin_pick_priority_30_14_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_29_14_sva_1 | Arbiter_16U_Roundrobin_pick_priority_28_14_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_29_14_sva_1 = weight_mem_read_arbxbar_arbiters_next_13_14_sva
      & (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[13]);
  assign Arbiter_16U_Roundrobin_pick_priority_30_14_sva_1 = weight_mem_read_arbxbar_arbiters_next_13_15_sva
      & (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[13]);
  assign Arbiter_16U_Roundrobin_pick_priority_26_14_sva_1 = weight_mem_read_arbxbar_arbiters_next_13_11_sva
      & (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[13]);
  assign Arbiter_16U_Roundrobin_pick_priority_28_14_sva_1 = weight_mem_read_arbxbar_arbiters_next_13_13_sva
      & (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[13]);
  assign Arbiter_16U_Roundrobin_pick_priority_21_14_sva_1 = weight_mem_read_arbxbar_arbiters_next_13_6_sva
      & (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[13]);
  assign Arbiter_16U_Roundrobin_pick_priority_23_14_sva_1 = weight_mem_read_arbxbar_arbiters_next_13_8_sva
      & (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[13]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_14_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_23_14_sva_1 | Arbiter_16U_Roundrobin_pick_priority_22_14_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_17_14_sva_1 = weight_mem_read_arbxbar_arbiters_next_13_2_sva
      & (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[13]);
  assign Arbiter_16U_Roundrobin_pick_priority_19_14_sva_1 = weight_mem_read_arbxbar_arbiters_next_13_4_sva
      & (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[13]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_14_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_19_14_sva_1 | Arbiter_16U_Roundrobin_pick_priority_18_14_sva_1;
  assign operator_4_false_operator_4_false_operator_4_false_or_mdf_14_sva_1 = Arbiter_16U_Roundrobin_pick_priority_23_14_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_14_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_14_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_14_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_22_14_sva_1 = weight_mem_read_arbxbar_arbiters_next_13_7_sva
      & (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[13]);
  assign Arbiter_16U_Roundrobin_pick_priority_18_14_sva_1 = weight_mem_read_arbxbar_arbiters_next_13_3_sva
      & (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[13]);
  assign Arbiter_16U_Roundrobin_pick_priority_20_14_sva_1 = weight_mem_read_arbxbar_arbiters_next_13_5_sva
      & (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[13]);
  assign Arbiter_16U_Roundrobin_pick_priority_24_14_sva_1 = weight_mem_read_arbxbar_arbiters_next_13_9_sva
      & (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[13]);
  assign operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_14_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[13]);
  assign operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_14_sva_1
      = (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[13]);
  assign operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_14_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[13])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[13]);
  assign operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_14_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[13]);
  assign operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_14_sva_1
      = (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[13]);
  assign operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_14_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[13])
      | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[13]);
  assign weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp
      = Arbiter_16U_Roundrobin_pick_priority_30_14_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_14_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_14_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_14_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_14_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_14_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_14_sva_1 | Arbiter_16U_Roundrobin_pick_priority_23_14_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_14_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_14_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_14_sva_1 | Arbiter_16U_Roundrobin_pick_priority_19_14_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_18_14_sva_1 | Arbiter_16U_Roundrobin_pick_priority_17_14_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_13_1_sva & (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[13]));
  assign Arbiter_16U_Roundrobin_pick_mux_3177_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_0,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_0,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_13_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_16_0_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3177_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3176_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_1,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_1,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_13_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_16_1_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3176_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3174_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_3,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_3,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_13_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_16_2_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3174_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3170_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_7,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_7,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_13_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3170_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_14;
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_14
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_14 & weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_14 & (~ weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_13
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_14 & weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_14 & (~ weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_12
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_14 & weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_14 & (~ weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_11
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_14 & weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_14 & (~ weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_10
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_14 & weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_14 & (~ weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_9
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_14 & weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_14 & (~ weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_8
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_14 & weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_14 & (~ weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_7
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_14 & weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_14 & (~ weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_6
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_14 & weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_14 & (~ weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_5
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_14 & weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_14 & (~ weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_4
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_14 & weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_14 & (~ weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_3
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_14 & weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_14 & (~ weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_2
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_14 & weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_14 & (~ weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_1
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_14 & weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_14 & (~ weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_0
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_14 & weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_14 & (~ weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_14_nl
      = Arbiter_16U_Roundrobin_pick_priority_29_15_sva_1 & (~ Arbiter_16U_Roundrobin_pick_priority_30_15_sva_1);
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_45_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_15_sva_1) &
      nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_30_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_46_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_15_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_30_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_48_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_15_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_32_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_49_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_15_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_32_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_50_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_15_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_33_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_51_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_15_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_33_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_52_nl
      = (~ operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_15_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_34_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_53_nl
      = operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_15_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_34_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_54_nl
      = (~ operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_15_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_35_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_55_nl
      = operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_15_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_35_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_56_nl
      = (~ operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_15_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_36_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_57_nl
      = operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_15_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_36_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_58_nl
      = (~ operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_15_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_37_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_59_nl
      = operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_15_sva_1
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_37_cse;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_15_lpi_1_dfm_mx0
      = MUX1HOT_s_1_15_2(Arbiter_16U_Roundrobin_pick_priority_25_15_sva_1, Arbiter_16U_Roundrobin_pick_priority_27_15_sva_1,
      nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_14_nl,
      Arbiter_16U_Roundrobin_pick_priority_17_15_sva_1, Arbiter_16U_Roundrobin_pick_priority_19_15_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_21_15_sva_1, Arbiter_16U_Roundrobin_pick_priority_23_15_sva_1,
      (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[14]), (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[14]),
      (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[14]), (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[14]),
      (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[14]), (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[14]),
      (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[14]), (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[14]),
      {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_45_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_46_nl
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_15_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_48_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_49_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_50_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_51_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_52_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_53_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_54_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_55_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_56_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_57_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_58_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_59_nl});
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_30_cse
      = (~ operator_3_false_operator_3_false_operator_3_false_or_mdf_15_sva_1) &
      weight_mem_read_arbxbar_xbar_for_3_15_operator_7_false_operator_7_false_operator_7_false_or_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_32_cse
      = (~ operator_4_false_operator_4_false_operator_4_false_or_mdf_15_sva_1) &
      and_dcpl_1043;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_33_cse
      = operator_4_false_operator_4_false_operator_4_false_or_mdf_15_sva_1 & and_dcpl_1043;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_34_cse
      = (~ operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_15_sva_1)
      & and_dcpl_1044;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_35_cse
      = operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_15_sva_1
      & and_dcpl_1044;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_36_cse
      = (~ operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_15_sva_1)
      & and_dcpl_1051;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_37_cse
      = operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_15_sva_1
      & and_dcpl_1051;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_15_lpi_1_dfm_mx0
      = MUX1HOT_s_1_8_2(operator_2_false_operator_2_false_operator_2_false_or_mdf_15_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_30_15_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_15_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_15_sva_1, operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_15_sva_1,
      operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_15_sva_1, operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_15_sva_1,
      operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_15_sva_1, {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_30_cse
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_15_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_32_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_33_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_34_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_35_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_36_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_37_cse});
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_15_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(operator_3_false_operator_3_false_operator_3_false_or_mdf_15_sva_1,
      operator_4_false_operator_4_false_operator_4_false_or_mdf_15_sva_1, operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_15_sva_1,
      operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_15_sva_1, {weight_mem_read_arbxbar_xbar_for_3_15_operator_7_false_operator_7_false_operator_7_false_or_cse
      , and_dcpl_1043 , and_dcpl_1044 , and_dcpl_1051});
  assign weight_mem_read_arbxbar_xbar_for_3_15_operator_7_false_operator_7_false_operator_7_false_or_cse
      = Arbiter_16U_Roundrobin_pick_priority_30_15_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_15_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_15_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_15_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_15_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_15_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_15_Arbiter_16U_Roundrobin_pick_priority_and_4_tmp;
  assign weight_mem_read_arbxbar_xbar_for_3_15_operator_8_false_operator_8_false_operator_8_false_or_nl
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[14])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[14])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[14])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[14]);
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_15_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_15_operator_8_false_operator_8_false_operator_8_false_or_nl,
      weight_mem_read_arbxbar_xbar_for_3_15_operator_7_false_operator_7_false_operator_7_false_or_cse,
      weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign Arbiter_16U_Roundrobin_pick_priority_25_15_sva_1 = weight_mem_read_arbxbar_arbiters_next_14_10_sva
      & (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[14]);
  assign Arbiter_16U_Roundrobin_pick_priority_27_15_sva_1 = weight_mem_read_arbxbar_arbiters_next_14_12_sva
      & (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[14]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_15_sva_1 = Arbiter_16U_Roundrobin_pick_priority_27_15_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_15_sva_1;
  assign operator_3_false_operator_3_false_operator_3_false_or_mdf_15_sva_1 = Arbiter_16U_Roundrobin_pick_priority_30_15_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_29_15_sva_1 | Arbiter_16U_Roundrobin_pick_priority_28_15_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_29_15_sva_1 = weight_mem_read_arbxbar_arbiters_next_14_14_sva
      & (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[14]);
  assign Arbiter_16U_Roundrobin_pick_priority_30_15_sva_1 = weight_mem_read_arbxbar_arbiters_next_14_15_sva
      & (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[14]);
  assign Arbiter_16U_Roundrobin_pick_priority_26_15_sva_1 = weight_mem_read_arbxbar_arbiters_next_14_11_sva
      & (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[14]);
  assign Arbiter_16U_Roundrobin_pick_priority_28_15_sva_1 = weight_mem_read_arbxbar_arbiters_next_14_13_sva
      & (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[14]);
  assign Arbiter_16U_Roundrobin_pick_priority_21_15_sva_1 = weight_mem_read_arbxbar_arbiters_next_14_6_sva
      & (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[14]);
  assign Arbiter_16U_Roundrobin_pick_priority_23_15_sva_1 = weight_mem_read_arbxbar_arbiters_next_14_8_sva
      & (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[14]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_15_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_23_15_sva_1 | Arbiter_16U_Roundrobin_pick_priority_22_15_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_17_15_sva_1 = weight_mem_read_arbxbar_arbiters_next_14_2_sva
      & (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[14]);
  assign Arbiter_16U_Roundrobin_pick_priority_19_15_sva_1 = weight_mem_read_arbxbar_arbiters_next_14_4_sva
      & (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[14]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_15_sva_1
      = Arbiter_16U_Roundrobin_pick_priority_19_15_sva_1 | Arbiter_16U_Roundrobin_pick_priority_18_15_sva_1;
  assign operator_4_false_operator_4_false_operator_4_false_or_mdf_15_sva_1 = Arbiter_16U_Roundrobin_pick_priority_23_15_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_15_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_15_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_15_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_22_15_sva_1 = weight_mem_read_arbxbar_arbiters_next_14_7_sva
      & (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[14]);
  assign Arbiter_16U_Roundrobin_pick_priority_18_15_sva_1 = weight_mem_read_arbxbar_arbiters_next_14_3_sva
      & (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[14]);
  assign Arbiter_16U_Roundrobin_pick_priority_20_15_sva_1 = weight_mem_read_arbxbar_arbiters_next_14_5_sva
      & (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[14]);
  assign weight_mem_read_arbxbar_xbar_for_3_15_Arbiter_16U_Roundrobin_pick_priority_and_4_tmp
      = weight_mem_read_arbxbar_arbiters_next_14_9_sva & (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[14]);
  assign operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_15_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[14]);
  assign operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_15_sva_1
      = (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[14]);
  assign operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_15_sva_1
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[14])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[14]);
  assign operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_15_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[14]);
  assign operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_15_sva_1
      = (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[14]);
  assign operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_15_sva_1
      = (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[14])
      | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[14]);
  assign weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp
      = Arbiter_16U_Roundrobin_pick_priority_30_15_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_15_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_15_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_15_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_15_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_15_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_15_Arbiter_16U_Roundrobin_pick_priority_and_4_tmp
      | Arbiter_16U_Roundrobin_pick_priority_23_15_sva_1 | Arbiter_16U_Roundrobin_pick_priority_22_15_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_21_15_sva_1 | Arbiter_16U_Roundrobin_pick_priority_20_15_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_19_15_sva_1 | Arbiter_16U_Roundrobin_pick_priority_18_15_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_17_15_sva_1 | (weight_mem_read_arbxbar_arbiters_next_14_1_sva
      & (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[14]));
  assign Arbiter_16U_Roundrobin_pick_mux_3191_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_0,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_0,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_14_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_17_0_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3191_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3190_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_1,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_1,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_14_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_17_1_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3190_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3188_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_3,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_3,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_14_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_17_2_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3188_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3184_nl = MUX_s_1_2_2(nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_7,
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_7,
      Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_14_tmp);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3184_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_14;
  assign weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_itm
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_15 & weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_15 & (~ weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_1_itm
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_15 & weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_15 & (~ weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_2_itm
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_15 & weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_15 & (~ weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_3_itm
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_15 & weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_15 & (~ weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_4_itm
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_15 & weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_15 & (~ weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_5_itm
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_15 & weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_15 & (~ weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_6_itm
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_15 & weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_15 & (~ weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_7_itm
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_15 & weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_15 & (~ weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_8_itm
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_15 & weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_15 & (~ weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_9_itm
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_15 & weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_15 & (~ weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_10_itm
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_15 & weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_15 & (~ weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_11_itm
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_15 & weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_15 & (~ weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_12_itm
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_15 & weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_15 & (~ weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_13_itm
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_15 & weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_15 & (~ weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_14_itm
      = (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_15 & weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp)
      | (Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_15 & (~ weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_15_nl
      = Arbiter_16U_Roundrobin_pick_priority_29_sva_1 & (~ Arbiter_16U_Roundrobin_pick_priority_30_sva_1);
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_15_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_sva_1) & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_16_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_18_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_2_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_19_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_2_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_20_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_3_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_21_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_3_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_22_nl
      = (~ operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_4_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_23_nl
      = operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_4_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_24_nl
      = (~ operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_5_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_25_nl
      = operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_5_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_26_nl
      = (~ operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_6_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_27_nl
      = operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_6_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_28_nl
      = (~ operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_sva_1)
      & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_7_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_29_nl
      = operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_sva_1 & nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_7_cse;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_lpi_1_dfm_mx0
      = MUX1HOT_s_1_15_2(Arbiter_16U_Roundrobin_pick_priority_25_sva_1, Arbiter_16U_Roundrobin_pick_priority_27_sva_1,
      nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_15_nl,
      Arbiter_16U_Roundrobin_pick_priority_17_sva_1, Arbiter_16U_Roundrobin_pick_priority_19_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_21_sva_1, Arbiter_16U_Roundrobin_pick_priority_23_sva_1,
      (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[15]), (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[15]),
      (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[15]), (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[15]),
      (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[15]), (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[15]),
      (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[15]), (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[15]),
      {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_15_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_16_nl
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_18_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_19_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_20_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_21_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_22_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_23_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_24_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_25_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_26_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_27_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_28_nl
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_29_nl});
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_cse
      = (~ operator_3_false_operator_3_false_operator_3_false_or_mdf_sva_1) & weight_mem_read_arbxbar_xbar_for_3_16_operator_7_false_operator_7_false_operator_7_false_or_cse;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_2_cse
      = (~ operator_4_false_operator_4_false_operator_4_false_or_mdf_sva_1) & and_dcpl_1066;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_3_cse
      = operator_4_false_operator_4_false_operator_4_false_or_mdf_sva_1 & and_dcpl_1066;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_4_cse
      = (~ operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_sva_1)
      & and_dcpl_1067;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_5_cse
      = operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_sva_1 & and_dcpl_1067;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_6_cse
      = (~ operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_sva_1)
      & and_dcpl_1074;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_7_cse
      = operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_sva_1 & and_dcpl_1074;
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_8_2(operator_2_false_operator_2_false_operator_2_false_or_mdf_sva_1,
      Arbiter_16U_Roundrobin_pick_priority_30_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_sva_1, operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_sva_1,
      operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_sva_1, operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_sva_1,
      operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_sva_1, {nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_cse
      , operator_3_false_operator_3_false_operator_3_false_or_mdf_sva_1 , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_2_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_3_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_4_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_5_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_6_cse
      , nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_7_cse});
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(operator_3_false_operator_3_false_operator_3_false_or_mdf_sva_1,
      operator_4_false_operator_4_false_operator_4_false_or_mdf_sva_1, operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_sva_1,
      operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_sva_1, {weight_mem_read_arbxbar_xbar_for_3_16_operator_7_false_operator_7_false_operator_7_false_or_cse
      , and_dcpl_1066 , and_dcpl_1067 , and_dcpl_1074});
  assign weight_mem_read_arbxbar_xbar_for_3_16_operator_7_false_operator_7_false_operator_7_false_or_cse
      = Arbiter_16U_Roundrobin_pick_priority_30_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_sva_1;
  assign weight_mem_read_arbxbar_xbar_for_3_16_operator_8_false_operator_8_false_operator_8_false_or_nl
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[15])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[15])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[15])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[15]);
  assign nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_for_3_16_operator_8_false_operator_8_false_operator_8_false_or_nl,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_7_false_operator_7_false_operator_7_false_or_cse,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign Arbiter_16U_Roundrobin_pick_priority_25_sva_1 = weight_mem_read_arbxbar_arbiters_next_15_10_sva
      & (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[15]);
  assign Arbiter_16U_Roundrobin_pick_priority_27_sva_1 = weight_mem_read_arbxbar_arbiters_next_15_12_sva
      & (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[15]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_sva_1 = Arbiter_16U_Roundrobin_pick_priority_27_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_sva_1;
  assign operator_3_false_operator_3_false_operator_3_false_or_mdf_sva_1 = Arbiter_16U_Roundrobin_pick_priority_30_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_29_sva_1 | Arbiter_16U_Roundrobin_pick_priority_28_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_29_sva_1 = weight_mem_read_arbxbar_arbiters_next_15_14_sva
      & (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[15]);
  assign Arbiter_16U_Roundrobin_pick_priority_30_sva_1 = weight_mem_read_arbxbar_arbiters_next_15_15_sva
      & (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[15]);
  assign Arbiter_16U_Roundrobin_pick_priority_26_sva_1 = weight_mem_read_arbxbar_arbiters_next_15_11_sva
      & (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[15]);
  assign Arbiter_16U_Roundrobin_pick_priority_28_sva_1 = weight_mem_read_arbxbar_arbiters_next_15_13_sva
      & (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[15]);
  assign Arbiter_16U_Roundrobin_pick_priority_21_sva_1 = weight_mem_read_arbxbar_arbiters_next_15_6_sva
      & (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[15]);
  assign Arbiter_16U_Roundrobin_pick_priority_23_sva_1 = weight_mem_read_arbxbar_arbiters_next_15_8_sva
      & (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[15]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_sva_1 =
      Arbiter_16U_Roundrobin_pick_priority_23_sva_1 | Arbiter_16U_Roundrobin_pick_priority_22_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_17_sva_1 = weight_mem_read_arbxbar_arbiters_next_15_2_sva
      & (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[15]);
  assign Arbiter_16U_Roundrobin_pick_priority_19_sva_1 = weight_mem_read_arbxbar_arbiters_next_15_4_sva
      & (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[15]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_sva_1 =
      Arbiter_16U_Roundrobin_pick_priority_19_sva_1 | Arbiter_16U_Roundrobin_pick_priority_18_sva_1;
  assign operator_4_false_operator_4_false_operator_4_false_or_mdf_sva_1 = Arbiter_16U_Roundrobin_pick_priority_23_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_sva_1;
  assign Arbiter_16U_Roundrobin_pick_priority_22_sva_1 = weight_mem_read_arbxbar_arbiters_next_15_7_sva
      & (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[15]);
  assign Arbiter_16U_Roundrobin_pick_priority_18_sva_1 = weight_mem_read_arbxbar_arbiters_next_15_3_sva
      & (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[15]);
  assign Arbiter_16U_Roundrobin_pick_priority_20_sva_1 = weight_mem_read_arbxbar_arbiters_next_15_5_sva
      & (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[15]);
  assign Arbiter_16U_Roundrobin_pick_priority_24_sva_1 = weight_mem_read_arbxbar_arbiters_next_15_9_sva
      & (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[15]);
  assign operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_sva_1 =
      (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[15]);
  assign operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_sva_1 =
      (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[15]);
  assign operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_sva_1 =
      (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[15])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[15]);
  assign operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_sva_1 =
      (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[15]);
  assign operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_sva_1 =
      (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[15]);
  assign operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_sva_1 =
      (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[15])
      | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[15]);
  assign weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp
      = Arbiter_16U_Roundrobin_pick_priority_30_sva_1 | Arbiter_16U_Roundrobin_pick_priority_29_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_28_sva_1 | Arbiter_16U_Roundrobin_pick_priority_27_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_26_sva_1 | Arbiter_16U_Roundrobin_pick_priority_25_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_24_sva_1 | Arbiter_16U_Roundrobin_pick_priority_23_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_22_sva_1 | Arbiter_16U_Roundrobin_pick_priority_21_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_20_sva_1 | Arbiter_16U_Roundrobin_pick_priority_19_sva_1
      | Arbiter_16U_Roundrobin_pick_priority_18_sva_1 | Arbiter_16U_Roundrobin_pick_priority_17_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_15_1_sva & (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[15]));
  assign Arbiter_16U_Roundrobin_pick_mux_3216_nl = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_11,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_11_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_2_2_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3216_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3218_nl = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_13,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_13_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_2_1_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3218_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_14;
  assign Arbiter_16U_Roundrobin_pick_mux_3219_nl = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_14,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_14_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign weight_mem_read_arbxbar_xbar_for_3_source_local_2_0_sva_1 = Arbiter_16U_Roundrobin_pick_mux_3219_nl
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_14;
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_lpi_1_dfm_1 = MUX_v_4_2_2(4'b0000,
      (weight_read_addrs_15_lpi_1_dfm_3[3:0]), weight_read_ack_15_lpi_1_dfm_15_mx0);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_15_lpi_1_dfm_1_3_1 =
      MUX_v_3_2_2(3'b000, (weight_read_addrs_14_15_1_lpi_1_dfm_3[2:0]), weight_read_ack_14_lpi_1_dfm_15_mx0);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_15_lpi_1_dfm_1_0 = (PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx1[0])
      & (~ pe_config_is_cluster_sva) & PECore_RunFSM_switch_lp_equal_tmp_5 & weight_read_ack_14_lpi_1_dfm_15_mx0;
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_14_lpi_1_dfm_1 = MUX_v_4_2_2(4'b0000,
      (weight_read_addrs_13_lpi_1_dfm_3[3:0]), weight_read_ack_13_lpi_1_dfm_15_mx0);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_13_3_2_lpi_1_dfm_1 =
      MUX_v_2_2_2(2'b00, (weight_read_addrs_12_15_2_lpi_1_dfm_3[1:0]), weight_read_ack_12_lpi_1_dfm_15_mx0);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_13_1_0_lpi_1_dfm_1 =
      (weight_read_addrs_8_2_0_lpi_1_dfm_1[1:0]) & ({{1{PECore_RunFSM_switch_lp_equal_tmp_5}},
      PECore_RunFSM_switch_lp_equal_tmp_5}) & ({{1{weight_read_ack_12_lpi_1_dfm_15_mx0}},
      weight_read_ack_12_lpi_1_dfm_15_mx0});
  assign weight_mem_run_1_if_for_if_and_697_nl = weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_236_tmp
      & (~(weight_mem_run_1_if_for_if_and_stg_2_4_15_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_2_3_sva_1));
  assign weight_read_ack_12_lpi_1_dfm_15_mx0 = MUX_s_1_2_2(weight_mem_run_1_if_for_if_and_697_nl,
      weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_236_tmp, or_dcpl_34);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_12_lpi_1_dfm_1 = MUX_v_4_2_2(4'b0000,
      (weight_read_addrs_11_lpi_1_dfm_3[3:0]), weight_read_ack_11_lpi_1_dfm_15_mx0);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_3_1_lpi_1_dfm_1 =
      MUX_v_3_2_2(3'b000, (weight_read_addrs_10_15_1_lpi_1_dfm_3[2:0]), weight_read_ack_10_lpi_1_dfm_15_mx0);
  assign weight_mem_run_1_if_for_if_and_693_nl = weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_234_tmp
      & (~(weight_mem_run_1_if_for_if_and_stg_2_2_15_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_2_3_sva_1));
  assign weight_read_ack_10_lpi_1_dfm_15_mx0 = MUX_s_1_2_2(weight_mem_run_1_if_for_if_and_693_nl,
      weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_234_tmp, or_dcpl_34);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_2_0_lpi_1_dfm_1 =
      weight_read_addrs_8_2_0_lpi_1_dfm_1 & ({{2{PECore_RunFSM_switch_lp_equal_tmp_5}},
      PECore_RunFSM_switch_lp_equal_tmp_5}) & ({{2{weight_read_ack_8_lpi_1_dfm_15_mx0}},
      weight_read_ack_8_lpi_1_dfm_15_mx0});
  assign weight_mem_run_1_if_for_if_and_689_nl = weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_232_tmp
      & (~(weight_mem_run_1_if_for_if_and_stg_2_0_15_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_2_3_sva_1));
  assign weight_read_ack_8_lpi_1_dfm_15_mx0 = MUX_s_1_2_2(weight_mem_run_1_if_for_if_and_689_nl,
      weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_232_tmp, or_dcpl_34);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_8_lpi_1_dfm_1 = MUX_v_4_2_2(4'b0000,
      (weight_read_addrs_7_lpi_1_dfm_2[3:0]), weight_read_ack_7_lpi_1_dfm_15_mx0);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_3_1_lpi_1_dfm_1 =
      MUX_v_3_2_2(3'b000, (weight_read_addrs_6_15_1_lpi_1_dfm_2[2:0]), weight_read_ack_6_lpi_1_dfm_15_mx0);
  assign weight_mem_run_1_if_for_if_and_690_nl = weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_230_tmp
      & (~(weight_mem_run_1_if_for_if_and_stg_2_6_15_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_2_3_sva_1)));
  assign weight_read_ack_6_lpi_1_dfm_15_mx0 = MUX_s_1_2_2(weight_mem_run_1_if_for_if_and_690_nl,
      weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_230_tmp, or_dcpl_34);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_6_lpi_1_dfm_1 = MUX_v_4_2_2(4'b0000,
      (weight_read_addrs_5_lpi_1_dfm_2[3:0]), weight_read_ack_5_lpi_1_dfm_15_mx0);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_5_3_2_lpi_1_dfm_1 =
      MUX_v_2_2_2(2'b00, (weight_read_addrs_4_15_2_lpi_1_dfm_2[1:0]), weight_read_ack_4_lpi_1_dfm_15_mx0);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_5_1_0_lpi_1_dfm_1 =
      MUX_v_2_2_2(2'b00, weight_read_addrs_4_1_0_lpi_1_dfm_1, weight_read_ack_4_lpi_1_dfm_15_mx0);
  assign weight_mem_run_1_if_for_if_and_694_nl = weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_228_tmp
      & (~(weight_mem_run_1_if_for_if_and_stg_2_4_15_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_2_3_sva_1)));
  assign weight_read_ack_4_lpi_1_dfm_15_mx0 = MUX_s_1_2_2(weight_mem_run_1_if_for_if_and_694_nl,
      weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_228_tmp, or_dcpl_34);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_4_lpi_1_dfm_1 = MUX_v_4_2_2(4'b0000,
      (weight_read_addrs_3_lpi_1_dfm_2[3:0]), weight_read_ack_3_lpi_1_dfm_15_mx0);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_3_1_lpi_1_dfm_1 =
      MUX_v_3_2_2(3'b000, (weight_read_addrs_2_15_1_lpi_1_dfm_2[2:0]), weight_read_ack_2_lpi_1_dfm_15_mx0);
  assign weight_mem_run_1_if_for_if_and_698_nl = weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_226_tmp
      & (~(weight_mem_run_1_if_for_if_and_stg_2_2_15_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_2_3_sva_1)));
  assign weight_read_ack_2_lpi_1_dfm_15_mx0 = MUX_s_1_2_2(weight_mem_run_1_if_for_if_and_698_nl,
      weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_226_tmp, or_dcpl_34);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_2_lpi_1_dfm_1 = MUX_v_4_2_2(4'b0000,
      (weight_read_addrs_1_lpi_1_dfm_2[3:0]), weight_read_ack_1_lpi_1_dfm_15_mx0);
  assign weight_mem_run_1_if_for_if_and_stg_2_1_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_3_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_2_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_3_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_3_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_3_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_4_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_3_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_5_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_3_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_6_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_3_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_7_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_3_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_0_sva_1 = ~(weight_mem_read_arbxbar_xbar_for_3_source_local_3_0_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_source_local_3_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_1_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_3_0_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_3_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_2_sva_1 = (~ weight_mem_read_arbxbar_xbar_for_3_source_local_3_0_sva_1)
      & weight_mem_read_arbxbar_xbar_for_3_source_local_3_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_3_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_3_0_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_3_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_1_1_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_1_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_4_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_2_1_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_1_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_4_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_3_1_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_1_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_4_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_4_1_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_1_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_4_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_5_1_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_1_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_4_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_6_1_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_1_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_4_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_7_1_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_1_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_4_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_0_1_sva_1 = ~(weight_mem_read_arbxbar_xbar_for_3_source_local_4_0_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_source_local_4_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_1_1_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_4_0_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_4_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_2_1_sva_1 = (~ weight_mem_read_arbxbar_xbar_for_3_source_local_4_0_sva_1)
      & weight_mem_read_arbxbar_xbar_for_3_source_local_4_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_3_1_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_4_0_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_4_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_1_2_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_2_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_5_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_2_2_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_2_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_5_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_3_2_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_2_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_5_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_4_2_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_2_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_5_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_5_2_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_2_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_5_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_6_2_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_2_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_5_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_7_2_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_2_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_5_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_0_2_sva_1 = ~(weight_mem_read_arbxbar_xbar_for_3_source_local_5_0_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_source_local_5_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_1_2_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_5_0_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_5_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_2_2_sva_1 = (~ weight_mem_read_arbxbar_xbar_for_3_source_local_5_0_sva_1)
      & weight_mem_read_arbxbar_xbar_for_3_source_local_5_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_3_2_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_5_0_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_5_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_1_3_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_3_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_6_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_2_3_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_3_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_6_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_3_3_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_3_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_6_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_4_3_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_3_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_6_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_5_3_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_3_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_6_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_6_3_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_3_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_6_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_7_3_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_3_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_6_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_0_3_sva_1 = ~(weight_mem_read_arbxbar_xbar_for_3_source_local_6_0_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_source_local_6_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_1_3_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_6_0_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_6_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_2_3_sva_1 = (~ weight_mem_read_arbxbar_xbar_for_3_source_local_6_0_sva_1)
      & weight_mem_read_arbxbar_xbar_for_3_source_local_6_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_3_3_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_6_0_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_6_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_1_4_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_4_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_7_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_2_4_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_4_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_7_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_3_4_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_4_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_7_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_4_4_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_4_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_7_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_5_4_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_4_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_7_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_6_4_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_4_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_7_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_7_4_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_4_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_7_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_0_4_sva_1 = ~(weight_mem_read_arbxbar_xbar_for_3_source_local_7_0_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_source_local_7_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_1_4_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_7_0_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_7_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_2_4_sva_1 = (~ weight_mem_read_arbxbar_xbar_for_3_source_local_7_0_sva_1)
      & weight_mem_read_arbxbar_xbar_for_3_source_local_7_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_3_4_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_7_0_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_7_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_1_5_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_5_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_8_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_2_5_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_5_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_8_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_3_5_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_5_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_8_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_4_5_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_5_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_8_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_5_5_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_5_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_8_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_6_5_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_5_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_8_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_7_5_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_5_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_8_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_0_5_sva_1 = ~(weight_mem_read_arbxbar_xbar_for_3_source_local_8_0_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_source_local_8_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_1_5_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_8_0_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_8_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_2_5_sva_1 = (~ weight_mem_read_arbxbar_xbar_for_3_source_local_8_0_sva_1)
      & weight_mem_read_arbxbar_xbar_for_3_source_local_8_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_3_5_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_8_0_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_8_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_1_6_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_6_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_9_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_2_6_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_6_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_9_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_3_6_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_6_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_9_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_4_6_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_6_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_9_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_5_6_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_6_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_9_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_6_6_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_6_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_9_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_7_6_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_6_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_9_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_0_6_sva_1 = ~(weight_mem_read_arbxbar_xbar_for_3_source_local_9_0_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_source_local_9_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_1_6_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_9_0_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_9_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_2_6_sva_1 = (~ weight_mem_read_arbxbar_xbar_for_3_source_local_9_0_sva_1)
      & weight_mem_read_arbxbar_xbar_for_3_source_local_9_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_3_6_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_9_0_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_9_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_1_7_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_7_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_10_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_2_7_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_7_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_10_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_3_7_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_7_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_10_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_4_7_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_7_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_10_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_5_7_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_7_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_10_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_6_7_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_7_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_10_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_7_7_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_7_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_10_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_0_7_sva_1 = ~(weight_mem_read_arbxbar_xbar_for_3_source_local_10_0_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_source_local_10_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_1_7_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_10_0_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_10_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_2_7_sva_1 = (~ weight_mem_read_arbxbar_xbar_for_3_source_local_10_0_sva_1)
      & weight_mem_read_arbxbar_xbar_for_3_source_local_10_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_3_7_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_10_0_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_10_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_1_8_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_8_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_11_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_2_8_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_8_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_11_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_3_8_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_8_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_11_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_4_8_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_8_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_11_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_5_8_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_8_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_11_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_6_8_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_8_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_11_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_7_8_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_8_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_11_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_0_8_sva_1 = ~(weight_mem_read_arbxbar_xbar_for_3_source_local_11_0_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_source_local_11_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_1_8_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_11_0_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_11_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_2_8_sva_1 = (~ weight_mem_read_arbxbar_xbar_for_3_source_local_11_0_sva_1)
      & weight_mem_read_arbxbar_xbar_for_3_source_local_11_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_3_8_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_11_0_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_11_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_1_9_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_9_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_12_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_2_9_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_9_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_12_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_3_9_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_9_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_12_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_4_9_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_9_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_12_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_5_9_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_9_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_12_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_6_9_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_9_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_12_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_7_9_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_9_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_12_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_0_9_sva_1 = ~(weight_mem_read_arbxbar_xbar_for_3_source_local_12_0_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_source_local_12_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_1_9_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_12_0_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_12_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_2_9_sva_1 = (~ weight_mem_read_arbxbar_xbar_for_3_source_local_12_0_sva_1)
      & weight_mem_read_arbxbar_xbar_for_3_source_local_12_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_3_9_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_12_0_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_12_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_1_10_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_10_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_13_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_2_10_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_10_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_13_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_3_10_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_10_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_13_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_4_10_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_10_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_13_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_5_10_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_10_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_13_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_6_10_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_10_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_13_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_7_10_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_10_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_13_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_0_10_sva_1 = ~(weight_mem_read_arbxbar_xbar_for_3_source_local_13_0_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_source_local_13_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_1_10_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_13_0_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_13_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_2_10_sva_1 = (~ weight_mem_read_arbxbar_xbar_for_3_source_local_13_0_sva_1)
      & weight_mem_read_arbxbar_xbar_for_3_source_local_13_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_3_10_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_13_0_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_13_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_1_11_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_11_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_14_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_2_11_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_11_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_14_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_3_11_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_11_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_14_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_4_11_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_11_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_14_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_5_11_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_11_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_14_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_6_11_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_11_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_14_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_7_11_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_11_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_14_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_0_11_sva_1 = ~(weight_mem_read_arbxbar_xbar_for_3_source_local_14_0_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_source_local_14_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_1_11_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_14_0_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_14_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_2_11_sva_1 = (~ weight_mem_read_arbxbar_xbar_for_3_source_local_14_0_sva_1)
      & weight_mem_read_arbxbar_xbar_for_3_source_local_14_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_3_11_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_14_0_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_14_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_1_12_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_12_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_15_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_2_12_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_12_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_15_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_3_12_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_12_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_15_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_4_12_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_12_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_15_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_5_12_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_12_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_15_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_6_12_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_12_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_15_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_7_12_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_12_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_15_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_0_12_sva_1 = ~(weight_mem_read_arbxbar_xbar_for_3_source_local_15_0_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_source_local_15_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_1_12_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_15_0_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_15_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_2_12_sva_1 = (~ weight_mem_read_arbxbar_xbar_for_3_source_local_15_0_sva_1)
      & weight_mem_read_arbxbar_xbar_for_3_source_local_15_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_3_12_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_15_0_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_15_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_1_13_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_13_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_16_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_2_13_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_13_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_16_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_3_13_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_13_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_16_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_4_13_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_13_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_16_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_5_13_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_13_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_16_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_6_13_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_13_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_16_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_7_13_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_13_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_16_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_0_13_sva_1 = ~(weight_mem_read_arbxbar_xbar_for_3_source_local_16_0_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_source_local_16_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_1_13_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_16_0_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_16_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_2_13_sva_1 = (~ weight_mem_read_arbxbar_xbar_for_3_source_local_16_0_sva_1)
      & weight_mem_read_arbxbar_xbar_for_3_source_local_16_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_3_13_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_16_0_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_16_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_1_14_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_14_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_17_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_2_14_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_14_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_17_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_3_14_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_14_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_17_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_2_4_14_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_14_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_17_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_5_14_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_14_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_17_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_6_14_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_14_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_17_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_2_7_14_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_14_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_17_2_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_0_14_sva_1 = ~(weight_mem_read_arbxbar_xbar_for_3_source_local_17_0_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_source_local_17_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_1_14_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_17_0_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_17_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_2_14_sva_1 = (~ weight_mem_read_arbxbar_xbar_for_3_source_local_17_0_sva_1)
      & weight_mem_read_arbxbar_xbar_for_3_source_local_17_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_3_14_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_17_0_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_17_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_703_nl = weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_239_tmp
      & (~(weight_mem_run_1_if_for_if_and_stg_2_7_15_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_2_3_sva_1));
  assign weight_read_ack_15_lpi_1_dfm_15_mx0 = MUX_s_1_2_2(weight_mem_run_1_if_for_if_and_703_nl,
      weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_239_tmp, or_dcpl_34);
  assign weight_mem_run_1_if_for_if_and_701_nl = weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_238_tmp
      & (~(weight_mem_run_1_if_for_if_and_stg_2_6_15_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_2_3_sva_1));
  assign weight_read_ack_14_lpi_1_dfm_15_mx0 = MUX_s_1_2_2(weight_mem_run_1_if_for_if_and_701_nl,
      weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_238_tmp, or_dcpl_34);
  assign weight_mem_run_1_if_for_if_and_699_nl = weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_237_tmp
      & (~(weight_mem_run_1_if_for_if_and_stg_2_5_15_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_2_3_sva_1));
  assign weight_read_ack_13_lpi_1_dfm_15_mx0 = MUX_s_1_2_2(weight_mem_run_1_if_for_if_and_699_nl,
      weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_237_tmp, or_dcpl_34);
  assign weight_mem_run_1_if_for_if_and_695_nl = weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_235_tmp
      & (~(weight_mem_run_1_if_for_if_and_stg_2_3_15_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_2_3_sva_1));
  assign weight_read_ack_11_lpi_1_dfm_15_mx0 = MUX_s_1_2_2(weight_mem_run_1_if_for_if_and_695_nl,
      weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_235_tmp, or_dcpl_34);
  assign weight_mem_run_1_if_for_if_and_688_nl = weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_231_tmp
      & (~(weight_mem_run_1_if_for_if_and_stg_2_7_15_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_2_3_sva_1)));
  assign weight_read_ack_7_lpi_1_dfm_15_mx0 = MUX_s_1_2_2(weight_mem_run_1_if_for_if_and_688_nl,
      weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_231_tmp, or_dcpl_34);
  assign weight_mem_run_1_if_for_if_and_692_nl = weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_229_tmp
      & (~(weight_mem_run_1_if_for_if_and_stg_2_5_15_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_2_3_sva_1)));
  assign weight_read_ack_5_lpi_1_dfm_15_mx0 = MUX_s_1_2_2(weight_mem_run_1_if_for_if_and_692_nl,
      weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_229_tmp, or_dcpl_34);
  assign weight_mem_run_1_if_for_if_and_696_nl = weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_227_tmp
      & (~(weight_mem_run_1_if_for_if_and_stg_2_3_15_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_2_3_sva_1)));
  assign weight_read_ack_3_lpi_1_dfm_15_mx0 = MUX_s_1_2_2(weight_mem_run_1_if_for_if_and_696_nl,
      weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_227_tmp, or_dcpl_34);
  assign weight_mem_run_1_if_for_if_and_700_nl = weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_225_tmp
      & (~(weight_mem_run_1_if_for_if_and_stg_2_1_15_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_2_3_sva_1)));
  assign weight_read_ack_1_lpi_1_dfm_15_mx0 = MUX_s_1_2_2(weight_mem_run_1_if_for_if_and_700_nl,
      weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_225_tmp, or_dcpl_34);
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_239_tmp = (~ pe_config_is_cluster_sva)
      & PECore_RunFSM_switch_lp_equal_tmp_5 & (nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_14
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_14) & (~(weight_mem_run_1_if_for_if_and_stg_2_7_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_1_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_7_1_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_2_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_7_2_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_3_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_7_3_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_4_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_7_4_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_5_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_7_5_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_6_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_7_6_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_7_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_7_7_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_8_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_7_8_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_9_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_7_9_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_10_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_7_10_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_11_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_7_11_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_12_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_7_12_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_13_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_7_13_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_14_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_7_14_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_15_lpi_1_dfm_1));
  assign weight_mem_run_1_if_for_if_and_stg_2_7_15_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_15_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_2_2_sva_1;
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_238_tmp = (~ pe_config_is_cluster_sva)
      & PECore_RunFSM_switch_lp_equal_tmp_5 & (nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_13
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_13) & (~(weight_mem_run_1_if_for_if_and_stg_2_6_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_1_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_6_1_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_2_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_6_2_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_3_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_6_3_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_4_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_6_4_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_5_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_6_5_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_6_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_6_6_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_7_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_6_7_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_8_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_6_8_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_9_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_6_9_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_10_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_6_10_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_11_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_6_11_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_12_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_6_12_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_13_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_6_13_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_14_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_6_14_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_15_lpi_1_dfm_1));
  assign weight_mem_run_1_if_for_if_and_stg_2_6_15_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_15_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_2_2_sva_1;
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_237_tmp = (~ pe_config_is_cluster_sva)
      & PECore_RunFSM_switch_lp_equal_tmp_5 & (nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_12
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_12) & (~(weight_mem_run_1_if_for_if_and_stg_2_5_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_1_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_5_1_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_2_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_5_2_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_3_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_5_3_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_4_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_5_4_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_5_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_5_5_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_6_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_5_6_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_7_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_5_7_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_8_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_5_8_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_9_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_5_9_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_10_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_5_10_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_11_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_5_11_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_12_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_5_12_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_13_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_5_13_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_14_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_5_14_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_15_lpi_1_dfm_1));
  assign weight_mem_run_1_if_for_if_and_stg_2_5_15_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_15_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_2_2_sva_1;
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_236_tmp = (~ pe_config_is_cluster_sva)
      & PECore_RunFSM_switch_lp_equal_tmp_5 & (nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_11
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_11) & (~(weight_mem_run_1_if_for_if_and_stg_2_4_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_1_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_4_1_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_2_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_4_2_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_3_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_4_3_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_4_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_4_4_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_5_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_4_5_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_6_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_4_6_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_7_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_4_7_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_8_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_4_8_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_9_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_4_9_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_10_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_4_10_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_11_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_4_11_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_12_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_4_12_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_13_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_4_13_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_14_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_4_14_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_15_lpi_1_dfm_1));
  assign weight_mem_run_1_if_for_if_and_stg_2_4_15_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_0_15_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_2_2_sva_1;
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_235_tmp = (~ pe_config_is_cluster_sva)
      & PECore_RunFSM_switch_lp_equal_tmp_5 & (nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_10
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_10) & (~(weight_mem_run_1_if_for_if_and_stg_2_3_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_1_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_3_1_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_2_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_3_2_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_3_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_3_3_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_4_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_3_4_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_5_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_3_5_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_6_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_3_6_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_7_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_3_7_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_8_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_3_8_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_9_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_3_9_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_10_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_3_10_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_11_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_3_11_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_12_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_3_12_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_13_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_3_13_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_14_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_3_14_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_15_lpi_1_dfm_1));
  assign weight_mem_run_1_if_for_if_and_stg_2_3_15_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_3_15_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_2_2_sva_1);
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_234_tmp = (~ pe_config_is_cluster_sva)
      & PECore_RunFSM_switch_lp_equal_tmp_5 & (nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_9
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_9) & (~(weight_mem_run_1_if_for_if_and_stg_2_2_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_1_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_2_1_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_2_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_2_2_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_3_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_2_3_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_4_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_2_4_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_5_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_2_5_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_6_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_2_6_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_7_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_2_7_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_8_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_2_8_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_9_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_2_9_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_10_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_2_10_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_11_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_2_11_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_12_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_2_12_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_13_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_2_13_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_14_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_2_14_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_15_lpi_1_dfm_1));
  assign weight_mem_run_1_if_for_if_and_stg_2_2_15_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_2_15_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_2_2_sva_1);
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_232_tmp = (~ pe_config_is_cluster_sva)
      & PECore_RunFSM_switch_lp_equal_tmp_5 & (nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_7
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_7) & (~(weight_mem_run_1_if_for_if_and_stg_2_0_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_1_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_0_1_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_2_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_0_2_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_3_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_0_3_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_4_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_0_4_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_5_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_0_5_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_6_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_0_6_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_7_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_0_7_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_8_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_0_8_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_9_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_0_9_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_10_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_0_10_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_11_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_0_11_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_12_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_0_12_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_13_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_0_13_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_14_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_0_14_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_15_lpi_1_dfm_1));
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_231_tmp = PECore_RunFSM_switch_lp_equal_tmp_5
      & (nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_6
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_6) & (~(weight_mem_run_1_if_for_if_and_stg_2_7_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_1_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_7_1_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_2_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_7_2_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_3_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_7_3_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_4_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_7_4_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_5_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_7_5_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_6_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_7_6_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_7_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_7_7_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_8_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_7_8_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_9_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_7_9_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_10_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_7_10_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_11_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_7_11_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_12_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_7_12_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_13_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_7_13_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_14_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_7_14_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_15_lpi_1_dfm_1));
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_230_tmp = PECore_RunFSM_switch_lp_equal_tmp_5
      & (nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_5
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_5) & (~(weight_mem_run_1_if_for_if_and_stg_2_6_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_1_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_6_1_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_2_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_6_2_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_3_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_6_3_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_4_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_6_4_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_5_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_6_5_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_6_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_6_6_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_7_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_6_7_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_8_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_6_8_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_9_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_6_9_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_10_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_6_10_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_11_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_6_11_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_12_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_6_12_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_13_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_6_13_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_14_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_6_14_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_15_lpi_1_dfm_1));
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_229_tmp = PECore_RunFSM_switch_lp_equal_tmp_5
      & (nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_4
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_4) & (~(weight_mem_run_1_if_for_if_and_stg_2_5_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_1_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_5_1_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_2_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_5_2_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_3_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_5_3_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_4_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_5_4_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_5_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_5_5_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_6_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_5_6_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_7_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_5_7_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_8_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_5_8_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_9_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_5_9_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_10_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_5_10_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_11_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_5_11_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_12_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_5_12_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_13_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_5_13_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_14_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_5_14_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_15_lpi_1_dfm_1));
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_228_tmp = PECore_RunFSM_switch_lp_equal_tmp_5
      & (nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_3
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_3) & (~(weight_mem_run_1_if_for_if_and_stg_2_4_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_1_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_4_1_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_2_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_4_2_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_3_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_4_3_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_4_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_4_4_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_5_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_4_5_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_6_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_4_6_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_7_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_4_7_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_8_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_4_8_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_9_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_4_9_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_10_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_4_10_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_11_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_4_11_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_12_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_4_12_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_13_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_4_13_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_14_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_4_14_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_15_lpi_1_dfm_1));
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_227_tmp = PECore_RunFSM_switch_lp_equal_tmp_5
      & (nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_2
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_2) & (~(weight_mem_run_1_if_for_if_and_stg_2_3_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_1_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_3_1_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_2_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_3_2_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_3_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_3_3_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_4_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_3_4_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_5_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_3_5_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_6_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_3_6_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_7_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_3_7_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_8_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_3_8_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_9_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_3_9_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_10_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_3_10_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_11_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_3_11_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_12_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_3_12_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_13_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_3_13_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_14_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_3_14_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_15_lpi_1_dfm_1));
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_226_tmp = PECore_RunFSM_switch_lp_equal_tmp_5
      & (nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_1
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_1) & (~(weight_mem_run_1_if_for_if_and_stg_2_2_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_1_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_2_1_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_2_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_2_2_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_3_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_2_3_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_4_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_2_4_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_5_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_2_5_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_6_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_2_6_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_7_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_2_7_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_8_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_2_8_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_9_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_2_9_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_10_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_2_10_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_11_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_2_11_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_12_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_2_12_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_13_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_2_13_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_14_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_2_14_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_15_lpi_1_dfm_1));
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_225_tmp = PECore_RunFSM_switch_lp_equal_tmp_5
      & (Arbiter_16U_Roundrobin_pick_return_15_1_1_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_15_1_2_lpi_1_dfm_3_0
      | Arbiter_16U_Roundrobin_pick_return_15_1_3_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_15_1_4_lpi_1_dfm_3_0
      | Arbiter_16U_Roundrobin_pick_return_15_1_5_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_15_1_6_lpi_1_dfm_3_0
      | Arbiter_16U_Roundrobin_pick_return_15_1_7_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_15_1_8_lpi_1_dfm_3_0
      | Arbiter_16U_Roundrobin_pick_return_15_1_9_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_15_1_10_lpi_1_dfm_3_0
      | Arbiter_16U_Roundrobin_pick_return_15_1_11_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_15_1_12_lpi_1_dfm_3_0
      | Arbiter_16U_Roundrobin_pick_return_15_1_13_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_15_1_14_lpi_1_dfm_3_0
      | Arbiter_16U_Roundrobin_pick_return_15_1_15_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_0)
      & (~(weight_mem_run_1_if_for_if_and_stg_2_1_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_1_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_1_1_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_2_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_1_2_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_3_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_1_3_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_4_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_1_4_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_5_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_1_5_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm_mx1) & weight_mem_run_1_if_for_land_6_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_1_6_sva_1 & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm_mx1)
      & weight_mem_run_1_if_for_land_7_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_1_7_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_8_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_1_8_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_9_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_1_9_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_10_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_1_10_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_11_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_1_11_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_12_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_1_12_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_13_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_1_13_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_14_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_1_14_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm_mx1) &
      weight_mem_run_1_if_for_land_15_lpi_1_dfm_1));
  assign weight_mem_run_1_if_for_if_and_stg_2_1_15_sva_1 = weight_mem_run_1_if_for_if_and_stg_1_1_15_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_2_2_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_0_15_sva_1 = ~(weight_mem_read_arbxbar_xbar_for_3_source_local_2_0_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_source_local_2_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_1_15_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_2_0_sva_1
      & (~ weight_mem_read_arbxbar_xbar_for_3_source_local_2_1_sva_1);
  assign weight_mem_run_1_if_for_if_and_stg_1_2_15_sva_1 = (~ weight_mem_read_arbxbar_xbar_for_3_source_local_2_0_sva_1)
      & weight_mem_read_arbxbar_xbar_for_3_source_local_2_1_sva_1;
  assign weight_mem_run_1_if_for_if_and_stg_1_3_15_sva_1 = weight_mem_read_arbxbar_xbar_for_3_source_local_2_0_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_2_1_sva_1;
  assign weight_write_addrs_lpi_1_dfm_6 = (rva_in_PopNB_mioi_idat_mxwt[147:132])
      & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
      & (signext_16_1(rva_in_PopNB_mioi_idat_mxwt[168])) & ({{15{rva_in_PopNB_mioi_ivld_mxwt}},
      rva_in_PopNB_mioi_ivld_mxwt}) & (signext_16_1(~ is_start_sva));
  assign weight_mem_read_arbxbar_xbar_for_3_1_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_1
      | Arbiter_16U_Roundrobin_pick_return_15_1_1_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_0_1_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_for_3_2_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_1
      | Arbiter_16U_Roundrobin_pick_return_15_1_2_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_0_2_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_for_3_3_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_1
      | Arbiter_16U_Roundrobin_pick_return_15_1_3_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_0_3_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_for_3_4_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_1
      | Arbiter_16U_Roundrobin_pick_return_15_1_4_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_0_4_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_for_3_5_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_1
      | Arbiter_16U_Roundrobin_pick_return_15_1_5_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_0_5_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_for_3_6_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_1
      | Arbiter_16U_Roundrobin_pick_return_15_1_6_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_0_6_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_for_3_7_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_1
      | Arbiter_16U_Roundrobin_pick_return_15_1_7_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_0_7_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_for_3_8_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_1
      | Arbiter_16U_Roundrobin_pick_return_15_1_8_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_0_8_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_for_3_9_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_1
      | Arbiter_16U_Roundrobin_pick_return_15_1_9_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_0_9_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_for_3_10_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_1
      | Arbiter_16U_Roundrobin_pick_return_15_1_10_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_0_10_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_for_3_11_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_1
      | Arbiter_16U_Roundrobin_pick_return_15_1_11_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_0_11_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_for_3_12_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_1
      | Arbiter_16U_Roundrobin_pick_return_15_1_12_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_0_12_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_for_3_13_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_1
      | Arbiter_16U_Roundrobin_pick_return_15_1_13_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_0_13_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_for_3_14_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_1
      | Arbiter_16U_Roundrobin_pick_return_15_1_14_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_0_14_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_for_3_15_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_13
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_12
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_11
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_10
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_9
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_7
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_6
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_5
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_4
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_3
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_2
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_1
      | Arbiter_16U_Roundrobin_pick_return_15_1_15_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_0_15_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_for_3_16_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      = Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_14 | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_13
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_12 | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_11
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_10 | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_9
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_8 | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_7
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_6 | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_5
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_4 | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_3
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_2 | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_1
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_0 | Arbiter_16U_Roundrobin_pick_return_0_lpi_1_dfm_2;
  assign PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_54_nl
      = MUX_s_1_2_2((rva_in_PopNB_mioi_idat_mxwt[8]), pe_config_is_zero_first_sva,
      PECore_DecodeAxiWrite_case_4_switch_lp_or_6_cse_1);
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_56_nl
      = MUX_s_1_2_2(pe_config_is_zero_first_sva, PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_54_nl,
      PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_31);
  assign PECore_DecodeAxi_if_mux_135_nl = MUX_s_1_2_2(pe_config_is_zero_first_sva,
      PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_56_nl,
      rva_in_PopNB_mioi_idat_mxwt[168]);
  assign PECore_DecodeAxi_mux_149_nl = MUX_s_1_2_2(pe_config_is_zero_first_sva, PECore_DecodeAxi_if_mux_135_nl,
      rva_in_PopNB_mioi_ivld_mxwt);
  assign pe_config_is_zero_first_sva_dfm_4_mx0 = MUX_s_1_2_2(PECore_DecodeAxi_mux_149_nl,
      pe_config_is_zero_first_sva, is_start_sva);
  assign pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_pe_config_UpdateInputCounter_if_nor_svs_1
      = ~((pe_config_input_counter_sva_dfm_4_mx0 != (operator_16_false_acc_tmp[7:0]))
      | (operator_16_false_acc_tmp[8]));
  assign PECore_UpdateFSM_switch_lp_or_nl = (~(or_dcpl_306 | pe_config_manager_counter_sva_dfm_4_mx0_0))
      | ((~ or_dcpl_310) & pe_config_manager_counter_sva_dfm_4_mx0_0);
  assign PECore_UpdateFSM_switch_lp_and_2_nl = or_dcpl_306 & (~ pe_config_manager_counter_sva_dfm_4_mx0_0);
  assign PECore_UpdateFSM_switch_lp_and_3_nl = or_dcpl_310 & pe_config_manager_counter_sva_dfm_4_mx0_0;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_mux1h_nl = MUX1HOT_v_8_3_2((rva_in_PopNB_mio_mrgout_dat_sva_1[39:32]),
      pe_manager_num_input_0_sva, pe_manager_num_input_1_sva, {PECore_UpdateFSM_switch_lp_or_nl
      , PECore_UpdateFSM_switch_lp_and_2_nl , PECore_UpdateFSM_switch_lp_and_3_nl});
  assign nl_operator_16_false_acc_tmp = conv_u2s_8_9(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_mux1h_nl)
      + 9'b111111111;
  assign operator_16_false_acc_tmp = nl_operator_16_false_acc_tmp[8:0];
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1
      = ~((pe_config_output_counter_sva_dfm_4_mx0 != (operator_8_false_acc_tmp[7:0]))
      | (operator_8_false_acc_tmp[8]));
  assign pe_config_UpdateManagerCounter_if_unequal_tmp = pe_config_manager_counter_sva_dfm_4_mx1
      != (operator_4_false_acc_tmp[3:0]);
  assign pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_nor_svs_1
      = ~(pe_config_UpdateManagerCounter_if_unequal_tmp | (operator_4_false_acc_tmp[4]));
  assign PECore_UpdateFSM_switch_lp_nor_6_cse = ~(state_2_0_sva_1 | state_2_0_sva_0);
  assign PECore_UpdateFSM_switch_lp_unequal_tmp_1 = ~(state_2_0_sva_2 & PECore_UpdateFSM_switch_lp_nor_6_cse);
  assign PECore_DecodeAxi_if_mux_68_nl = MUX_v_8_2_2((rva_in_PopNB_mio_mrgout_dat_sva_1[47:40]),
      pe_config_num_output_sva, or_dcpl_334);
  assign nl_operator_8_false_acc_tmp = conv_u2s_8_9(PECore_DecodeAxi_if_mux_68_nl)
      + 9'b111111111;
  assign operator_8_false_acc_tmp = nl_operator_8_false_acc_tmp[8:0];
  assign PECore_DecodeAxi_if_mux_69_nl = MUX_v_4_2_2((rva_in_PopNB_mio_mrgout_dat_sva_1[35:32]),
      pe_config_num_manager_sva, or_dcpl_334);
  assign nl_operator_4_false_acc_tmp = conv_u2s_4_5(PECore_DecodeAxi_if_mux_69_nl)
      + 5'b11111;
  assign operator_4_false_acc_tmp = nl_operator_4_false_acc_tmp[4:0];
  assign weight_mem_read_arbxbar_xbar_for_3_1_operator_31_false_operator_31_false_operator_31_false_or_seb
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[0]);
  assign Arbiter_16U_Roundrobin_pick_return_15_1_1_lpi_1_dfm_3_0 = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_0
      & weight_mem_read_arbxbar_xbar_for_3_1_operator_31_false_operator_31_false_operator_31_false_or_seb;
  assign weight_mem_read_arbxbar_xbar_for_3_2_operator_31_false_operator_31_false_operator_31_false_or_seb
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[1]);
  assign Arbiter_16U_Roundrobin_pick_return_15_1_2_lpi_1_dfm_3_0 = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_0
      & weight_mem_read_arbxbar_xbar_for_3_2_operator_31_false_operator_31_false_operator_31_false_or_seb;
  assign weight_mem_read_arbxbar_xbar_for_3_3_operator_31_false_operator_31_false_operator_31_false_or_seb
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[2]);
  assign Arbiter_16U_Roundrobin_pick_return_15_1_3_lpi_1_dfm_3_0 = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_0
      & weight_mem_read_arbxbar_xbar_for_3_3_operator_31_false_operator_31_false_operator_31_false_or_seb;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_4_lpi_1_dfm_3_0 = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_0
      & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_3_tmp;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_5_lpi_1_dfm_3_0 = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_0
      & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_4_tmp;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_6_lpi_1_dfm_3_0 = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_0
      & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_5_tmp;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_7_lpi_1_dfm_3_0 = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_0
      & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_6_tmp;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_8_lpi_1_dfm_3_0 = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_0
      & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_7_tmp;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_9_lpi_1_dfm_3_0 = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_0
      & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_8_tmp;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_10_lpi_1_dfm_3_0 = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_0
      & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_9_tmp;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_11_lpi_1_dfm_3_0 = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_0
      & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_10_tmp;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_12_lpi_1_dfm_3_0 = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_0
      & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_11_tmp;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_13_lpi_1_dfm_3_0 = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_0
      & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_12_tmp;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_14_lpi_1_dfm_3_0 = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_0
      & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_13_tmp;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_15_lpi_1_dfm_3_0 = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_0
      & Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_14_tmp;
  assign weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse
      = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[15])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[15])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[15])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[15])
      | (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[15])
      | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[15])
      | (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[15])
      | (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[15]);
  assign Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_14 = weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_itm
      & weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_13 = weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_1_itm
      & weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_12 = weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_2_itm
      & weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_11 = weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_3_itm
      & weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_10 = weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_4_itm
      & weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_9 = weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_5_itm
      & weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_8 = weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_6_itm
      & weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_7 = weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_7_itm
      & weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_6 = weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_8_itm
      & weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_5 = weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_9_itm
      & weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_4 = weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_10_itm
      & weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_3 = weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_11_itm
      & weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_2 = weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_12_itm
      & weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_1 = weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_13_itm
      & weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse;
  assign Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_0 = weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_14_itm
      & weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse;
  assign Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_14_tmp
      = (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[14])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[14])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[14])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[14])
      | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[14])
      | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[14])
      | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[14])
      | (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[14]);
  assign Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_13_tmp
      = (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[13])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[13])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[13])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[13])
      | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[13])
      | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[13])
      | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[13])
      | (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[13]);
  assign Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_12_tmp
      = (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[12])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[12])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[12])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[12])
      | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[12])
      | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[12])
      | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[12])
      | (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[12]);
  assign Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_11_tmp
      = (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[11])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[11])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[11])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[11])
      | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[11])
      | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[11])
      | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[11])
      | (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[11]);
  assign Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_10_tmp
      = (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[10])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[10])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[10])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[10])
      | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[10])
      | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[10])
      | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[10])
      | (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[10]);
  assign Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_9_tmp
      = (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[9])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[9])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[9])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[9])
      | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[9])
      | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[9])
      | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[9])
      | (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[9]);
  assign Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_8_tmp
      = (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[8])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[8])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[8])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[8])
      | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[8])
      | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[8])
      | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[8])
      | (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[8]);
  assign Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_7_tmp
      = (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]);
  assign Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_6_tmp
      = (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]);
  assign Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_5_tmp
      = (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]);
  assign Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_4_tmp
      = (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]);
  assign Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_3_tmp
      = (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_9_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_for_8_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_7_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_for_6_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_5_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_for_4_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_3_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_for_2_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]);
  assign weight_read_req_valid_8_lpi_1_dfm_1 = (~ pe_config_is_cluster_sva) & PECore_RunFSM_switch_lp_equal_tmp_5;
  assign weight_read_addrs_10_0_lpi_1_dfm_2 = (weight_read_addrs_8_2_0_lpi_1_dfm_1[0])
      & PECore_RunFSM_switch_lp_equal_tmp_5;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_2;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_3;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_4;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_5;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_6;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_7;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_8;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_9;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_10;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_11;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_12;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_13;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_2;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_3;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_4;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_5;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_6;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_7;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_8;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_9;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_10;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_11;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_12;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_13;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_2;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_3;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_4;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_5;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_6;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_7;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_8;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_9;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_10;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_11;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_12;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_13;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_2;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_3;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_4;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_5;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_6;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_7;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_8;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_9;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_10;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_11;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_12;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_13;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_2;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_3;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_4;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_5;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_6;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_7;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_8;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_9;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_10;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_11;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_12;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_13;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_2;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_3;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_4;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_5;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_6;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_7;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_8;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_9;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_10;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_11;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_12;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_13;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_2;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_3;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_4;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_5;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_6;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_7;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_8;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_9;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_10;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_11;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_12;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_13;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_2;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_3;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_4;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_5;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_6;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_7;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_8;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_9;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_10;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_11;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_12;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_13;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_2;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_3;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_4;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_5;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_6;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_7;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_8;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_9;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_10;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_11;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_12;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_13;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_2;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_3;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_4;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_5;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_6;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_7;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_8;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_9;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_10;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_11;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_12;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_13;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_2;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_3;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_4;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_5;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_6;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_7;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_8;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_9;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_10;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_11;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_12;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_13;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_2;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_3;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_4;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_5;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_6;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_7;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_8;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_9;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_10;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_11;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_12;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_13;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_2;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_3;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_4;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_5;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_6;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_7;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_8;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_9;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_10;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_11;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_12;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_13;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_2;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_3;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_4;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_5;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_6;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_7;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_8;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_9;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_10;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_11;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_12;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_13;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_2;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_3;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_4;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_5;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_6;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_7;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_8;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_9;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_10;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_11;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_12;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
      = nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_14
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_13;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_12_itm;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_11_itm;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_10_itm;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_9_itm;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_8_itm;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_7_itm;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_6_itm;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_5_itm;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_4_itm;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_3_itm;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      = Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      | weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_2_itm;
  assign Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      = weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_itm
      | weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_1_itm;
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_10_lpi_1_dfm_1 = MUX_v_4_2_2(4'b0000,
      (weight_read_addrs_9_lpi_1_dfm_3[3:0]), weight_read_ack_9_lpi_1_dfm_15_mx0);
  assign weight_mem_run_1_if_for_if_and_691_nl = weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_233_tmp
      & (~(weight_mem_run_1_if_for_if_and_stg_2_1_15_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_2_3_sva_1));
  assign weight_read_ack_9_lpi_1_dfm_15_mx0 = MUX_s_1_2_2(weight_mem_run_1_if_for_if_and_691_nl,
      weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_233_tmp, or_dcpl_34);
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_233_tmp = (~ pe_config_is_cluster_sva)
      & PECore_RunFSM_switch_lp_equal_tmp_5 & (nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_8
      | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_8
      | Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_8) & (~(weight_mem_run_1_if_for_if_and_stg_2_1_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_1_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_1_1_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_2_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_1_2_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_3_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_1_3_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_4_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_1_4_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_5_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_1_5_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_6_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_1_6_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_7_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_1_7_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_8_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_1_8_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_9_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_1_9_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_10_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_1_10_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_11_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_1_11_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_12_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_1_12_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_13_lpi_1_dfm_1))
      & (~(weight_mem_run_1_if_for_if_and_stg_2_1_13_sva_1 & weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm_mx1
      & weight_mem_run_1_if_for_land_14_lpi_1_dfm_1)) & (~(weight_mem_run_1_if_for_if_and_stg_2_1_14_sva_1
      & weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm_mx1 & weight_mem_run_1_if_for_land_15_lpi_1_dfm_1));
  assign Arbiter_16U_Roundrobin_pick_if_1_not_241 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_14_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_14_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_14_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_14_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_not_243 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_not_245 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_6_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_not_247 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_not_249 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_2_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_not_251 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_1_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_not_253 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_10_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_10_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_10_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_10_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_not_255 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_15_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_15_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_15_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_15_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_not_257 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_5_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_not_259 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_4_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_not_261 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_8_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_8_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_8_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_8_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_not_263 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_11_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_11_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_11_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_11_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_not_265 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_13_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_13_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_13_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_13_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_not_267 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_9_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_9_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_9_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_9_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_not_269 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_7_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_not_271 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_12_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_12_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_12_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_12_lpi_1_dfm_mx0;
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_31 = (rva_in_PopNB_mioi_idat_mxwt[150])
      & PECore_DecodeAxiRead_switch_lp_nor_2_itm_mx0w0;
  assign PECore_DecodeAxiWrite_case_4_switch_lp_nor_7_tmp = ~((rva_in_PopNB_mioi_idat_mxwt[147:133]!=15'b000000000000000));
  assign PECore_DecodeAxiWrite_case_4_switch_lp_nor_9_tmp = ~((rva_in_PopNB_mioi_idat_mxwt[147])
      | (rva_in_PopNB_mioi_idat_mxwt[146]) | (rva_in_PopNB_mioi_idat_mxwt[145]) |
      (rva_in_PopNB_mioi_idat_mxwt[144]) | (rva_in_PopNB_mioi_idat_mxwt[143]) | (rva_in_PopNB_mioi_idat_mxwt[142])
      | (rva_in_PopNB_mioi_idat_mxwt[141]) | (rva_in_PopNB_mioi_idat_mxwt[140]) |
      (rva_in_PopNB_mioi_idat_mxwt[139]) | (rva_in_PopNB_mioi_idat_mxwt[138]) | (rva_in_PopNB_mioi_idat_mxwt[137])
      | (rva_in_PopNB_mioi_idat_mxwt[136]) | (rva_in_PopNB_mioi_idat_mxwt[135]) |
      (rva_in_PopNB_mioi_idat_mxwt[133]));
  assign PECore_DecodeAxiWrite_case_4_switch_lp_nor_11_tmp = ~((rva_in_PopNB_mioi_idat_mxwt[147])
      | (rva_in_PopNB_mioi_idat_mxwt[146]) | (rva_in_PopNB_mioi_idat_mxwt[145]) |
      (rva_in_PopNB_mioi_idat_mxwt[144]) | (rva_in_PopNB_mioi_idat_mxwt[143]) | (rva_in_PopNB_mioi_idat_mxwt[142])
      | (rva_in_PopNB_mioi_idat_mxwt[141]) | (rva_in_PopNB_mioi_idat_mxwt[140]) |
      (rva_in_PopNB_mioi_idat_mxwt[139]) | (rva_in_PopNB_mioi_idat_mxwt[138]) | (rva_in_PopNB_mioi_idat_mxwt[137])
      | (rva_in_PopNB_mioi_idat_mxwt[136]) | (rva_in_PopNB_mioi_idat_mxwt[135]) |
      (rva_in_PopNB_mioi_idat_mxwt[133]) | (rva_in_PopNB_mioi_idat_mxwt[132]));
  assign PECore_DecodeAxiWrite_case_4_switch_lp_nor_13_tmp = ~((rva_in_PopNB_mioi_idat_mxwt[147:134]!=14'b00000000000000));
  assign PECore_DecodeAxiWrite_case_4_switch_lp_nor_15_tmp = ~((rva_in_PopNB_mioi_idat_mxwt[147])
      | (rva_in_PopNB_mioi_idat_mxwt[146]) | (rva_in_PopNB_mioi_idat_mxwt[145]) |
      (rva_in_PopNB_mioi_idat_mxwt[144]) | (rva_in_PopNB_mioi_idat_mxwt[143]) | (rva_in_PopNB_mioi_idat_mxwt[142])
      | (rva_in_PopNB_mioi_idat_mxwt[141]) | (rva_in_PopNB_mioi_idat_mxwt[140]) |
      (rva_in_PopNB_mioi_idat_mxwt[139]) | (rva_in_PopNB_mioi_idat_mxwt[138]) | (rva_in_PopNB_mioi_idat_mxwt[137])
      | (rva_in_PopNB_mioi_idat_mxwt[136]) | (rva_in_PopNB_mioi_idat_mxwt[135]) |
      (rva_in_PopNB_mioi_idat_mxwt[134]) | (rva_in_PopNB_mioi_idat_mxwt[132]));
  assign nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_1_sva_mx0w2 = conv_u2u_3_4(input_mem_banks_write_if_for_if_mux_cse[6:4])
      + conv_u2u_3_4(PECore_RunBias_if_for_if_bias_tmp2_mux_17);
  assign adpfloat_tmp_to_fixed_20U_14U_acc_sdt_1_sva_mx0w2 = nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_1_sva_mx0w2[3:0];
  assign nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_12_sva_mx0w1 = conv_u2u_3_4(input_mem_banks_write_if_for_if_mux_cse[94:92])
      + conv_u2u_3_4(PECore_RunBias_if_for_if_bias_tmp2_mux_17);
  assign adpfloat_tmp_to_fixed_20U_14U_acc_sdt_12_sva_mx0w1 = nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_12_sva_mx0w1[3:0];
  assign nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_2_sva_mx0w1 = conv_u2u_3_4(input_mem_banks_write_if_for_if_mux_cse[14:12])
      + conv_u2u_3_4(PECore_RunBias_if_for_if_bias_tmp2_mux_17);
  assign adpfloat_tmp_to_fixed_20U_14U_acc_sdt_2_sva_mx0w1 = nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_2_sva_mx0w1[3:0];
  assign nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_3_sva_mx0w1 = conv_u2u_3_4(input_mem_banks_write_if_for_if_mux_cse[22:20])
      + conv_u2u_3_4(PECore_RunBias_if_for_if_bias_tmp2_mux_17);
  assign adpfloat_tmp_to_fixed_20U_14U_acc_sdt_3_sva_mx0w1 = nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_3_sva_mx0w1[3:0];
  assign nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_4_sva_mx0w1 = conv_u2u_3_4(input_mem_banks_write_if_for_if_mux_cse[30:28])
      + conv_u2u_3_4(PECore_RunBias_if_for_if_bias_tmp2_mux_17);
  assign adpfloat_tmp_to_fixed_20U_14U_acc_sdt_4_sva_mx0w1 = nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_4_sva_mx0w1[3:0];
  assign nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_5_sva_mx0w1 = conv_u2u_3_4(input_mem_banks_write_if_for_if_mux_cse[38:36])
      + conv_u2u_3_4(PECore_RunBias_if_for_if_bias_tmp2_mux_17);
  assign adpfloat_tmp_to_fixed_20U_14U_acc_sdt_5_sva_mx0w1 = nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_5_sva_mx0w1[3:0];
  assign nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_8_sva_mx0w1 = conv_u2u_3_4(input_mem_banks_write_if_for_if_mux_cse[62:60])
      + conv_u2u_3_4(PECore_RunBias_if_for_if_bias_tmp2_mux_17);
  assign adpfloat_tmp_to_fixed_20U_14U_acc_sdt_8_sva_mx0w1 = nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_8_sva_mx0w1[3:0];
  assign nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_9_sva_mx0w1 = conv_u2u_3_4(input_mem_banks_write_if_for_if_mux_cse[70:68])
      + conv_u2u_3_4(PECore_RunBias_if_for_if_bias_tmp2_mux_17);
  assign adpfloat_tmp_to_fixed_20U_14U_acc_sdt_9_sva_mx0w1 = nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_9_sva_mx0w1[3:0];
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_12_mx1w2
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_2_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_2_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_123_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_11_mx1w2
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_3_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_3_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_123_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_13_mx1w2
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_1_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_1_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_123_ftd_1);
  assign rva_out_reg_data_and_2_cse = crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm
      & (fsm_output[2]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_0_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_0_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_130_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_1_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_1_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_130_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_2_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_2_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_130_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_3_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_3_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_130_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_4_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_4_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_130_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_5_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_5_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_130_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_6_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_6_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_130_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_7_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_7_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_130_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_8_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_8_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_130_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_9_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_9_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_130_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_10_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_10_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_130_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_11_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_11_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_130_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_12_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_12_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_130_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_13_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_13_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_130_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_14_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_14_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_130_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_15_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_15_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_130_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm});
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_260_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[0]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_0_0_lpi_1_dfm_2 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data0_rsci_q_d[7:0]), weight_mem_write_arbxbar_xbar_for_1_for_not_260_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_262_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[1]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_1_0_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data1_rsci_q_d[7:0]), weight_mem_write_arbxbar_xbar_for_1_for_not_262_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_264_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[2]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_2_0_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data2_rsci_q_d[7:0]), weight_mem_write_arbxbar_xbar_for_1_for_not_264_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_266_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[3]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_3_0_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data3_rsci_q_d[7:0]), weight_mem_write_arbxbar_xbar_for_1_for_not_266_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_268_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[4]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_4_0_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data4_rsci_q_d[7:0]), weight_mem_write_arbxbar_xbar_for_1_for_not_268_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_270_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[5]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_5_0_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data5_rsci_q_d[7:0]), weight_mem_write_arbxbar_xbar_for_1_for_not_270_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_272_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[6]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_6_0_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data6_rsci_q_d[7:0]), weight_mem_write_arbxbar_xbar_for_1_for_not_272_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_274_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[7]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_7_0_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data7_rsci_q_d[7:0]), weight_mem_write_arbxbar_xbar_for_1_for_not_274_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_276_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[8]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_8_0_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data8_rsci_q_d[7:0]), weight_mem_write_arbxbar_xbar_for_1_for_not_276_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_278_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[9]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_9_0_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data9_rsci_q_d[7:0]), weight_mem_write_arbxbar_xbar_for_1_for_not_278_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_280_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[10]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_10_0_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data10_rsci_q_d[7:0]), weight_mem_write_arbxbar_xbar_for_1_for_not_280_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_282_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[11]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_11_0_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data11_rsci_q_d[7:0]), weight_mem_write_arbxbar_xbar_for_1_for_not_282_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_284_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[12]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_12_0_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data12_rsci_q_d[7:0]), weight_mem_write_arbxbar_xbar_for_1_for_not_284_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_286_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[13]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_13_0_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data13_rsci_q_d[7:0]), weight_mem_write_arbxbar_xbar_for_1_for_not_286_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_256_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[14]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_14_0_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data14_rsci_q_d[7:0]), weight_mem_write_arbxbar_xbar_for_1_for_not_256_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_258_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[15]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_15_0_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data15_rsci_q_d[7:0]), weight_mem_write_arbxbar_xbar_for_1_for_not_258_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_332_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[0]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_0_1_lpi_1_dfm_2 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data0_rsci_q_d[15:8]), weight_mem_write_arbxbar_xbar_for_1_for_not_332_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_347_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[1]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_1_1_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data1_rsci_q_d[15:8]), weight_mem_write_arbxbar_xbar_for_1_for_not_347_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_362_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[2]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_2_1_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data2_rsci_q_d[15:8]), weight_mem_write_arbxbar_xbar_for_1_for_not_362_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_377_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[3]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_3_1_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data3_rsci_q_d[15:8]), weight_mem_write_arbxbar_xbar_for_1_for_not_377_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_392_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[4]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_4_1_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data4_rsci_q_d[15:8]), weight_mem_write_arbxbar_xbar_for_1_for_not_392_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_407_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[5]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_5_1_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data5_rsci_q_d[15:8]), weight_mem_write_arbxbar_xbar_for_1_for_not_407_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_422_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[6]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_6_1_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data6_rsci_q_d[15:8]), weight_mem_write_arbxbar_xbar_for_1_for_not_422_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_437_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[7]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_7_1_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data7_rsci_q_d[15:8]), weight_mem_write_arbxbar_xbar_for_1_for_not_437_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_452_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[8]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_8_1_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data8_rsci_q_d[15:8]), weight_mem_write_arbxbar_xbar_for_1_for_not_452_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_467_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[9]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_9_1_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data9_rsci_q_d[15:8]), weight_mem_write_arbxbar_xbar_for_1_for_not_467_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_482_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[10]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_10_1_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data10_rsci_q_d[15:8]), weight_mem_write_arbxbar_xbar_for_1_for_not_482_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_497_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[11]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_11_1_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data11_rsci_q_d[15:8]), weight_mem_write_arbxbar_xbar_for_1_for_not_497_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_512_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[12]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_12_1_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data12_rsci_q_d[15:8]), weight_mem_write_arbxbar_xbar_for_1_for_not_512_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_527_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[13]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_13_1_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data13_rsci_q_d[15:8]), weight_mem_write_arbxbar_xbar_for_1_for_not_527_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_302_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[14]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_14_1_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data14_rsci_q_d[15:8]), weight_mem_write_arbxbar_xbar_for_1_for_not_302_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_317_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[15]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_15_1_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data15_rsci_q_d[15:8]), weight_mem_write_arbxbar_xbar_for_1_for_not_317_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_331_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[0]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_0_2_lpi_1_dfm_2 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data0_rsci_q_d[23:16]), weight_mem_write_arbxbar_xbar_for_1_for_not_331_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_346_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[1]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_1_2_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data1_rsci_q_d[23:16]), weight_mem_write_arbxbar_xbar_for_1_for_not_346_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_361_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[2]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_2_2_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data2_rsci_q_d[23:16]), weight_mem_write_arbxbar_xbar_for_1_for_not_361_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_376_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[3]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_3_2_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data3_rsci_q_d[23:16]), weight_mem_write_arbxbar_xbar_for_1_for_not_376_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_391_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[4]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_4_2_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data4_rsci_q_d[23:16]), weight_mem_write_arbxbar_xbar_for_1_for_not_391_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_406_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[5]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_5_2_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data5_rsci_q_d[23:16]), weight_mem_write_arbxbar_xbar_for_1_for_not_406_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_421_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[6]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_6_2_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data6_rsci_q_d[23:16]), weight_mem_write_arbxbar_xbar_for_1_for_not_421_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_436_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[7]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_7_2_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data7_rsci_q_d[23:16]), weight_mem_write_arbxbar_xbar_for_1_for_not_436_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_451_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[8]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_8_2_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data8_rsci_q_d[23:16]), weight_mem_write_arbxbar_xbar_for_1_for_not_451_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_466_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[9]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_9_2_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data9_rsci_q_d[23:16]), weight_mem_write_arbxbar_xbar_for_1_for_not_466_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_481_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[10]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_10_2_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data10_rsci_q_d[23:16]), weight_mem_write_arbxbar_xbar_for_1_for_not_481_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_496_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[11]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_11_2_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data11_rsci_q_d[23:16]), weight_mem_write_arbxbar_xbar_for_1_for_not_496_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_511_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[12]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_12_2_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data12_rsci_q_d[23:16]), weight_mem_write_arbxbar_xbar_for_1_for_not_511_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_526_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[13]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_13_2_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data13_rsci_q_d[23:16]), weight_mem_write_arbxbar_xbar_for_1_for_not_526_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_301_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[14]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_14_2_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data14_rsci_q_d[23:16]), weight_mem_write_arbxbar_xbar_for_1_for_not_301_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_316_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[15]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_15_2_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data15_rsci_q_d[23:16]), weight_mem_write_arbxbar_xbar_for_1_for_not_316_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_330_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[0]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_0_3_lpi_1_dfm_2 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data0_rsci_q_d[31:24]), weight_mem_write_arbxbar_xbar_for_1_for_not_330_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_345_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[1]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_1_3_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data1_rsci_q_d[31:24]), weight_mem_write_arbxbar_xbar_for_1_for_not_345_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_360_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[2]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_2_3_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data2_rsci_q_d[31:24]), weight_mem_write_arbxbar_xbar_for_1_for_not_360_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_375_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[3]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_3_3_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data3_rsci_q_d[31:24]), weight_mem_write_arbxbar_xbar_for_1_for_not_375_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_390_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[4]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_4_3_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data4_rsci_q_d[31:24]), weight_mem_write_arbxbar_xbar_for_1_for_not_390_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_405_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[5]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_5_3_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data5_rsci_q_d[31:24]), weight_mem_write_arbxbar_xbar_for_1_for_not_405_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_420_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[6]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_6_3_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data6_rsci_q_d[31:24]), weight_mem_write_arbxbar_xbar_for_1_for_not_420_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_435_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[7]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_7_3_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data7_rsci_q_d[31:24]), weight_mem_write_arbxbar_xbar_for_1_for_not_435_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_450_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[8]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_8_3_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data8_rsci_q_d[31:24]), weight_mem_write_arbxbar_xbar_for_1_for_not_450_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_465_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[9]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_9_3_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data9_rsci_q_d[31:24]), weight_mem_write_arbxbar_xbar_for_1_for_not_465_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_480_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[10]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_10_3_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data10_rsci_q_d[31:24]), weight_mem_write_arbxbar_xbar_for_1_for_not_480_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_495_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[11]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_11_3_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data11_rsci_q_d[31:24]), weight_mem_write_arbxbar_xbar_for_1_for_not_495_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_510_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[12]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_12_3_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data12_rsci_q_d[31:24]), weight_mem_write_arbxbar_xbar_for_1_for_not_510_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_525_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[13]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_13_3_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data13_rsci_q_d[31:24]), weight_mem_write_arbxbar_xbar_for_1_for_not_525_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_300_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[14]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_14_3_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data14_rsci_q_d[31:24]), weight_mem_write_arbxbar_xbar_for_1_for_not_300_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_315_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[15]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_15_3_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data15_rsci_q_d[31:24]), weight_mem_write_arbxbar_xbar_for_1_for_not_315_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_329_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[0]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_0_4_lpi_1_dfm_2 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data0_rsci_q_d[39:32]), weight_mem_write_arbxbar_xbar_for_1_for_not_329_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_344_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[1]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_1_4_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data1_rsci_q_d[39:32]), weight_mem_write_arbxbar_xbar_for_1_for_not_344_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_359_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[2]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_2_4_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data2_rsci_q_d[39:32]), weight_mem_write_arbxbar_xbar_for_1_for_not_359_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_374_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[3]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_3_4_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data3_rsci_q_d[39:32]), weight_mem_write_arbxbar_xbar_for_1_for_not_374_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_389_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[4]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_4_4_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data4_rsci_q_d[39:32]), weight_mem_write_arbxbar_xbar_for_1_for_not_389_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_404_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[5]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_5_4_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data5_rsci_q_d[39:32]), weight_mem_write_arbxbar_xbar_for_1_for_not_404_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_419_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[6]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_6_4_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data6_rsci_q_d[39:32]), weight_mem_write_arbxbar_xbar_for_1_for_not_419_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_434_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[7]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_7_4_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data7_rsci_q_d[39:32]), weight_mem_write_arbxbar_xbar_for_1_for_not_434_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_449_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[8]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_8_4_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data8_rsci_q_d[39:32]), weight_mem_write_arbxbar_xbar_for_1_for_not_449_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_464_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[9]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_9_4_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data9_rsci_q_d[39:32]), weight_mem_write_arbxbar_xbar_for_1_for_not_464_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_479_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[10]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_10_4_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data10_rsci_q_d[39:32]), weight_mem_write_arbxbar_xbar_for_1_for_not_479_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_494_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[11]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_11_4_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data11_rsci_q_d[39:32]), weight_mem_write_arbxbar_xbar_for_1_for_not_494_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_509_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[12]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_12_4_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data12_rsci_q_d[39:32]), weight_mem_write_arbxbar_xbar_for_1_for_not_509_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_524_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[13]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_13_4_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data13_rsci_q_d[39:32]), weight_mem_write_arbxbar_xbar_for_1_for_not_524_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_299_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[14]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_14_4_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data14_rsci_q_d[39:32]), weight_mem_write_arbxbar_xbar_for_1_for_not_299_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_314_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[15]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_15_4_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data15_rsci_q_d[39:32]), weight_mem_write_arbxbar_xbar_for_1_for_not_314_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_328_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[0]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_0_5_lpi_1_dfm_2 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data0_rsci_q_d[47:40]), weight_mem_write_arbxbar_xbar_for_1_for_not_328_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_343_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[1]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_1_5_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data1_rsci_q_d[47:40]), weight_mem_write_arbxbar_xbar_for_1_for_not_343_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_358_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[2]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_2_5_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data2_rsci_q_d[47:40]), weight_mem_write_arbxbar_xbar_for_1_for_not_358_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_373_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[3]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_3_5_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data3_rsci_q_d[47:40]), weight_mem_write_arbxbar_xbar_for_1_for_not_373_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_388_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[4]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_4_5_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data4_rsci_q_d[47:40]), weight_mem_write_arbxbar_xbar_for_1_for_not_388_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_403_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[5]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_5_5_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data5_rsci_q_d[47:40]), weight_mem_write_arbxbar_xbar_for_1_for_not_403_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_418_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[6]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_6_5_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data6_rsci_q_d[47:40]), weight_mem_write_arbxbar_xbar_for_1_for_not_418_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_433_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[7]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_7_5_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data7_rsci_q_d[47:40]), weight_mem_write_arbxbar_xbar_for_1_for_not_433_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_448_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[8]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_8_5_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data8_rsci_q_d[47:40]), weight_mem_write_arbxbar_xbar_for_1_for_not_448_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_463_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[9]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_9_5_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data9_rsci_q_d[47:40]), weight_mem_write_arbxbar_xbar_for_1_for_not_463_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_478_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[10]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_10_5_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data10_rsci_q_d[47:40]), weight_mem_write_arbxbar_xbar_for_1_for_not_478_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_493_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[11]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_11_5_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data11_rsci_q_d[47:40]), weight_mem_write_arbxbar_xbar_for_1_for_not_493_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_508_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[12]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_12_5_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data12_rsci_q_d[47:40]), weight_mem_write_arbxbar_xbar_for_1_for_not_508_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_523_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[13]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_13_5_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data13_rsci_q_d[47:40]), weight_mem_write_arbxbar_xbar_for_1_for_not_523_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_298_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[14]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_14_5_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data14_rsci_q_d[47:40]), weight_mem_write_arbxbar_xbar_for_1_for_not_298_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_313_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[15]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_15_5_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data15_rsci_q_d[47:40]), weight_mem_write_arbxbar_xbar_for_1_for_not_313_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_327_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[0]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_0_6_lpi_1_dfm_2 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data0_rsci_q_d[55:48]), weight_mem_write_arbxbar_xbar_for_1_for_not_327_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_342_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[1]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_1_6_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data1_rsci_q_d[55:48]), weight_mem_write_arbxbar_xbar_for_1_for_not_342_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_357_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[2]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_2_6_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data2_rsci_q_d[55:48]), weight_mem_write_arbxbar_xbar_for_1_for_not_357_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_372_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[3]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_3_6_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data3_rsci_q_d[55:48]), weight_mem_write_arbxbar_xbar_for_1_for_not_372_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_387_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[4]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_4_6_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data4_rsci_q_d[55:48]), weight_mem_write_arbxbar_xbar_for_1_for_not_387_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_402_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[5]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_5_6_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data5_rsci_q_d[55:48]), weight_mem_write_arbxbar_xbar_for_1_for_not_402_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_417_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[6]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_6_6_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data6_rsci_q_d[55:48]), weight_mem_write_arbxbar_xbar_for_1_for_not_417_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_432_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[7]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_7_6_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data7_rsci_q_d[55:48]), weight_mem_write_arbxbar_xbar_for_1_for_not_432_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_447_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[8]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_8_6_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data8_rsci_q_d[55:48]), weight_mem_write_arbxbar_xbar_for_1_for_not_447_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_462_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[9]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_9_6_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data9_rsci_q_d[55:48]), weight_mem_write_arbxbar_xbar_for_1_for_not_462_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_477_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[10]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_10_6_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data10_rsci_q_d[55:48]), weight_mem_write_arbxbar_xbar_for_1_for_not_477_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_492_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[11]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_11_6_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data11_rsci_q_d[55:48]), weight_mem_write_arbxbar_xbar_for_1_for_not_492_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_507_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[12]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_12_6_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data12_rsci_q_d[55:48]), weight_mem_write_arbxbar_xbar_for_1_for_not_507_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_522_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[13]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_13_6_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data13_rsci_q_d[55:48]), weight_mem_write_arbxbar_xbar_for_1_for_not_522_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_297_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[14]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_14_6_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data14_rsci_q_d[55:48]), weight_mem_write_arbxbar_xbar_for_1_for_not_297_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_312_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[15]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_15_6_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data15_rsci_q_d[55:48]), weight_mem_write_arbxbar_xbar_for_1_for_not_312_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_326_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[0]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_0_7_lpi_1_dfm_2 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data0_rsci_q_d[63:56]), weight_mem_write_arbxbar_xbar_for_1_for_not_326_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_341_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[1]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_1_7_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data1_rsci_q_d[63:56]), weight_mem_write_arbxbar_xbar_for_1_for_not_341_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_356_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[2]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_2_7_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data2_rsci_q_d[63:56]), weight_mem_write_arbxbar_xbar_for_1_for_not_356_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_371_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[3]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_3_7_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data3_rsci_q_d[63:56]), weight_mem_write_arbxbar_xbar_for_1_for_not_371_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_386_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[4]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_4_7_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data4_rsci_q_d[63:56]), weight_mem_write_arbxbar_xbar_for_1_for_not_386_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_401_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[5]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_5_7_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data5_rsci_q_d[63:56]), weight_mem_write_arbxbar_xbar_for_1_for_not_401_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_416_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[6]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_6_7_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data6_rsci_q_d[63:56]), weight_mem_write_arbxbar_xbar_for_1_for_not_416_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_431_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[7]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_7_7_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data7_rsci_q_d[63:56]), weight_mem_write_arbxbar_xbar_for_1_for_not_431_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_446_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[8]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_8_7_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data8_rsci_q_d[63:56]), weight_mem_write_arbxbar_xbar_for_1_for_not_446_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_461_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[9]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_9_7_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data9_rsci_q_d[63:56]), weight_mem_write_arbxbar_xbar_for_1_for_not_461_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_476_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[10]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_10_7_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data10_rsci_q_d[63:56]), weight_mem_write_arbxbar_xbar_for_1_for_not_476_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_491_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[11]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_11_7_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data11_rsci_q_d[63:56]), weight_mem_write_arbxbar_xbar_for_1_for_not_491_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_506_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[12]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_12_7_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data12_rsci_q_d[63:56]), weight_mem_write_arbxbar_xbar_for_1_for_not_506_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_521_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[13]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_13_7_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data13_rsci_q_d[63:56]), weight_mem_write_arbxbar_xbar_for_1_for_not_521_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_296_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[14]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_14_7_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data14_rsci_q_d[63:56]), weight_mem_write_arbxbar_xbar_for_1_for_not_296_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_311_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[15]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_15_7_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data15_rsci_q_d[63:56]), weight_mem_write_arbxbar_xbar_for_1_for_not_311_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_325_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[0]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_0_8_lpi_1_dfm_2 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data0_rsci_q_d[71:64]), weight_mem_write_arbxbar_xbar_for_1_for_not_325_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_340_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[1]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_1_8_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data1_rsci_q_d[71:64]), weight_mem_write_arbxbar_xbar_for_1_for_not_340_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_355_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[2]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_2_8_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data2_rsci_q_d[71:64]), weight_mem_write_arbxbar_xbar_for_1_for_not_355_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_370_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[3]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_3_8_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data3_rsci_q_d[71:64]), weight_mem_write_arbxbar_xbar_for_1_for_not_370_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_385_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[4]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_4_8_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data4_rsci_q_d[71:64]), weight_mem_write_arbxbar_xbar_for_1_for_not_385_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_400_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[5]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_5_8_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data5_rsci_q_d[71:64]), weight_mem_write_arbxbar_xbar_for_1_for_not_400_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_415_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[6]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_6_8_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data6_rsci_q_d[71:64]), weight_mem_write_arbxbar_xbar_for_1_for_not_415_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_430_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[7]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_7_8_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data7_rsci_q_d[71:64]), weight_mem_write_arbxbar_xbar_for_1_for_not_430_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_445_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[8]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_8_8_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data8_rsci_q_d[71:64]), weight_mem_write_arbxbar_xbar_for_1_for_not_445_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_460_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[9]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_9_8_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data9_rsci_q_d[71:64]), weight_mem_write_arbxbar_xbar_for_1_for_not_460_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_475_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[10]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_10_8_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data10_rsci_q_d[71:64]), weight_mem_write_arbxbar_xbar_for_1_for_not_475_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_490_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[11]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_11_8_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data11_rsci_q_d[71:64]), weight_mem_write_arbxbar_xbar_for_1_for_not_490_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_505_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[12]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_12_8_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data12_rsci_q_d[71:64]), weight_mem_write_arbxbar_xbar_for_1_for_not_505_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_520_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[13]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_13_8_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data13_rsci_q_d[71:64]), weight_mem_write_arbxbar_xbar_for_1_for_not_520_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_295_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[14]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_14_8_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data14_rsci_q_d[71:64]), weight_mem_write_arbxbar_xbar_for_1_for_not_295_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_310_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[15]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_15_8_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data15_rsci_q_d[71:64]), weight_mem_write_arbxbar_xbar_for_1_for_not_310_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_324_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[0]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_0_9_lpi_1_dfm_2 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data0_rsci_q_d[79:72]), weight_mem_write_arbxbar_xbar_for_1_for_not_324_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_339_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[1]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_1_9_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data1_rsci_q_d[79:72]), weight_mem_write_arbxbar_xbar_for_1_for_not_339_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_354_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[2]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_2_9_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data2_rsci_q_d[79:72]), weight_mem_write_arbxbar_xbar_for_1_for_not_354_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_369_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[3]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_3_9_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data3_rsci_q_d[79:72]), weight_mem_write_arbxbar_xbar_for_1_for_not_369_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_384_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[4]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_4_9_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data4_rsci_q_d[79:72]), weight_mem_write_arbxbar_xbar_for_1_for_not_384_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_399_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[5]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_5_9_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data5_rsci_q_d[79:72]), weight_mem_write_arbxbar_xbar_for_1_for_not_399_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_414_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[6]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_6_9_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data6_rsci_q_d[79:72]), weight_mem_write_arbxbar_xbar_for_1_for_not_414_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_429_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[7]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_7_9_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data7_rsci_q_d[79:72]), weight_mem_write_arbxbar_xbar_for_1_for_not_429_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_444_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[8]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_8_9_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data8_rsci_q_d[79:72]), weight_mem_write_arbxbar_xbar_for_1_for_not_444_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_459_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[9]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_9_9_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data9_rsci_q_d[79:72]), weight_mem_write_arbxbar_xbar_for_1_for_not_459_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_474_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[10]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_10_9_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data10_rsci_q_d[79:72]), weight_mem_write_arbxbar_xbar_for_1_for_not_474_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_489_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[11]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_11_9_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data11_rsci_q_d[79:72]), weight_mem_write_arbxbar_xbar_for_1_for_not_489_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_504_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[12]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_12_9_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data12_rsci_q_d[79:72]), weight_mem_write_arbxbar_xbar_for_1_for_not_504_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_519_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[13]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_13_9_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data13_rsci_q_d[79:72]), weight_mem_write_arbxbar_xbar_for_1_for_not_519_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_294_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[14]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_14_9_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data14_rsci_q_d[79:72]), weight_mem_write_arbxbar_xbar_for_1_for_not_294_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_309_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[15]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_15_9_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data15_rsci_q_d[79:72]), weight_mem_write_arbxbar_xbar_for_1_for_not_309_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_323_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[0]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_0_10_lpi_1_dfm_2 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data0_rsci_q_d[87:80]), weight_mem_write_arbxbar_xbar_for_1_for_not_323_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_338_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[1]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_1_10_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data1_rsci_q_d[87:80]), weight_mem_write_arbxbar_xbar_for_1_for_not_338_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_353_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[2]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_2_10_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data2_rsci_q_d[87:80]), weight_mem_write_arbxbar_xbar_for_1_for_not_353_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_368_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[3]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_3_10_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data3_rsci_q_d[87:80]), weight_mem_write_arbxbar_xbar_for_1_for_not_368_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_383_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[4]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_4_10_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data4_rsci_q_d[87:80]), weight_mem_write_arbxbar_xbar_for_1_for_not_383_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_398_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[5]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_5_10_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data5_rsci_q_d[87:80]), weight_mem_write_arbxbar_xbar_for_1_for_not_398_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_413_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[6]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_6_10_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data6_rsci_q_d[87:80]), weight_mem_write_arbxbar_xbar_for_1_for_not_413_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_428_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[7]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_7_10_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data7_rsci_q_d[87:80]), weight_mem_write_arbxbar_xbar_for_1_for_not_428_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_443_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[8]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_8_10_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data8_rsci_q_d[87:80]), weight_mem_write_arbxbar_xbar_for_1_for_not_443_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_458_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[9]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_9_10_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data9_rsci_q_d[87:80]), weight_mem_write_arbxbar_xbar_for_1_for_not_458_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_473_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[10]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_10_10_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data10_rsci_q_d[87:80]), weight_mem_write_arbxbar_xbar_for_1_for_not_473_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_488_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[11]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_11_10_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data11_rsci_q_d[87:80]), weight_mem_write_arbxbar_xbar_for_1_for_not_488_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_503_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[12]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_12_10_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data12_rsci_q_d[87:80]), weight_mem_write_arbxbar_xbar_for_1_for_not_503_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_518_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[13]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_13_10_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data13_rsci_q_d[87:80]), weight_mem_write_arbxbar_xbar_for_1_for_not_518_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_293_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[14]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_14_10_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data14_rsci_q_d[87:80]), weight_mem_write_arbxbar_xbar_for_1_for_not_293_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_308_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[15]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_15_10_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data15_rsci_q_d[87:80]), weight_mem_write_arbxbar_xbar_for_1_for_not_308_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_322_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[0]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_0_11_lpi_1_dfm_2 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data0_rsci_q_d[95:88]), weight_mem_write_arbxbar_xbar_for_1_for_not_322_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_337_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[1]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_1_11_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data1_rsci_q_d[95:88]), weight_mem_write_arbxbar_xbar_for_1_for_not_337_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_352_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[2]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_2_11_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data2_rsci_q_d[95:88]), weight_mem_write_arbxbar_xbar_for_1_for_not_352_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_367_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[3]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_3_11_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data3_rsci_q_d[95:88]), weight_mem_write_arbxbar_xbar_for_1_for_not_367_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_382_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[4]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_4_11_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data4_rsci_q_d[95:88]), weight_mem_write_arbxbar_xbar_for_1_for_not_382_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_397_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[5]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_5_11_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data5_rsci_q_d[95:88]), weight_mem_write_arbxbar_xbar_for_1_for_not_397_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_412_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[6]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_6_11_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data6_rsci_q_d[95:88]), weight_mem_write_arbxbar_xbar_for_1_for_not_412_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_427_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[7]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_7_11_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data7_rsci_q_d[95:88]), weight_mem_write_arbxbar_xbar_for_1_for_not_427_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_442_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[8]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_8_11_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data8_rsci_q_d[95:88]), weight_mem_write_arbxbar_xbar_for_1_for_not_442_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_457_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[9]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_9_11_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data9_rsci_q_d[95:88]), weight_mem_write_arbxbar_xbar_for_1_for_not_457_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_472_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[10]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_10_11_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data10_rsci_q_d[95:88]), weight_mem_write_arbxbar_xbar_for_1_for_not_472_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_487_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[11]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_11_11_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data11_rsci_q_d[95:88]), weight_mem_write_arbxbar_xbar_for_1_for_not_487_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_502_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[12]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_12_11_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data12_rsci_q_d[95:88]), weight_mem_write_arbxbar_xbar_for_1_for_not_502_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_517_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[13]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_13_11_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data13_rsci_q_d[95:88]), weight_mem_write_arbxbar_xbar_for_1_for_not_517_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_292_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[14]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_14_11_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data14_rsci_q_d[95:88]), weight_mem_write_arbxbar_xbar_for_1_for_not_292_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_307_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[15]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_15_11_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data15_rsci_q_d[95:88]), weight_mem_write_arbxbar_xbar_for_1_for_not_307_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_321_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[0]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_0_12_lpi_1_dfm_2 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data0_rsci_q_d[103:96]), weight_mem_write_arbxbar_xbar_for_1_for_not_321_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_336_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[1]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_1_12_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data1_rsci_q_d[103:96]), weight_mem_write_arbxbar_xbar_for_1_for_not_336_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_351_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[2]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_2_12_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data2_rsci_q_d[103:96]), weight_mem_write_arbxbar_xbar_for_1_for_not_351_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_366_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[3]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_3_12_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data3_rsci_q_d[103:96]), weight_mem_write_arbxbar_xbar_for_1_for_not_366_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_381_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[4]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_4_12_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data4_rsci_q_d[103:96]), weight_mem_write_arbxbar_xbar_for_1_for_not_381_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_396_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[5]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_5_12_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data5_rsci_q_d[103:96]), weight_mem_write_arbxbar_xbar_for_1_for_not_396_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_411_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[6]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_6_12_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data6_rsci_q_d[103:96]), weight_mem_write_arbxbar_xbar_for_1_for_not_411_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_426_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[7]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_7_12_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data7_rsci_q_d[103:96]), weight_mem_write_arbxbar_xbar_for_1_for_not_426_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_441_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[8]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_8_12_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data8_rsci_q_d[103:96]), weight_mem_write_arbxbar_xbar_for_1_for_not_441_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_456_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[9]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_9_12_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data9_rsci_q_d[103:96]), weight_mem_write_arbxbar_xbar_for_1_for_not_456_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_471_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[10]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_10_12_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data10_rsci_q_d[103:96]), weight_mem_write_arbxbar_xbar_for_1_for_not_471_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_486_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[11]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_11_12_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data11_rsci_q_d[103:96]), weight_mem_write_arbxbar_xbar_for_1_for_not_486_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_501_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[12]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_12_12_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data12_rsci_q_d[103:96]), weight_mem_write_arbxbar_xbar_for_1_for_not_501_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_516_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[13]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_13_12_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data13_rsci_q_d[103:96]), weight_mem_write_arbxbar_xbar_for_1_for_not_516_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_291_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[14]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_14_12_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data14_rsci_q_d[103:96]), weight_mem_write_arbxbar_xbar_for_1_for_not_291_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_306_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[15]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_15_12_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data15_rsci_q_d[103:96]), weight_mem_write_arbxbar_xbar_for_1_for_not_306_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_320_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[0]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_0_13_lpi_1_dfm_2 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data0_rsci_q_d[111:104]), weight_mem_write_arbxbar_xbar_for_1_for_not_320_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_335_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[1]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_1_13_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data1_rsci_q_d[111:104]), weight_mem_write_arbxbar_xbar_for_1_for_not_335_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_350_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[2]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_2_13_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data2_rsci_q_d[111:104]), weight_mem_write_arbxbar_xbar_for_1_for_not_350_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_365_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[3]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_3_13_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data3_rsci_q_d[111:104]), weight_mem_write_arbxbar_xbar_for_1_for_not_365_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_380_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[4]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_4_13_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data4_rsci_q_d[111:104]), weight_mem_write_arbxbar_xbar_for_1_for_not_380_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_395_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[5]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_5_13_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data5_rsci_q_d[111:104]), weight_mem_write_arbxbar_xbar_for_1_for_not_395_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_410_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[6]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_6_13_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data6_rsci_q_d[111:104]), weight_mem_write_arbxbar_xbar_for_1_for_not_410_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_425_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[7]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_7_13_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data7_rsci_q_d[111:104]), weight_mem_write_arbxbar_xbar_for_1_for_not_425_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_440_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[8]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_8_13_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data8_rsci_q_d[111:104]), weight_mem_write_arbxbar_xbar_for_1_for_not_440_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_455_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[9]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_9_13_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data9_rsci_q_d[111:104]), weight_mem_write_arbxbar_xbar_for_1_for_not_455_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_470_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[10]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_10_13_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data10_rsci_q_d[111:104]), weight_mem_write_arbxbar_xbar_for_1_for_not_470_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_485_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[11]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_11_13_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data11_rsci_q_d[111:104]), weight_mem_write_arbxbar_xbar_for_1_for_not_485_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_500_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[12]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_12_13_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data12_rsci_q_d[111:104]), weight_mem_write_arbxbar_xbar_for_1_for_not_500_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_515_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[13]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_13_13_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data13_rsci_q_d[111:104]), weight_mem_write_arbxbar_xbar_for_1_for_not_515_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_290_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[14]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_14_13_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data14_rsci_q_d[111:104]), weight_mem_write_arbxbar_xbar_for_1_for_not_290_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_305_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[15]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_15_13_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data15_rsci_q_d[111:104]), weight_mem_write_arbxbar_xbar_for_1_for_not_305_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_319_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[0]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_0_14_lpi_1_dfm_2 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data0_rsci_q_d[119:112]), weight_mem_write_arbxbar_xbar_for_1_for_not_319_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_334_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[1]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_1_14_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data1_rsci_q_d[119:112]), weight_mem_write_arbxbar_xbar_for_1_for_not_334_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_349_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[2]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_2_14_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data2_rsci_q_d[119:112]), weight_mem_write_arbxbar_xbar_for_1_for_not_349_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_364_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[3]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_3_14_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data3_rsci_q_d[119:112]), weight_mem_write_arbxbar_xbar_for_1_for_not_364_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_379_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[4]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_4_14_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data4_rsci_q_d[119:112]), weight_mem_write_arbxbar_xbar_for_1_for_not_379_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_394_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[5]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_5_14_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data5_rsci_q_d[119:112]), weight_mem_write_arbxbar_xbar_for_1_for_not_394_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_409_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[6]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_6_14_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data6_rsci_q_d[119:112]), weight_mem_write_arbxbar_xbar_for_1_for_not_409_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_424_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[7]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_7_14_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data7_rsci_q_d[119:112]), weight_mem_write_arbxbar_xbar_for_1_for_not_424_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_439_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[8]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_8_14_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data8_rsci_q_d[119:112]), weight_mem_write_arbxbar_xbar_for_1_for_not_439_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_454_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[9]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_9_14_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data9_rsci_q_d[119:112]), weight_mem_write_arbxbar_xbar_for_1_for_not_454_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_469_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[10]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_10_14_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data10_rsci_q_d[119:112]), weight_mem_write_arbxbar_xbar_for_1_for_not_469_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_484_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[11]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_11_14_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data11_rsci_q_d[119:112]), weight_mem_write_arbxbar_xbar_for_1_for_not_484_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_499_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[12]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_12_14_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data12_rsci_q_d[119:112]), weight_mem_write_arbxbar_xbar_for_1_for_not_499_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_514_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[13]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_13_14_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data13_rsci_q_d[119:112]), weight_mem_write_arbxbar_xbar_for_1_for_not_514_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_289_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[14]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_14_14_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data14_rsci_q_d[119:112]), weight_mem_write_arbxbar_xbar_for_1_for_not_289_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_304_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[15]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_15_14_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data15_rsci_q_d[119:112]), weight_mem_write_arbxbar_xbar_for_1_for_not_304_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_318_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[0]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_0_15_lpi_1_dfm_2 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data0_rsci_q_d[127:120]), weight_mem_write_arbxbar_xbar_for_1_for_not_318_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_333_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[1]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_1_15_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data1_rsci_q_d[127:120]), weight_mem_write_arbxbar_xbar_for_1_for_not_333_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_348_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[2]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_2_15_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data2_rsci_q_d[127:120]), weight_mem_write_arbxbar_xbar_for_1_for_not_348_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_363_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[3]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_3_15_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data3_rsci_q_d[127:120]), weight_mem_write_arbxbar_xbar_for_1_for_not_363_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_378_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[4]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_4_15_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data4_rsci_q_d[127:120]), weight_mem_write_arbxbar_xbar_for_1_for_not_378_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_393_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[5]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_5_15_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data5_rsci_q_d[127:120]), weight_mem_write_arbxbar_xbar_for_1_for_not_393_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_408_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[6]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_6_15_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data6_rsci_q_d[127:120]), weight_mem_write_arbxbar_xbar_for_1_for_not_408_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_423_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[7]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_7_15_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data7_rsci_q_d[127:120]), weight_mem_write_arbxbar_xbar_for_1_for_not_423_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_438_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[8]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_8_15_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data8_rsci_q_d[127:120]), weight_mem_write_arbxbar_xbar_for_1_for_not_438_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_453_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[9]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_9_15_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data9_rsci_q_d[127:120]), weight_mem_write_arbxbar_xbar_for_1_for_not_453_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_468_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[10]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_10_15_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data10_rsci_q_d[127:120]), weight_mem_write_arbxbar_xbar_for_1_for_not_468_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_483_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[11]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_11_15_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data11_rsci_q_d[127:120]), weight_mem_write_arbxbar_xbar_for_1_for_not_483_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_498_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[12]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_12_15_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data12_rsci_q_d[127:120]), weight_mem_write_arbxbar_xbar_for_1_for_not_498_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_513_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[13]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_13_15_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data13_rsci_q_d[127:120]), weight_mem_write_arbxbar_xbar_for_1_for_not_513_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_288_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[14]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_14_15_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data14_rsci_q_d[127:120]), weight_mem_write_arbxbar_xbar_for_1_for_not_288_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_303_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva[15]);
  assign weight_mem_run_1_bankread_rsp_rdata_data_15_15_lpi_1_dfm_3 = MUX_v_8_2_2(8'b00000000,
      (weight_mem_banks_bank_array_impl_data15_rsci_q_d[127:120]), weight_mem_write_arbxbar_xbar_for_1_for_not_303_nl);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_0_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_0_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_132_itm[1:0]) , (PECore_RunMac_if_mux_131_itm[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_1_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_1_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_132_itm[1:0]) , (PECore_RunMac_if_mux_131_itm[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_2_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_2_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_132_itm[1:0]) , (PECore_RunMac_if_mux_131_itm[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_3_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_3_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_132_itm[1:0]) , (PECore_RunMac_if_mux_131_itm[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_4_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_4_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_132_itm[1:0]) , (PECore_RunMac_if_mux_131_itm[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_5_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_5_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_132_itm[1:0]) , (PECore_RunMac_if_mux_131_itm[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_6_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_6_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_132_itm[1:0]) , (PECore_RunMac_if_mux_131_itm[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_7_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_7_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_132_itm[1:0]) , (PECore_RunMac_if_mux_131_itm[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_8_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_8_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_132_itm[1:0]) , (PECore_RunMac_if_mux_131_itm[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_9_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_9_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_132_itm[1:0]) , (PECore_RunMac_if_mux_131_itm[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_10_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_10_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_132_itm[1:0]) , (PECore_RunMac_if_mux_131_itm[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_11_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_11_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_132_itm[1:0]) , (PECore_RunMac_if_mux_131_itm[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_12_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_12_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_132_itm[1:0]) , (PECore_RunMac_if_mux_131_itm[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_13_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_13_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_132_itm[1:0]) , (PECore_RunMac_if_mux_131_itm[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_14_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_14_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_132_itm[1:0]) , (PECore_RunMac_if_mux_131_itm[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_15_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_15_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_132_itm[1:0]) , (PECore_RunMac_if_mux_131_itm[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_0_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_0_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_133_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_1_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_1_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_133_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_2_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_2_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_133_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_3_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_3_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_133_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_4_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_4_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_133_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_5_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_5_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_133_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_6_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_6_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_133_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_7_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_7_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_133_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_8_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_8_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_133_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_9_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_9_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_133_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_10_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_10_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_133_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_11_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_11_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_133_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_12_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_12_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_133_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_13_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_13_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_133_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_14_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_14_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_133_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_15_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_15_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_133_itm[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_0_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_0_lpi_1_dfm_3,
      {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm , (PECore_RunMac_if_mux_135_itm[2:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_1_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_1_lpi_1_dfm_3,
      {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm , (PECore_RunMac_if_mux_135_itm[2:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_2_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_2_lpi_1_dfm_3,
      {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm , (PECore_RunMac_if_mux_135_itm[2:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_3_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_3_lpi_1_dfm_3,
      {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm , (PECore_RunMac_if_mux_135_itm[2:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_4_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_4_lpi_1_dfm_3,
      {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm , (PECore_RunMac_if_mux_135_itm[2:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_5_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_5_lpi_1_dfm_3,
      {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm , (PECore_RunMac_if_mux_135_itm[2:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_6_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_6_lpi_1_dfm_3,
      {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm , (PECore_RunMac_if_mux_135_itm[2:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_7_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_7_lpi_1_dfm_3,
      {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm , (PECore_RunMac_if_mux_135_itm[2:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_8_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_8_lpi_1_dfm_3,
      {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm , (PECore_RunMac_if_mux_135_itm[2:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_9_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_9_lpi_1_dfm_3,
      {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm , (PECore_RunMac_if_mux_135_itm[2:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_10_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_10_lpi_1_dfm_3,
      {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm , (PECore_RunMac_if_mux_135_itm[2:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_11_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_11_lpi_1_dfm_3,
      {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm , (PECore_RunMac_if_mux_135_itm[2:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_12_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_12_lpi_1_dfm_3,
      {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm , (PECore_RunMac_if_mux_135_itm[2:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_13_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_13_lpi_1_dfm_3,
      {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm , (PECore_RunMac_if_mux_135_itm[2:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_14_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_14_lpi_1_dfm_3,
      {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm , (PECore_RunMac_if_mux_135_itm[2:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_15_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_15_lpi_1_dfm_3,
      {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm , (PECore_RunMac_if_mux_135_itm[2:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_0_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_0_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_13_itm[1:0]) , (reg_PECore_RunMac_if_mux_10_ftd_1[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_1_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_1_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_13_itm[1:0]) , (reg_PECore_RunMac_if_mux_10_ftd_1[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_2_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_2_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_13_itm[1:0]) , (reg_PECore_RunMac_if_mux_10_ftd_1[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_3_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_3_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_13_itm[1:0]) , (reg_PECore_RunMac_if_mux_10_ftd_1[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_4_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_4_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_13_itm[1:0]) , (reg_PECore_RunMac_if_mux_10_ftd_1[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_5_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_5_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_13_itm[1:0]) , (reg_PECore_RunMac_if_mux_10_ftd_1[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_6_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_6_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_13_itm[1:0]) , (reg_PECore_RunMac_if_mux_10_ftd_1[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_7_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_7_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_13_itm[1:0]) , (reg_PECore_RunMac_if_mux_10_ftd_1[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_8_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_8_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_13_itm[1:0]) , (reg_PECore_RunMac_if_mux_10_ftd_1[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_9_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_9_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_13_itm[1:0]) , (reg_PECore_RunMac_if_mux_10_ftd_1[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_10_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_10_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_13_itm[1:0]) , (reg_PECore_RunMac_if_mux_10_ftd_1[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_11_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_11_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_13_itm[1:0]) , (reg_PECore_RunMac_if_mux_10_ftd_1[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_12_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_12_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_13_itm[1:0]) , (reg_PECore_RunMac_if_mux_10_ftd_1[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_13_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_13_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_13_itm[1:0]) , (reg_PECore_RunMac_if_mux_10_ftd_1[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_14_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_14_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_13_itm[1:0]) , (reg_PECore_RunMac_if_mux_10_ftd_1[1:0])});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_15_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_15_lpi_1_dfm_3,
      {(PECore_RunMac_if_mux_13_itm[1:0]) , (reg_PECore_RunMac_if_mux_10_ftd_1[1:0])});
  assign nl_operator_4_false_acc_psp_1_sva_1 = 4'b1011 + conv_u2u_3_4(adpfloat_tmp_to_fixed_20U_14U_acc_sdt_1_sva_mx0w2[3:1]);
  assign operator_4_false_acc_psp_1_sva_1 = nl_operator_4_false_acc_psp_1_sva_1[3:0];
  assign nl_operator_4_false_acc_psp_2_sva_1 = 4'b1011 + conv_u2u_3_4(adpfloat_tmp_to_fixed_20U_14U_acc_sdt_2_sva_mx0w1[3:1]);
  assign operator_4_false_acc_psp_2_sva_1 = nl_operator_4_false_acc_psp_2_sva_1[3:0];
  assign nl_operator_4_false_acc_psp_3_sva_1 = 4'b1011 + conv_u2u_3_4(adpfloat_tmp_to_fixed_20U_14U_acc_sdt_3_sva_mx0w1[3:1]);
  assign operator_4_false_acc_psp_3_sva_1 = nl_operator_4_false_acc_psp_3_sva_1[3:0];
  assign nl_operator_4_false_acc_psp_4_sva_1 = 4'b1011 + conv_u2u_3_4(adpfloat_tmp_to_fixed_20U_14U_acc_sdt_4_sva_mx0w1[3:1]);
  assign operator_4_false_acc_psp_4_sva_1 = nl_operator_4_false_acc_psp_4_sva_1[3:0];
  assign nl_operator_4_false_acc_psp_5_sva_1 = 4'b1011 + conv_u2u_3_4(adpfloat_tmp_to_fixed_20U_14U_acc_sdt_5_sva_mx0w1[3:1]);
  assign operator_4_false_acc_psp_5_sva_1 = nl_operator_4_false_acc_psp_5_sva_1[3:0];
  assign nl_operator_4_false_acc_psp_8_sva_1 = 4'b1011 + conv_u2u_3_4(adpfloat_tmp_to_fixed_20U_14U_acc_sdt_8_sva_mx0w1[3:1]);
  assign operator_4_false_acc_psp_8_sva_1 = nl_operator_4_false_acc_psp_8_sva_1[3:0];
  assign nl_operator_4_false_acc_psp_9_sva_1 = 4'b1011 + conv_u2u_3_4(adpfloat_tmp_to_fixed_20U_14U_acc_sdt_9_sva_mx0w1[3:1]);
  assign operator_4_false_acc_psp_9_sva_1 = nl_operator_4_false_acc_psp_9_sva_1[3:0];
  assign nl_operator_4_false_acc_psp_12_sva_1 = 4'b1011 + conv_u2u_3_4(adpfloat_tmp_to_fixed_20U_14U_acc_sdt_12_sva_mx0w1[3:1]);
  assign operator_4_false_acc_psp_12_sva_1 = nl_operator_4_false_acc_psp_12_sva_1[3:0];
  assign nl_operator_4_false_acc_psp_13_sva_1 = 4'b1011 + conv_u2u_3_4(z_out_50[3:1]);
  assign operator_4_false_acc_psp_13_sva_1 = nl_operator_4_false_acc_psp_13_sva_1[3:0];
  assign nl_operator_4_false_acc_psp_14_sva_1 = 4'b1011 + conv_u2u_3_4(adpfloat_tmp_to_fixed_20U_14U_acc_sdt_14_sva_1[3:1]);
  assign operator_4_false_acc_psp_14_sva_1 = nl_operator_4_false_acc_psp_14_sva_1[3:0];
  assign nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_14_sva_1 = conv_u2u_3_4(input_mem_banks_write_if_for_if_mux_cse[110:108])
      + conv_u2u_3_4(PECore_RunBias_if_for_if_bias_tmp2_mux_17);
  assign adpfloat_tmp_to_fixed_20U_14U_acc_sdt_14_sva_1 = nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_14_sva_1[3:0];
  assign nl_operator_4_false_acc_psp_15_sva_1 = 4'b1011 + conv_u2u_3_4(adpfloat_tmp_to_fixed_20U_14U_acc_sdt_15_sva_1[3:1]);
  assign operator_4_false_acc_psp_15_sva_1 = nl_operator_4_false_acc_psp_15_sva_1[3:0];
  assign nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_15_sva_1 = conv_u2u_3_4(input_mem_banks_write_if_for_if_mux_cse[118:116])
      + conv_u2u_3_4(PECore_RunBias_if_for_if_bias_tmp2_mux_17);
  assign adpfloat_tmp_to_fixed_20U_14U_acc_sdt_15_sva_1 = nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_15_sva_1[3:0];
  assign nl_operator_4_false_acc_psp_sva_1 = 4'b1011 + conv_u2u_3_4(adpfloat_tmp_to_fixed_20U_14U_acc_sdt_sva_1[3:1]);
  assign operator_4_false_acc_psp_sva_1 = nl_operator_4_false_acc_psp_sva_1[3:0];
  assign nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_sva_1 = conv_u2u_3_4(input_mem_banks_write_if_for_if_mux_cse[126:124])
      + conv_u2u_3_4(PECore_RunBias_if_for_if_bias_tmp2_mux_17);
  assign adpfloat_tmp_to_fixed_20U_14U_acc_sdt_sva_1 = nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_sva_1[3:0];
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_12_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_12_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_123_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_13_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_13_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_123_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_14_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_14_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_123_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_2
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_15_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_15_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_123_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_10_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_10_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_123_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_11_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_11_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_123_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_8_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_8_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_123_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_9_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_9_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_123_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_6_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_6_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_123_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_7_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_7_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_123_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_5_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_5_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_123_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_4_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_4_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_123_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_15
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_13_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_13_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_125_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_17
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_12_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_12_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_125_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_19
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_11_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_11_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_125_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_21
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_10_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_10_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_125_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_23
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_9_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_9_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_125_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_25
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_8_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_8_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_125_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_27
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_7_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_7_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_125_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_29
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_6_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_6_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_125_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_31
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_5_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_5_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_125_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_33
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_4_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_4_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_125_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_35
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_3_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_3_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_125_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_37
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_2_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_2_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_125_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_39
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_1_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_1_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_125_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_41
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_0_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_0_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_125_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_14_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_14_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_124_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_13_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_13_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_124_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_12_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_12_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_124_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_11_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_11_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_124_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_10_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_10_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_124_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_9_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_9_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_124_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_8_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_8_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_124_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_7_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_7_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_124_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_6_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_6_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_124_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_5_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_5_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_124_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_4_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_4_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_124_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_3_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_3_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_124_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_2_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_2_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_124_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_1_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_1_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_124_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_0_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_0_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_124_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_14_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_14_lpi_1_dfm_3,
      PECore_RunMac_if_mux_134_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_13_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_13_lpi_1_dfm_3,
      PECore_RunMac_if_mux_134_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_12_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_12_lpi_1_dfm_3,
      PECore_RunMac_if_mux_134_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_11_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_11_lpi_1_dfm_3,
      PECore_RunMac_if_mux_134_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_10_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_10_lpi_1_dfm_3,
      PECore_RunMac_if_mux_134_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_9_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_9_lpi_1_dfm_3,
      PECore_RunMac_if_mux_134_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_8_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_8_lpi_1_dfm_3,
      PECore_RunMac_if_mux_134_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_7_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_7_lpi_1_dfm_3,
      PECore_RunMac_if_mux_134_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_6_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_6_lpi_1_dfm_3,
      PECore_RunMac_if_mux_134_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_5_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_5_lpi_1_dfm_3,
      PECore_RunMac_if_mux_134_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_4_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_4_lpi_1_dfm_3,
      PECore_RunMac_if_mux_134_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_3_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_3_lpi_1_dfm_3,
      PECore_RunMac_if_mux_134_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_2_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_2_lpi_1_dfm_3,
      PECore_RunMac_if_mux_134_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_1_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_1_lpi_1_dfm_3,
      PECore_RunMac_if_mux_134_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_0_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_0_lpi_1_dfm_3,
      PECore_RunMac_if_mux_134_itm[3:0]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_14_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_14_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_129_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_13_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_13_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_129_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_12_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_12_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_129_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_11_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_11_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_129_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_10_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_10_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_129_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_9_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_9_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_129_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_8_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_8_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_129_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_14_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_14_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_128_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_13_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_13_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_128_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_12_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_12_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_128_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_11_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_11_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_128_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_10_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_10_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_128_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_9_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_9_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_128_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_8_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_8_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_128_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_7_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_7_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_128_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_6_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_6_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_128_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_5_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_5_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_128_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_4_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_4_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_128_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_3_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_3_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_128_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_2_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_2_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_128_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_1_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_1_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_128_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_0_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_0_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_128_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_14_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_14_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_127_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_13_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_13_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_127_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_12_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_12_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_127_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_11_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_11_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_127_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_10_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_10_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_127_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_9_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_9_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_127_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_8_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_8_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_127_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_7_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_7_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_127_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_6_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_6_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_127_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_5_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_5_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_127_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_4_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_4_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_127_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_3_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_3_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_127_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_2_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_2_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_127_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_1_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_1_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_127_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_0_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_0_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_127_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_0_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_0_lpi_1_dfm_3,
      {(reg_PECore_RunMac_if_mux_1_ftd_1[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_1_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_1_lpi_1_dfm_3,
      {(reg_PECore_RunMac_if_mux_1_ftd_1[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_2_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_2_lpi_1_dfm_3,
      {(reg_PECore_RunMac_if_mux_1_ftd_1[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_3_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_3_lpi_1_dfm_3,
      {(reg_PECore_RunMac_if_mux_1_ftd_1[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_4_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_4_lpi_1_dfm_3,
      {(reg_PECore_RunMac_if_mux_1_ftd_1[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_5_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_5_lpi_1_dfm_3,
      {(reg_PECore_RunMac_if_mux_1_ftd_1[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_6_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_6_lpi_1_dfm_3,
      {(reg_PECore_RunMac_if_mux_1_ftd_1[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_7_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_7_lpi_1_dfm_3,
      {(reg_PECore_RunMac_if_mux_1_ftd_1[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_8_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_8_lpi_1_dfm_3,
      {(reg_PECore_RunMac_if_mux_1_ftd_1[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_9_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_9_lpi_1_dfm_3,
      {(reg_PECore_RunMac_if_mux_1_ftd_1[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_10_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_10_lpi_1_dfm_3,
      {(reg_PECore_RunMac_if_mux_1_ftd_1[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_11_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_11_lpi_1_dfm_3,
      {(reg_PECore_RunMac_if_mux_1_ftd_1[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_12_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_12_lpi_1_dfm_3,
      {(reg_PECore_RunMac_if_mux_1_ftd_1[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_13_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_13_lpi_1_dfm_3,
      {(reg_PECore_RunMac_if_mux_1_ftd_1[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_14_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_14_lpi_1_dfm_3,
      {(reg_PECore_RunMac_if_mux_1_ftd_1[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_15_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_15_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_15_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_15_lpi_1_dfm_3,
      {(reg_PECore_RunMac_if_mux_1_ftd_1[2:0]) , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm});
  assign nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_6_sva_1 = conv_u2u_3_4(input_mem_banks_write_if_for_if_mux_cse[46:44])
      + conv_u2u_3_4(PECore_RunBias_if_for_if_bias_tmp2_mux_17);
  assign adpfloat_tmp_to_fixed_20U_14U_acc_sdt_6_sva_1 = nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_6_sva_1[3:0];
  assign nl_operator_4_false_acc_psp_6_sva_1 = 4'b1011 + conv_u2u_3_4(adpfloat_tmp_to_fixed_20U_14U_acc_sdt_6_sva_1[3:1]);
  assign operator_4_false_acc_psp_6_sva_1 = nl_operator_4_false_acc_psp_6_sva_1[3:0];
  assign nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_7_sva_1 = conv_u2u_3_4(input_mem_banks_write_if_for_if_mux_cse[54:52])
      + conv_u2u_3_4(PECore_RunBias_if_for_if_bias_tmp2_mux_17);
  assign adpfloat_tmp_to_fixed_20U_14U_acc_sdt_7_sva_1 = nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_7_sva_1[3:0];
  assign nl_operator_4_false_acc_psp_7_sva_1 = 4'b1011 + conv_u2u_3_4(adpfloat_tmp_to_fixed_20U_14U_acc_sdt_7_sva_1[3:1]);
  assign operator_4_false_acc_psp_7_sva_1 = nl_operator_4_false_acc_psp_7_sva_1[3:0];
  assign nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_10_sva_1 = conv_u2u_3_4(input_mem_banks_write_if_for_if_mux_cse[78:76])
      + conv_u2u_3_4(PECore_RunBias_if_for_if_bias_tmp2_mux_17);
  assign adpfloat_tmp_to_fixed_20U_14U_acc_sdt_10_sva_1 = nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_10_sva_1[3:0];
  assign nl_operator_4_false_acc_psp_10_sva_1 = 4'b1011 + conv_u2u_3_4(adpfloat_tmp_to_fixed_20U_14U_acc_sdt_10_sva_1[3:1]);
  assign operator_4_false_acc_psp_10_sva_1 = nl_operator_4_false_acc_psp_10_sva_1[3:0];
  assign nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_11_sva_1 = conv_u2u_3_4(input_mem_banks_write_if_for_if_mux_cse[86:84])
      + conv_u2u_3_4(PECore_RunBias_if_for_if_bias_tmp2_mux_17);
  assign adpfloat_tmp_to_fixed_20U_14U_acc_sdt_11_sva_1 = nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_11_sva_1[3:0];
  assign nl_operator_4_false_acc_psp_11_sva_1 = 4'b1011 + conv_u2u_3_4(adpfloat_tmp_to_fixed_20U_14U_acc_sdt_11_sva_1[3:1]);
  assign operator_4_false_acc_psp_11_sva_1 = nl_operator_4_false_acc_psp_11_sva_1[3:0];
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_14_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_14_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_14_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_14_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_11_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_13_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_13_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_13_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_13_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_11_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_12_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_12_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_12_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_12_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_11_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_11_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_11_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_11_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_11_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_11_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_10_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_10_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_10_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_10_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_11_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_9_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_9_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_9_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_9_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_11_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_8_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_8_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_8_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_8_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_11_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_7_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_7_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_11_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_6_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_6_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_11_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_5_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_5_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_11_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_4_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_4_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_11_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_3_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_3_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_11_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_2_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_2_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_11_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_1_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_1_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_11_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_0_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_0_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_11_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_7_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_7_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_7_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_7_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_129_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_6_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_6_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_6_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_6_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_129_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_5_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_5_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_5_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_5_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_129_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_4_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_4_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_4_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_4_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_129_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_3_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_3_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_3_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_3_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_129_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_2_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_2_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_2_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_2_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_129_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_1_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_1_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_1_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_1_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_129_ftd_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44
      = MUX_v_8_16_2(weight_mem_run_1_bankread_rsp_rdata_data_0_0_lpi_1_dfm_2, weight_mem_run_1_bankread_rsp_rdata_data_1_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_2_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_3_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_4_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_5_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_6_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_7_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_8_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_9_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_10_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_11_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_12_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_13_0_lpi_1_dfm_3,
      weight_mem_run_1_bankread_rsp_rdata_data_14_0_lpi_1_dfm_3, weight_mem_run_1_bankread_rsp_rdata_data_15_0_lpi_1_dfm_3,
      reg_PECore_RunMac_if_mux_129_ftd_1);
  assign PECore_RunBias_if_for_if_bias_tmp2_mux_17 = MUX_v_3_2_2(pe_manager_adplfloat_bias_bias_0_sva,
      pe_manager_adplfloat_bias_bias_1_sva, reg_PECore_RunMac_if_mux_142_ftd_1[0]);
  assign PECore_PushAxiRsp_if_asn_66 = ~(input_mem_banks_load_store_for_else_and_cse_1
      | crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm);
  assign PECore_PushAxiRsp_if_asn_68 = input_mem_banks_load_store_for_else_and_cse_1
      & (~ crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm);
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_5 = (rva_in_PopNB_mio_mrgout_dat_sva[150])
      & PECore_DecodeAxiRead_switch_lp_nor_2_itm;
  assign PECore_DecodeAxiRead_switch_lp_nor_10_cse_1 = ~(PECore_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva
      | PECore_CheckStart_start_reg_sva | PECore_DecodeAxiRead_switch_lp_nor_tmp);
  assign PECore_PushAxiRsp_if_asn_70 = ~(input_mem_banks_load_store_for_else_and_cse
      | crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm);
  assign Arbiter_16U_Roundrobin_pick_mux_2460_tmp_14 = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign Arbiter_16U_Roundrobin_pick_mux_2460_tmp_13 = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_1,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_1_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign Arbiter_16U_Roundrobin_pick_mux_2460_tmp_12 = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_2,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_2_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign Arbiter_16U_Roundrobin_pick_mux_2460_tmp_11 = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_3,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_3_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign Arbiter_16U_Roundrobin_pick_mux_2460_tmp_10 = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_4,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_4_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign Arbiter_16U_Roundrobin_pick_mux_2460_tmp_9 = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_5,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_5_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign Arbiter_16U_Roundrobin_pick_mux_2460_tmp_8 = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_6,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_6_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign Arbiter_16U_Roundrobin_pick_mux_2460_tmp_7 = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_7,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_7_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign Arbiter_16U_Roundrobin_pick_mux_2460_tmp_6 = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_8,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_8_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign Arbiter_16U_Roundrobin_pick_mux_2460_tmp_5 = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_9,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_9_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign Arbiter_16U_Roundrobin_pick_mux_2460_tmp_4 = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_10,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_10_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign Arbiter_16U_Roundrobin_pick_mux_2460_tmp_3 = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_11,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_11_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign Arbiter_16U_Roundrobin_pick_mux_2460_tmp_2 = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_12,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_12_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign Arbiter_16U_Roundrobin_pick_mux_2460_tmp_1 = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_13,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_13_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign Arbiter_16U_Roundrobin_pick_mux_2460_tmp_0 = MUX_s_1_2_2(reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_14,
      weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_14_itm,
      weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse);
  assign or_tmp_18 = (rva_in_PopNB_mioi_idat_mxwt[168]) | is_start_sva | (rva_in_PopNB_mioi_idat_mxwt[151:148]!=4'b0110)
      | (~ rva_in_PopNB_mioi_ivld_mxwt);
  assign or_tmp_20 = (~ (rva_in_PopNB_mioi_idat_mxwt[168])) | is_start_sva | (rva_in_PopNB_mioi_idat_mxwt[151:148]!=4'b0110)
      | (~ rva_in_PopNB_mioi_ivld_mxwt);
  assign or_dcpl = state_2_0_sva_0 | state_2_0_sva_1;
  assign or_dcpl_34 = ~((weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]) & weight_mem_read_arbxbar_xbar_for_3_16_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp);
  assign and_dcpl_135 = (~ state_2_0_sva_2) & state_2_0_sva_1;
  assign and_dcpl_210 = is_start_sva & (~ state_2_0_sva_0);
  assign and_dcpl_211 = and_dcpl_135 & and_dcpl_210;
  assign or_tmp_545 = (~ PECore_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva)
      | (rva_in_PopNB_mio_mrgout_dat_sva[168]);
  assign or_55_cse = state_2_0_sva_2 | state_2_0_sva_1 | (~ input_port_PopNB_mioi_ivld_mxwt)
      | state_2_0_sva_0;
  assign nand_199_cse = ~((rva_in_PopNB_mioi_idat_mxwt[150]) & rva_in_PopNB_mioi_ivld_mxwt);
  assign or_dcpl_247 = state_2_0_sva_0 | (~ is_start_sva);
  assign and_dcpl_414 = and_5335_cse & (~ reg_PECore_RunMac_asn_15_itm_1_ftd);
  assign or_dcpl_251 = (fsm_output[4:3]!=2'b00);
  assign or_tmp_1286 = is_start_sva | (rva_in_PopNB_mioi_idat_mxwt[151:148]!=4'b0110)
      | (~ rva_in_PopNB_mioi_ivld_mxwt);
  assign or_dcpl_285 = (rva_in_PopNB_mioi_idat_mxwt[148]) | (~ (rva_in_PopNB_mioi_idat_mxwt[168]));
  assign or_dcpl_286 = or_dcpl_285 | is_start_sva;
  assign and_dcpl_437 = and_dcpl_414 & reg_PECore_RunMac_asn_15_itm_1_ftd_2 & PECore_DecodeAxiRead_case_4_switch_lp_and_2_itm;
  assign and_dcpl_439 = and_dcpl_414 & reg_PECore_RunMac_asn_15_itm_1_ftd_2 & (~
      PECore_DecodeAxiRead_case_4_switch_lp_and_2_itm);
  assign or_dcpl_295 = (~ and_5335_cse) | reg_PECore_RunMac_asn_15_itm_1_ftd | (~
      reg_PECore_RunMac_asn_15_itm_1_ftd_2);
  assign and_dcpl_440 = reg_PECore_RunMac_asn_15_itm_1_ftd_2 & while_stage_0_2;
  assign or_dcpl_300 = (rva_in_PopNB_mioi_idat_mxwt[149:148]!=2'b00);
  assign or_dcpl_301 = or_dcpl_300 | (~ (rva_in_PopNB_mioi_idat_mxwt[168])) | is_start_sva;
  assign or_dcpl_302 = (rva_in_PopNB_mioi_idat_mxwt[151:150]!=2'b01);
  assign or_dcpl_306 = (~ PECore_DecodeAxiWrite_case_4_switch_lp_nor_15_tmp) | (~
      (rva_in_PopNB_mioi_idat_mxwt[133])) | (~ rva_in_PopNB_mioi_ivld_mxwt) | or_dcpl_302
      | or_dcpl_301;
  assign or_dcpl_310 = (~ (rva_in_PopNB_mioi_idat_mxwt[134])) | (~ PECore_DecodeAxiWrite_case_4_switch_lp_nor_11_tmp)
      | (~ rva_in_PopNB_mioi_ivld_mxwt) | or_dcpl_302 | or_dcpl_301;
  assign or_dcpl_313 = or_dcpl_300 | (~ (rva_in_PopNB_mioi_idat_mxwt[168])) | (~
      (rva_in_PopNB_mioi_idat_mxwt[132])) | is_start_sva;
  assign or_dcpl_327 = (rva_in_PopNB_mioi_idat_mxwt[151]) | (rva_in_PopNB_mioi_idat_mxwt[149]);
  assign or_dcpl_334 = nand_199_cse | or_dcpl_327 | or_dcpl_285 | (~ PECore_DecodeAxiWrite_case_4_switch_lp_nor_7_tmp)
      | (~ (rva_in_PopNB_mioi_idat_mxwt[132])) | is_start_sva;
  assign or_dcpl_362 = ~(state_2_0_sva_0 & is_start_sva);
  assign or_dcpl_363 = or_500_cse | (~ is_start_sva);
  assign or_dcpl_364 = or_dcpl_363 | or_dcpl_362;
  assign or_dcpl_365 = or_500_cse | or_dcpl_362;
  assign or_dcpl_369 = ~((~ or_dcpl_363) & pe_config_is_bias_sva & state_2_0_sva_0);
  assign and_dcpl_700 = and_dcpl_135 & pe_config_is_bias_sva & state_2_0_sva_0;
  assign and_dcpl_702 = and_dcpl_135 & (~ pe_config_is_bias_sva) & state_2_0_sva_0;
  assign or_dcpl_370 = or_500_cse | (~ state_2_0_sva_0);
  assign and_dcpl_704 = pe_config_is_cluster_sva & is_start_sva;
  assign and_dcpl_705 = (~ pe_config_is_cluster_sva) & is_start_sva;
  assign and_dcpl_706 = pe_config_is_cluster_sva & (~ state_2_0_sva_0);
  assign and_dcpl_707 = and_dcpl_706 & is_start_sva;
  assign and_dcpl_708 = ~(pe_config_is_cluster_sva | state_2_0_sva_0);
  assign and_dcpl_709 = and_dcpl_708 & is_start_sva;
  assign or_dcpl_374 = nand_199_cse | or_dcpl_327;
  assign or_dcpl_375 = or_dcpl_374 | or_dcpl_286;
  assign or_dcpl_378 = or_dcpl_374 | (~ (rva_in_PopNB_mioi_idat_mxwt[148])) | (rva_in_PopNB_mioi_idat_mxwt[168])
      | is_start_sva;
  assign and_dcpl_725 = (~((weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[0]) &
      weight_mem_read_arbxbar_arbiters_next_0_10_sva)) & (~((weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[0])
      & weight_mem_read_arbxbar_arbiters_next_0_9_sva)) & (~((weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[0])
      & weight_mem_read_arbxbar_arbiters_next_0_11_sva)) & (~((weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[0])
      & weight_mem_read_arbxbar_arbiters_next_0_12_sva)) & (~((weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[0])
      & weight_mem_read_arbxbar_arbiters_next_0_13_sva)) & (~((weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[0])
      & weight_mem_read_arbxbar_arbiters_next_0_14_sva)) & (~((weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[0])
      & weight_mem_read_arbxbar_arbiters_next_0_15_sva)) & weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  assign and_dcpl_726 = ~((~((weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[0]))) | weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_733 = ~((weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[0])
      | weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_748 = (~((weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[1]) &
      weight_mem_read_arbxbar_arbiters_next_1_9_sva)) & (~((weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[1])
      & weight_mem_read_arbxbar_arbiters_next_1_11_sva)) & (~((weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[1])
      & weight_mem_read_arbxbar_arbiters_next_1_12_sva)) & (~((weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[1])
      & weight_mem_read_arbxbar_arbiters_next_1_10_sva)) & (~((weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[1])
      & weight_mem_read_arbxbar_arbiters_next_1_13_sva)) & (~((weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[1])
      & weight_mem_read_arbxbar_arbiters_next_1_15_sva)) & (~((weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[1])
      & weight_mem_read_arbxbar_arbiters_next_1_14_sva)) & weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  assign and_dcpl_749 = ~((~((weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[1]))) | weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_756 = ~((weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[1])
      | weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_771 = (~((weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[2]) &
      weight_mem_read_arbxbar_arbiters_next_2_11_sva)) & (~((weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[2])
      & weight_mem_read_arbxbar_arbiters_next_2_9_sva)) & (~((weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[2])
      & weight_mem_read_arbxbar_arbiters_next_2_10_sva)) & (~((weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[2])
      & weight_mem_read_arbxbar_arbiters_next_2_13_sva)) & (~((weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[2])
      & weight_mem_read_arbxbar_arbiters_next_2_14_sva)) & (~((weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[2])
      & weight_mem_read_arbxbar_arbiters_next_2_12_sva)) & (~((weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[2])
      & weight_mem_read_arbxbar_arbiters_next_2_15_sva)) & weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  assign and_dcpl_772 = ~((~((weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]) |
      (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[2]))) | weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_779 = ~((weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[2])
      | weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_794 = (~((weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[3]) &
      weight_mem_read_arbxbar_arbiters_next_3_9_sva)) & (~((weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[3])
      & weight_mem_read_arbxbar_arbiters_next_3_10_sva)) & (~((weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[3])
      & weight_mem_read_arbxbar_arbiters_next_3_12_sva)) & (~((weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[3])
      & weight_mem_read_arbxbar_arbiters_next_3_13_sva)) & (~((weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[3])
      & weight_mem_read_arbxbar_arbiters_next_3_11_sva)) & (~((weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[3])
      & weight_mem_read_arbxbar_arbiters_next_3_14_sva)) & (~((weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[3])
      & weight_mem_read_arbxbar_arbiters_next_3_15_sva)) & weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  assign and_dcpl_795 = ~((~((weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[3]))) | weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_802 = ~((weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[3])
      | weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_817 = (~((weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[4]) &
      weight_mem_read_arbxbar_arbiters_next_4_11_sva)) & (~((weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[4])
      & weight_mem_read_arbxbar_arbiters_next_4_9_sva)) & (~((weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[4])
      & weight_mem_read_arbxbar_arbiters_next_4_10_sva)) & (~((weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[4])
      & weight_mem_read_arbxbar_arbiters_next_4_12_sva)) & (~((weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[4])
      & weight_mem_read_arbxbar_arbiters_next_4_13_sva)) & (~((weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[4])
      & weight_mem_read_arbxbar_arbiters_next_4_15_sva)) & (~((weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[4])
      & weight_mem_read_arbxbar_arbiters_next_4_14_sva)) & weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  assign and_dcpl_818 = ~((~((weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[4]))) | weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_825 = ~((weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[4])
      | weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_840 = (~((weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[5]) &
      weight_mem_read_arbxbar_arbiters_next_5_14_sva)) & (~((weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[5])
      & weight_mem_read_arbxbar_arbiters_next_5_9_sva)) & (~((weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[5])
      & weight_mem_read_arbxbar_arbiters_next_5_11_sva)) & (~((weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[5])
      & weight_mem_read_arbxbar_arbiters_next_5_12_sva)) & (~((weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[5])
      & weight_mem_read_arbxbar_arbiters_next_5_13_sva)) & (~((weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[5])
      & weight_mem_read_arbxbar_arbiters_next_5_10_sva)) & (~((weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[5])
      & weight_mem_read_arbxbar_arbiters_next_5_15_sva)) & weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  assign and_dcpl_841 = ~((~((weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[5]))) | weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_848 = ~((weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[5])
      | weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_863 = (~(weight_mem_read_arbxbar_arbiters_next_6_10_sva & (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[6])))
      & (~((weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_9_sva))
      & (~((weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_11_sva))
      & (~((weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_12_sva))
      & (~((weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_13_sva))
      & (~((weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_15_sva))
      & (~((weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_14_sva))
      & weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  assign and_dcpl_864 = ~((~((weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]) |
      (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[6]))) | weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_871 = ~((weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[6])
      | weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_886 = (~(weight_mem_read_arbxbar_arbiters_next_7_9_sva & (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[7])))
      & (~((weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_10_sva))
      & (~((weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_13_sva))
      & (~((weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_11_sva))
      & (~((weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_12_sva))
      & (~((weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_15_sva))
      & (~((weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_14_sva))
      & weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  assign and_dcpl_887 = ~((~((weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]) |
      (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[7]))) | weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_894 = ~((weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[7])
      | weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_909 = (~((weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[8]) &
      weight_mem_read_arbxbar_arbiters_next_8_13_sva)) & (~((weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[8])
      & weight_mem_read_arbxbar_arbiters_next_8_9_sva)) & (~((weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[8])
      & weight_mem_read_arbxbar_arbiters_next_8_12_sva)) & (~((weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[8])
      & weight_mem_read_arbxbar_arbiters_next_8_11_sva)) & (~((weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[8])
      & weight_mem_read_arbxbar_arbiters_next_8_10_sva)) & (~((weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[8])
      & weight_mem_read_arbxbar_arbiters_next_8_14_sva)) & (~((weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[8])
      & weight_mem_read_arbxbar_arbiters_next_8_15_sva)) & weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  assign and_dcpl_910 = ~((~((weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[8])
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[8])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[8])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[8])
      | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[8]))) | weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_917 = ~((weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[8])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[8])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[8])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[8]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[8])
      | weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_932 = (~((weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[9]) &
      weight_mem_read_arbxbar_arbiters_next_9_15_sva)) & (~((weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[9])
      & weight_mem_read_arbxbar_arbiters_next_9_9_sva)) & (~((weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[9])
      & weight_mem_read_arbxbar_arbiters_next_9_10_sva)) & (~((weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[9])
      & weight_mem_read_arbxbar_arbiters_next_9_13_sva)) & (~((weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[9])
      & weight_mem_read_arbxbar_arbiters_next_9_12_sva)) & (~((weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[9])
      & weight_mem_read_arbxbar_arbiters_next_9_11_sva)) & (~((weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[9])
      & weight_mem_read_arbxbar_arbiters_next_9_14_sva)) & weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  assign and_dcpl_933 = ~((~((weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[9])
      | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[9])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[9])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[9])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[9]))) | weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_939 = ~((weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[9])
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[9])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[9])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[9]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[9])
      | weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_954 = (~((weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[10]) &
      weight_mem_read_arbxbar_arbiters_next_10_10_sva)) & (~((weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[10])
      & weight_mem_read_arbxbar_arbiters_next_10_15_sva)) & (~((weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[10])
      & weight_mem_read_arbxbar_arbiters_next_10_13_sva)) & (~((weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[10])
      & weight_mem_read_arbxbar_arbiters_next_10_9_sva)) & (~((weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[10])
      & weight_mem_read_arbxbar_arbiters_next_10_14_sva)) & (~((weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[10])
      & weight_mem_read_arbxbar_arbiters_next_10_11_sva)) & (~((weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[10])
      & weight_mem_read_arbxbar_arbiters_next_10_12_sva)) & weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  assign and_dcpl_955 = ~((~((weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[10])
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[10])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[10])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[10])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[10]))) | weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_962 = ~((weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[10]) |
      (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[10])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[10])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[10]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[10])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[10]) | weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_977 = (~((weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[11]) &
      weight_mem_read_arbxbar_arbiters_next_11_10_sva)) & (~((weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[11])
      & weight_mem_read_arbxbar_arbiters_next_11_15_sva)) & (~((weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[11])
      & weight_mem_read_arbxbar_arbiters_next_11_14_sva)) & (~((weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[11])
      & weight_mem_read_arbxbar_arbiters_next_11_9_sva)) & (~((weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[11])
      & weight_mem_read_arbxbar_arbiters_next_11_12_sva)) & (~((weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[11])
      & weight_mem_read_arbxbar_arbiters_next_11_11_sva)) & (~((weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[11])
      & weight_mem_read_arbxbar_arbiters_next_11_13_sva)) & weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  assign and_dcpl_978 = ~((~((weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[11])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[11])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[11])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[11])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[11]))) | weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_985 = ~((weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[11])
      | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[11])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[11])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[11]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[11])
      | weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_1000 = (~(weight_mem_read_arbxbar_arbiters_next_12_10_sva & (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[12])))
      & (~(weight_mem_read_arbxbar_arbiters_next_12_9_sva & (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[12])))
      & (~((weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[12]) & weight_mem_read_arbxbar_arbiters_next_12_12_sva))
      & (~((weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[12]) & weight_mem_read_arbxbar_arbiters_next_12_13_sva))
      & (~((weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[12]) & weight_mem_read_arbxbar_arbiters_next_12_14_sva))
      & (~((weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[12]) & weight_mem_read_arbxbar_arbiters_next_12_15_sva))
      & (~((weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[12]) & weight_mem_read_arbxbar_arbiters_next_12_11_sva))
      & weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  assign and_dcpl_1001 = ~((~((weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[12])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[12])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[12])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[12])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[12]))) | weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_1008 = ~((weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[12]) |
      (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[12])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[12])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[12]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[12])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[12]) | weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_1023 = (~((weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[13])
      & weight_mem_read_arbxbar_arbiters_next_13_10_sva)) & (~(weight_mem_read_arbxbar_arbiters_next_13_9_sva
      & (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[13]))) & (~(weight_mem_read_arbxbar_arbiters_next_13_11_sva
      & (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[13]))) & (~((weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[13])
      & weight_mem_read_arbxbar_arbiters_next_13_12_sva)) & (~((weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[13])
      & weight_mem_read_arbxbar_arbiters_next_13_13_sva)) & (~((weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[13])
      & weight_mem_read_arbxbar_arbiters_next_13_15_sva)) & (~((weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[13])
      & weight_mem_read_arbxbar_arbiters_next_13_14_sva)) & weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  assign and_dcpl_1024 = ~((~((weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[13])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[13])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[13])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[13])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[13]))) | weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_1029 = ~((weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[13]) |
      (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[13])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[13])
      | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[13]) | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[13])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[13]) | weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_1043 = (~((weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[14])
      & weight_mem_read_arbxbar_arbiters_next_14_15_sva)) & (~((weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[14])
      & weight_mem_read_arbxbar_arbiters_next_14_14_sva)) & (~((weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[14])
      & weight_mem_read_arbxbar_arbiters_next_14_13_sva)) & (~((weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[14])
      & weight_mem_read_arbxbar_arbiters_next_14_10_sva)) & (~((weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[14])
      & weight_mem_read_arbxbar_arbiters_next_14_12_sva)) & (~((weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[14])
      & weight_mem_read_arbxbar_arbiters_next_14_11_sva)) & (~ weight_mem_read_arbxbar_xbar_for_3_15_Arbiter_16U_Roundrobin_pick_priority_and_4_tmp)
      & weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  assign and_dcpl_1044 = ~((~((weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[14])
      | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[14])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[14])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[14])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[14]))) | weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_1051 = ~((weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[14]) |
      (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[14])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[14])
      | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[14]) | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[14])
      | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[14]) | weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_1066 = (~((weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[15])
      & weight_mem_read_arbxbar_arbiters_next_15_15_sva)) & (~((weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[15])
      & weight_mem_read_arbxbar_arbiters_next_15_10_sva)) & (~((weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[15])
      & weight_mem_read_arbxbar_arbiters_next_15_9_sva)) & (~((weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[15])
      & weight_mem_read_arbxbar_arbiters_next_15_11_sva)) & (~((weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[15])
      & weight_mem_read_arbxbar_arbiters_next_15_14_sva)) & (~((weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[15])
      & weight_mem_read_arbxbar_arbiters_next_15_13_sva)) & (~((weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[15])
      & weight_mem_read_arbxbar_arbiters_next_15_12_sva)) & weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  assign and_dcpl_1067 = ~((~((weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[15])
      | (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[15])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[15])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[15])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[15]))) | weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_dcpl_1074 = ~((weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[15]) |
      (weight_mem_read_arbxbar_xbar_for_16_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_11_lshift_tmp[15])
      | (weight_mem_read_arbxbar_xbar_for_10_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_12_lshift_tmp[15])
      | (weight_mem_read_arbxbar_xbar_for_15_lshift_tmp[15]) | (weight_mem_read_arbxbar_xbar_for_14_lshift_tmp[15])
      | (weight_mem_read_arbxbar_xbar_for_13_lshift_tmp[15]) | weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp);
  assign and_2164_cse = ~((fsm_output[0]) | (fsm_output[4]));
  assign or_tmp_1334 = (fsm_output[1:0]!=2'b00);
  assign or_tmp_1655 = w_axi_rsp_lpi_1_dfm_1 & (~ crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm)
      & (~ is_start_sva) & (fsm_output[3]);
  assign and_2907_cse = and_dcpl_414 & (~ reg_PECore_RunMac_asn_15_itm_1_ftd_2) &
      while_stage_0_2 & (fsm_output[1]);
  assign or_tmp_2232 = (~ (fsm_output[1])) | is_start_sva;
  assign and_4616_cse = (fsm_output[3:2]!=2'b00);
  assign or_tmp_2557 = or_dcpl_251 | (((~((~(and_dcpl_135 & is_start_sva & state_2_0_sva_0))
      & while_asn_41_itm_1)) | (~ reg_PECore_RunMac_asn_15_itm_1_ftd_1) | reg_PECore_RunMac_asn_15_itm_1_ftd
      | (~(reg_PECore_RunMac_asn_15_itm_1_ftd_2 & while_stage_0_2))) & (fsm_output[1]));
  assign or_3399_cse = (fsm_output[3]) | (fsm_output[1]);
  assign PECore_RunBias_if_accum_vector_out_data_and_15_rgt = and_dcpl_414 & and_dcpl_440
      & (~ PECore_DecodeAxiRead_case_4_switch_lp_and_2_itm) & (~ nor_499_cse);
  assign PECore_RunBias_if_accum_vector_out_data_and_17_cse = PECoreRun_wen & ((and_dcpl_414
      & and_dcpl_440 & PECore_DecodeAxiRead_case_4_switch_lp_and_2_itm & (~ nor_499_cse))
      | PECore_RunBias_if_accum_vector_out_data_and_15_rgt);
  assign weight_mem_banks_bank_array_impl_data0_rsci_d_d = {while_while_and_18_itm
      , weight_write_data_data_mux1h_14_rmff , weight_write_data_data_mux1h_13_rmff
      , weight_write_data_data_mux1h_12_rmff , weight_write_data_data_mux1h_11_rmff
      , weight_write_data_data_mux1h_10_rmff , weight_write_data_data_mux1h_9_rmff
      , weight_write_data_data_mux1h_8_rmff , weight_write_data_data_mux1h_7_rmff
      , weight_write_data_data_mux1h_6_rmff , weight_write_data_data_mux1h_5_rmff
      , weight_write_data_data_mux1h_4_rmff , weight_write_data_data_mux1h_3_rmff
      , weight_write_data_data_mux1h_2_rmff , weight_write_data_data_mux1h_1_rmff
      , weight_write_data_data_mux1h_rmff};
  assign weight_mem_banks_bank_array_impl_data0_rsci_radr_d = MUX_v_12_16_2(weight_read_addrs_0_15_4_lpi_1_dfm_5_mx0,
      (weight_read_addrs_1_lpi_1_dfm_2[15:4]), (weight_read_addrs_2_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_3_lpi_1_dfm_2[15:4]), (weight_read_addrs_4_15_2_lpi_1_dfm_2[13:2]),
      (weight_read_addrs_5_lpi_1_dfm_2[15:4]), (weight_read_addrs_6_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_7_lpi_1_dfm_2[15:4]), (weight_read_addrs_8_15_3_lpi_1_dfm_3[12:1]),
      (weight_read_addrs_9_lpi_1_dfm_3[15:4]), (weight_read_addrs_10_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_11_lpi_1_dfm_3[15:4]), (weight_read_addrs_12_15_2_lpi_1_dfm_3[13:2]),
      (weight_read_addrs_13_lpi_1_dfm_3[15:4]), (weight_read_addrs_14_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_15_lpi_1_dfm_3[15:4]), {weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_3_2_sva_1 , weight_mem_read_arbxbar_xbar_for_3_source_local_3_1_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_3_0_sva_1});
  assign weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_pff = weight_write_addrs_lpi_1_dfm_6[15:4];
  assign weight_mem_banks_bank_array_impl_data0_rsci_we_d_pff = and_3039_cse;
  assign weight_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = or_1405_cse;
  assign weight_mem_banks_bank_array_impl_data1_rsci_d_d = {while_while_and_18_itm
      , weight_write_data_data_mux1h_14_rmff , weight_write_data_data_mux1h_13_rmff
      , weight_write_data_data_mux1h_12_rmff , weight_write_data_data_mux1h_11_rmff
      , weight_write_data_data_mux1h_10_rmff , weight_write_data_data_mux1h_9_rmff
      , weight_write_data_data_mux1h_8_rmff , weight_write_data_data_mux1h_7_rmff
      , weight_write_data_data_mux1h_6_rmff , weight_write_data_data_mux1h_5_rmff
      , weight_write_data_data_mux1h_4_rmff , weight_write_data_data_mux1h_3_rmff
      , weight_write_data_data_mux1h_2_rmff , weight_write_data_data_mux1h_1_rmff
      , weight_write_data_data_mux1h_rmff};
  assign weight_mem_banks_bank_array_impl_data1_rsci_radr_d = MUX_v_12_16_2(weight_read_addrs_0_15_4_lpi_1_dfm_5_mx0,
      (weight_read_addrs_1_lpi_1_dfm_2[15:4]), (weight_read_addrs_2_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_3_lpi_1_dfm_2[15:4]), (weight_read_addrs_4_15_2_lpi_1_dfm_2[13:2]),
      (weight_read_addrs_5_lpi_1_dfm_2[15:4]), (weight_read_addrs_6_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_7_lpi_1_dfm_2[15:4]), (weight_read_addrs_8_15_3_lpi_1_dfm_3[12:1]),
      (weight_read_addrs_9_lpi_1_dfm_3[15:4]), (weight_read_addrs_10_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_11_lpi_1_dfm_3[15:4]), (weight_read_addrs_12_15_2_lpi_1_dfm_3[13:2]),
      (weight_read_addrs_13_lpi_1_dfm_3[15:4]), (weight_read_addrs_14_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_15_lpi_1_dfm_3[15:4]), {weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_4_2_sva_1 , weight_mem_read_arbxbar_xbar_for_3_source_local_4_1_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_4_0_sva_1});
  assign weight_mem_banks_bank_array_impl_data1_rsci_we_d_pff = and_3035_cse;
  assign weight_mem_banks_bank_array_impl_data1_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = or_1409_cse;
  assign weight_mem_banks_bank_array_impl_data2_rsci_d_d = {while_while_and_18_itm
      , weight_write_data_data_mux1h_14_rmff , weight_write_data_data_mux1h_13_rmff
      , weight_write_data_data_mux1h_12_rmff , weight_write_data_data_mux1h_11_rmff
      , weight_write_data_data_mux1h_10_rmff , weight_write_data_data_mux1h_9_rmff
      , weight_write_data_data_mux1h_8_rmff , weight_write_data_data_mux1h_7_rmff
      , weight_write_data_data_mux1h_6_rmff , weight_write_data_data_mux1h_5_rmff
      , weight_write_data_data_mux1h_4_rmff , weight_write_data_data_mux1h_3_rmff
      , weight_write_data_data_mux1h_2_rmff , weight_write_data_data_mux1h_1_rmff
      , weight_write_data_data_mux1h_rmff};
  assign weight_mem_banks_bank_array_impl_data2_rsci_radr_d = MUX_v_12_16_2(weight_read_addrs_0_15_4_lpi_1_dfm_5_mx0,
      (weight_read_addrs_1_lpi_1_dfm_2[15:4]), (weight_read_addrs_2_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_3_lpi_1_dfm_2[15:4]), (weight_read_addrs_4_15_2_lpi_1_dfm_2[13:2]),
      (weight_read_addrs_5_lpi_1_dfm_2[15:4]), (weight_read_addrs_6_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_7_lpi_1_dfm_2[15:4]), (weight_read_addrs_8_15_3_lpi_1_dfm_3[12:1]),
      (weight_read_addrs_9_lpi_1_dfm_3[15:4]), (weight_read_addrs_10_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_11_lpi_1_dfm_3[15:4]), (weight_read_addrs_12_15_2_lpi_1_dfm_3[13:2]),
      (weight_read_addrs_13_lpi_1_dfm_3[15:4]), (weight_read_addrs_14_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_15_lpi_1_dfm_3[15:4]), {weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_5_2_sva_1 , weight_mem_read_arbxbar_xbar_for_3_source_local_5_1_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_5_0_sva_1});
  assign weight_mem_banks_bank_array_impl_data2_rsci_we_d_pff = and_3031_cse;
  assign weight_mem_banks_bank_array_impl_data2_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = or_1413_cse;
  assign weight_mem_banks_bank_array_impl_data3_rsci_d_d = {while_while_and_18_itm
      , weight_write_data_data_mux1h_14_rmff , weight_write_data_data_mux1h_13_rmff
      , weight_write_data_data_mux1h_12_rmff , weight_write_data_data_mux1h_11_rmff
      , weight_write_data_data_mux1h_10_rmff , weight_write_data_data_mux1h_9_rmff
      , weight_write_data_data_mux1h_8_rmff , weight_write_data_data_mux1h_7_rmff
      , weight_write_data_data_mux1h_6_rmff , weight_write_data_data_mux1h_5_rmff
      , weight_write_data_data_mux1h_4_rmff , weight_write_data_data_mux1h_3_rmff
      , weight_write_data_data_mux1h_2_rmff , weight_write_data_data_mux1h_1_rmff
      , weight_write_data_data_mux1h_rmff};
  assign weight_mem_banks_bank_array_impl_data3_rsci_radr_d = MUX_v_12_16_2(weight_read_addrs_0_15_4_lpi_1_dfm_5_mx0,
      (weight_read_addrs_1_lpi_1_dfm_2[15:4]), (weight_read_addrs_2_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_3_lpi_1_dfm_2[15:4]), (weight_read_addrs_4_15_2_lpi_1_dfm_2[13:2]),
      (weight_read_addrs_5_lpi_1_dfm_2[15:4]), (weight_read_addrs_6_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_7_lpi_1_dfm_2[15:4]), (weight_read_addrs_8_15_3_lpi_1_dfm_3[12:1]),
      (weight_read_addrs_9_lpi_1_dfm_3[15:4]), (weight_read_addrs_10_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_11_lpi_1_dfm_3[15:4]), (weight_read_addrs_12_15_2_lpi_1_dfm_3[13:2]),
      (weight_read_addrs_13_lpi_1_dfm_3[15:4]), (weight_read_addrs_14_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_15_lpi_1_dfm_3[15:4]), {weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_6_2_sva_1 , weight_mem_read_arbxbar_xbar_for_3_source_local_6_1_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_6_0_sva_1});
  assign weight_mem_banks_bank_array_impl_data3_rsci_we_d_pff = and_3027_cse;
  assign weight_mem_banks_bank_array_impl_data3_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = or_1417_cse;
  assign weight_mem_banks_bank_array_impl_data4_rsci_d_d = {while_while_and_18_itm
      , weight_write_data_data_mux1h_14_rmff , weight_write_data_data_mux1h_13_rmff
      , weight_write_data_data_mux1h_12_rmff , weight_write_data_data_mux1h_11_rmff
      , weight_write_data_data_mux1h_10_rmff , weight_write_data_data_mux1h_9_rmff
      , weight_write_data_data_mux1h_8_rmff , weight_write_data_data_mux1h_7_rmff
      , weight_write_data_data_mux1h_6_rmff , weight_write_data_data_mux1h_5_rmff
      , weight_write_data_data_mux1h_4_rmff , weight_write_data_data_mux1h_3_rmff
      , weight_write_data_data_mux1h_2_rmff , weight_write_data_data_mux1h_1_rmff
      , weight_write_data_data_mux1h_rmff};
  assign weight_mem_banks_bank_array_impl_data4_rsci_radr_d = MUX_v_12_16_2(weight_read_addrs_0_15_4_lpi_1_dfm_5_mx0,
      (weight_read_addrs_1_lpi_1_dfm_2[15:4]), (weight_read_addrs_2_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_3_lpi_1_dfm_2[15:4]), (weight_read_addrs_4_15_2_lpi_1_dfm_2[13:2]),
      (weight_read_addrs_5_lpi_1_dfm_2[15:4]), (weight_read_addrs_6_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_7_lpi_1_dfm_2[15:4]), (weight_read_addrs_8_15_3_lpi_1_dfm_3[12:1]),
      (weight_read_addrs_9_lpi_1_dfm_3[15:4]), (weight_read_addrs_10_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_11_lpi_1_dfm_3[15:4]), (weight_read_addrs_12_15_2_lpi_1_dfm_3[13:2]),
      (weight_read_addrs_13_lpi_1_dfm_3[15:4]), (weight_read_addrs_14_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_15_lpi_1_dfm_3[15:4]), {weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_7_2_sva_1 , weight_mem_read_arbxbar_xbar_for_3_source_local_7_1_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_7_0_sva_1});
  assign weight_mem_banks_bank_array_impl_data4_rsci_we_d_pff = and_3023_cse;
  assign weight_mem_banks_bank_array_impl_data4_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = or_1421_cse;
  assign weight_mem_banks_bank_array_impl_data5_rsci_d_d = {while_while_and_18_itm
      , weight_write_data_data_mux1h_14_rmff , weight_write_data_data_mux1h_13_rmff
      , weight_write_data_data_mux1h_12_rmff , weight_write_data_data_mux1h_11_rmff
      , weight_write_data_data_mux1h_10_rmff , weight_write_data_data_mux1h_9_rmff
      , weight_write_data_data_mux1h_8_rmff , weight_write_data_data_mux1h_7_rmff
      , weight_write_data_data_mux1h_6_rmff , weight_write_data_data_mux1h_5_rmff
      , weight_write_data_data_mux1h_4_rmff , weight_write_data_data_mux1h_3_rmff
      , weight_write_data_data_mux1h_2_rmff , weight_write_data_data_mux1h_1_rmff
      , weight_write_data_data_mux1h_rmff};
  assign weight_mem_banks_bank_array_impl_data5_rsci_radr_d = MUX_v_12_16_2(weight_read_addrs_0_15_4_lpi_1_dfm_5_mx0,
      (weight_read_addrs_1_lpi_1_dfm_2[15:4]), (weight_read_addrs_2_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_3_lpi_1_dfm_2[15:4]), (weight_read_addrs_4_15_2_lpi_1_dfm_2[13:2]),
      (weight_read_addrs_5_lpi_1_dfm_2[15:4]), (weight_read_addrs_6_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_7_lpi_1_dfm_2[15:4]), (weight_read_addrs_8_15_3_lpi_1_dfm_3[12:1]),
      (weight_read_addrs_9_lpi_1_dfm_3[15:4]), (weight_read_addrs_10_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_11_lpi_1_dfm_3[15:4]), (weight_read_addrs_12_15_2_lpi_1_dfm_3[13:2]),
      (weight_read_addrs_13_lpi_1_dfm_3[15:4]), (weight_read_addrs_14_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_15_lpi_1_dfm_3[15:4]), {weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_8_2_sva_1 , weight_mem_read_arbxbar_xbar_for_3_source_local_8_1_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_8_0_sva_1});
  assign weight_mem_banks_bank_array_impl_data5_rsci_we_d_pff = and_3019_cse;
  assign weight_mem_banks_bank_array_impl_data5_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = or_1425_cse;
  assign weight_mem_banks_bank_array_impl_data6_rsci_d_d = {while_while_and_18_itm
      , weight_write_data_data_mux1h_14_rmff , weight_write_data_data_mux1h_13_rmff
      , weight_write_data_data_mux1h_12_rmff , weight_write_data_data_mux1h_11_rmff
      , weight_write_data_data_mux1h_10_rmff , weight_write_data_data_mux1h_9_rmff
      , weight_write_data_data_mux1h_8_rmff , weight_write_data_data_mux1h_7_rmff
      , weight_write_data_data_mux1h_6_rmff , weight_write_data_data_mux1h_5_rmff
      , weight_write_data_data_mux1h_4_rmff , weight_write_data_data_mux1h_3_rmff
      , weight_write_data_data_mux1h_2_rmff , weight_write_data_data_mux1h_1_rmff
      , weight_write_data_data_mux1h_rmff};
  assign weight_mem_banks_bank_array_impl_data6_rsci_radr_d = MUX_v_12_16_2(weight_read_addrs_0_15_4_lpi_1_dfm_5_mx0,
      (weight_read_addrs_1_lpi_1_dfm_2[15:4]), (weight_read_addrs_2_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_3_lpi_1_dfm_2[15:4]), (weight_read_addrs_4_15_2_lpi_1_dfm_2[13:2]),
      (weight_read_addrs_5_lpi_1_dfm_2[15:4]), (weight_read_addrs_6_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_7_lpi_1_dfm_2[15:4]), (weight_read_addrs_8_15_3_lpi_1_dfm_3[12:1]),
      (weight_read_addrs_9_lpi_1_dfm_3[15:4]), (weight_read_addrs_10_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_11_lpi_1_dfm_3[15:4]), (weight_read_addrs_12_15_2_lpi_1_dfm_3[13:2]),
      (weight_read_addrs_13_lpi_1_dfm_3[15:4]), (weight_read_addrs_14_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_15_lpi_1_dfm_3[15:4]), {weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_9_2_sva_1 , weight_mem_read_arbxbar_xbar_for_3_source_local_9_1_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_9_0_sva_1});
  assign weight_mem_banks_bank_array_impl_data6_rsci_we_d_pff = and_3015_cse;
  assign weight_mem_banks_bank_array_impl_data6_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = or_1429_cse;
  assign weight_mem_banks_bank_array_impl_data7_rsci_d_d = {while_while_and_18_itm
      , weight_write_data_data_mux1h_14_rmff , weight_write_data_data_mux1h_13_rmff
      , weight_write_data_data_mux1h_12_rmff , weight_write_data_data_mux1h_11_rmff
      , weight_write_data_data_mux1h_10_rmff , weight_write_data_data_mux1h_9_rmff
      , weight_write_data_data_mux1h_8_rmff , weight_write_data_data_mux1h_7_rmff
      , weight_write_data_data_mux1h_6_rmff , weight_write_data_data_mux1h_5_rmff
      , weight_write_data_data_mux1h_4_rmff , weight_write_data_data_mux1h_3_rmff
      , weight_write_data_data_mux1h_2_rmff , weight_write_data_data_mux1h_1_rmff
      , weight_write_data_data_mux1h_rmff};
  assign weight_mem_banks_bank_array_impl_data7_rsci_radr_d = MUX_v_12_16_2(weight_read_addrs_0_15_4_lpi_1_dfm_5_mx0,
      (weight_read_addrs_1_lpi_1_dfm_2[15:4]), (weight_read_addrs_2_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_3_lpi_1_dfm_2[15:4]), (weight_read_addrs_4_15_2_lpi_1_dfm_2[13:2]),
      (weight_read_addrs_5_lpi_1_dfm_2[15:4]), (weight_read_addrs_6_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_7_lpi_1_dfm_2[15:4]), (weight_read_addrs_8_15_3_lpi_1_dfm_3[12:1]),
      (weight_read_addrs_9_lpi_1_dfm_3[15:4]), (weight_read_addrs_10_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_11_lpi_1_dfm_3[15:4]), (weight_read_addrs_12_15_2_lpi_1_dfm_3[13:2]),
      (weight_read_addrs_13_lpi_1_dfm_3[15:4]), (weight_read_addrs_14_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_15_lpi_1_dfm_3[15:4]), {weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_10_2_sva_1 , weight_mem_read_arbxbar_xbar_for_3_source_local_10_1_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_10_0_sva_1});
  assign weight_mem_banks_bank_array_impl_data7_rsci_we_d_pff = and_3011_cse;
  assign weight_mem_banks_bank_array_impl_data7_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = or_1433_cse;
  assign weight_mem_banks_bank_array_impl_data8_rsci_d_d = {while_while_and_18_itm
      , weight_write_data_data_mux1h_14_rmff , weight_write_data_data_mux1h_13_rmff
      , weight_write_data_data_mux1h_12_rmff , weight_write_data_data_mux1h_11_rmff
      , weight_write_data_data_mux1h_10_rmff , weight_write_data_data_mux1h_9_rmff
      , weight_write_data_data_mux1h_8_rmff , weight_write_data_data_mux1h_7_rmff
      , weight_write_data_data_mux1h_6_rmff , weight_write_data_data_mux1h_5_rmff
      , weight_write_data_data_mux1h_4_rmff , weight_write_data_data_mux1h_3_rmff
      , weight_write_data_data_mux1h_2_rmff , weight_write_data_data_mux1h_1_rmff
      , weight_write_data_data_mux1h_rmff};
  assign weight_mem_banks_bank_array_impl_data8_rsci_radr_d = MUX_v_12_16_2(weight_read_addrs_0_15_4_lpi_1_dfm_5_mx0,
      (weight_read_addrs_1_lpi_1_dfm_2[15:4]), (weight_read_addrs_2_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_3_lpi_1_dfm_2[15:4]), (weight_read_addrs_4_15_2_lpi_1_dfm_2[13:2]),
      (weight_read_addrs_5_lpi_1_dfm_2[15:4]), (weight_read_addrs_6_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_7_lpi_1_dfm_2[15:4]), (weight_read_addrs_8_15_3_lpi_1_dfm_3[12:1]),
      (weight_read_addrs_9_lpi_1_dfm_3[15:4]), (weight_read_addrs_10_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_11_lpi_1_dfm_3[15:4]), (weight_read_addrs_12_15_2_lpi_1_dfm_3[13:2]),
      (weight_read_addrs_13_lpi_1_dfm_3[15:4]), (weight_read_addrs_14_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_15_lpi_1_dfm_3[15:4]), {weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_11_2_sva_1 , weight_mem_read_arbxbar_xbar_for_3_source_local_11_1_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_11_0_sva_1});
  assign weight_mem_banks_bank_array_impl_data8_rsci_we_d_pff = and_3007_cse;
  assign weight_mem_banks_bank_array_impl_data8_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = or_1437_cse;
  assign weight_mem_banks_bank_array_impl_data9_rsci_d_d = {while_while_and_18_itm
      , weight_write_data_data_mux1h_14_rmff , weight_write_data_data_mux1h_13_rmff
      , weight_write_data_data_mux1h_12_rmff , weight_write_data_data_mux1h_11_rmff
      , weight_write_data_data_mux1h_10_rmff , weight_write_data_data_mux1h_9_rmff
      , weight_write_data_data_mux1h_8_rmff , weight_write_data_data_mux1h_7_rmff
      , weight_write_data_data_mux1h_6_rmff , weight_write_data_data_mux1h_5_rmff
      , weight_write_data_data_mux1h_4_rmff , weight_write_data_data_mux1h_3_rmff
      , weight_write_data_data_mux1h_2_rmff , weight_write_data_data_mux1h_1_rmff
      , weight_write_data_data_mux1h_rmff};
  assign weight_mem_banks_bank_array_impl_data9_rsci_radr_d = MUX_v_12_16_2(weight_read_addrs_0_15_4_lpi_1_dfm_5_mx0,
      (weight_read_addrs_1_lpi_1_dfm_2[15:4]), (weight_read_addrs_2_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_3_lpi_1_dfm_2[15:4]), (weight_read_addrs_4_15_2_lpi_1_dfm_2[13:2]),
      (weight_read_addrs_5_lpi_1_dfm_2[15:4]), (weight_read_addrs_6_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_7_lpi_1_dfm_2[15:4]), (weight_read_addrs_8_15_3_lpi_1_dfm_3[12:1]),
      (weight_read_addrs_9_lpi_1_dfm_3[15:4]), (weight_read_addrs_10_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_11_lpi_1_dfm_3[15:4]), (weight_read_addrs_12_15_2_lpi_1_dfm_3[13:2]),
      (weight_read_addrs_13_lpi_1_dfm_3[15:4]), (weight_read_addrs_14_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_15_lpi_1_dfm_3[15:4]), {weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_12_2_sva_1 , weight_mem_read_arbxbar_xbar_for_3_source_local_12_1_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_12_0_sva_1});
  assign weight_mem_banks_bank_array_impl_data9_rsci_we_d_pff = and_3003_cse;
  assign weight_mem_banks_bank_array_impl_data9_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = or_1441_cse;
  assign weight_mem_banks_bank_array_impl_data10_rsci_d_d = {while_while_and_18_itm
      , weight_write_data_data_mux1h_14_rmff , weight_write_data_data_mux1h_13_rmff
      , weight_write_data_data_mux1h_12_rmff , weight_write_data_data_mux1h_11_rmff
      , weight_write_data_data_mux1h_10_rmff , weight_write_data_data_mux1h_9_rmff
      , weight_write_data_data_mux1h_8_rmff , weight_write_data_data_mux1h_7_rmff
      , weight_write_data_data_mux1h_6_rmff , weight_write_data_data_mux1h_5_rmff
      , weight_write_data_data_mux1h_4_rmff , weight_write_data_data_mux1h_3_rmff
      , weight_write_data_data_mux1h_2_rmff , weight_write_data_data_mux1h_1_rmff
      , weight_write_data_data_mux1h_rmff};
  assign weight_mem_banks_bank_array_impl_data10_rsci_radr_d = MUX_v_12_16_2(weight_read_addrs_0_15_4_lpi_1_dfm_5_mx0,
      (weight_read_addrs_1_lpi_1_dfm_2[15:4]), (weight_read_addrs_2_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_3_lpi_1_dfm_2[15:4]), (weight_read_addrs_4_15_2_lpi_1_dfm_2[13:2]),
      (weight_read_addrs_5_lpi_1_dfm_2[15:4]), (weight_read_addrs_6_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_7_lpi_1_dfm_2[15:4]), (weight_read_addrs_8_15_3_lpi_1_dfm_3[12:1]),
      (weight_read_addrs_9_lpi_1_dfm_3[15:4]), (weight_read_addrs_10_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_11_lpi_1_dfm_3[15:4]), (weight_read_addrs_12_15_2_lpi_1_dfm_3[13:2]),
      (weight_read_addrs_13_lpi_1_dfm_3[15:4]), (weight_read_addrs_14_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_15_lpi_1_dfm_3[15:4]), {weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_13_2_sva_1 , weight_mem_read_arbxbar_xbar_for_3_source_local_13_1_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_13_0_sva_1});
  assign weight_mem_banks_bank_array_impl_data10_rsci_we_d_pff = and_2999_cse;
  assign weight_mem_banks_bank_array_impl_data10_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = or_1445_cse;
  assign weight_mem_banks_bank_array_impl_data11_rsci_d_d = {while_while_and_18_itm
      , weight_write_data_data_mux1h_14_rmff , weight_write_data_data_mux1h_13_rmff
      , weight_write_data_data_mux1h_12_rmff , weight_write_data_data_mux1h_11_rmff
      , weight_write_data_data_mux1h_10_rmff , weight_write_data_data_mux1h_9_rmff
      , weight_write_data_data_mux1h_8_rmff , weight_write_data_data_mux1h_7_rmff
      , weight_write_data_data_mux1h_6_rmff , weight_write_data_data_mux1h_5_rmff
      , weight_write_data_data_mux1h_4_rmff , weight_write_data_data_mux1h_3_rmff
      , weight_write_data_data_mux1h_2_rmff , weight_write_data_data_mux1h_1_rmff
      , weight_write_data_data_mux1h_rmff};
  assign weight_mem_banks_bank_array_impl_data11_rsci_radr_d = MUX_v_12_16_2(weight_read_addrs_0_15_4_lpi_1_dfm_5_mx0,
      (weight_read_addrs_1_lpi_1_dfm_2[15:4]), (weight_read_addrs_2_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_3_lpi_1_dfm_2[15:4]), (weight_read_addrs_4_15_2_lpi_1_dfm_2[13:2]),
      (weight_read_addrs_5_lpi_1_dfm_2[15:4]), (weight_read_addrs_6_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_7_lpi_1_dfm_2[15:4]), (weight_read_addrs_8_15_3_lpi_1_dfm_3[12:1]),
      (weight_read_addrs_9_lpi_1_dfm_3[15:4]), (weight_read_addrs_10_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_11_lpi_1_dfm_3[15:4]), (weight_read_addrs_12_15_2_lpi_1_dfm_3[13:2]),
      (weight_read_addrs_13_lpi_1_dfm_3[15:4]), (weight_read_addrs_14_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_15_lpi_1_dfm_3[15:4]), {weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_14_2_sva_1 , weight_mem_read_arbxbar_xbar_for_3_source_local_14_1_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_14_0_sva_1});
  assign weight_mem_banks_bank_array_impl_data11_rsci_we_d_pff = and_2995_cse;
  assign weight_mem_banks_bank_array_impl_data11_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = or_1449_cse;
  assign weight_mem_banks_bank_array_impl_data12_rsci_d_d = {while_while_and_18_itm
      , weight_write_data_data_mux1h_14_rmff , weight_write_data_data_mux1h_13_rmff
      , weight_write_data_data_mux1h_12_rmff , weight_write_data_data_mux1h_11_rmff
      , weight_write_data_data_mux1h_10_rmff , weight_write_data_data_mux1h_9_rmff
      , weight_write_data_data_mux1h_8_rmff , weight_write_data_data_mux1h_7_rmff
      , weight_write_data_data_mux1h_6_rmff , weight_write_data_data_mux1h_5_rmff
      , weight_write_data_data_mux1h_4_rmff , weight_write_data_data_mux1h_3_rmff
      , weight_write_data_data_mux1h_2_rmff , weight_write_data_data_mux1h_1_rmff
      , weight_write_data_data_mux1h_rmff};
  assign weight_mem_banks_bank_array_impl_data12_rsci_radr_d = MUX_v_12_16_2(weight_read_addrs_0_15_4_lpi_1_dfm_5_mx0,
      (weight_read_addrs_1_lpi_1_dfm_2[15:4]), (weight_read_addrs_2_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_3_lpi_1_dfm_2[15:4]), (weight_read_addrs_4_15_2_lpi_1_dfm_2[13:2]),
      (weight_read_addrs_5_lpi_1_dfm_2[15:4]), (weight_read_addrs_6_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_7_lpi_1_dfm_2[15:4]), (weight_read_addrs_8_15_3_lpi_1_dfm_3[12:1]),
      (weight_read_addrs_9_lpi_1_dfm_3[15:4]), (weight_read_addrs_10_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_11_lpi_1_dfm_3[15:4]), (weight_read_addrs_12_15_2_lpi_1_dfm_3[13:2]),
      (weight_read_addrs_13_lpi_1_dfm_3[15:4]), (weight_read_addrs_14_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_15_lpi_1_dfm_3[15:4]), {weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_15_2_sva_1 , weight_mem_read_arbxbar_xbar_for_3_source_local_15_1_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_15_0_sva_1});
  assign weight_mem_banks_bank_array_impl_data12_rsci_we_d_pff = and_2991_cse;
  assign weight_mem_banks_bank_array_impl_data12_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = or_1453_cse;
  assign weight_mem_banks_bank_array_impl_data13_rsci_d_d = {while_while_and_18_itm
      , weight_write_data_data_mux1h_14_rmff , weight_write_data_data_mux1h_13_rmff
      , weight_write_data_data_mux1h_12_rmff , weight_write_data_data_mux1h_11_rmff
      , weight_write_data_data_mux1h_10_rmff , weight_write_data_data_mux1h_9_rmff
      , weight_write_data_data_mux1h_8_rmff , weight_write_data_data_mux1h_7_rmff
      , weight_write_data_data_mux1h_6_rmff , weight_write_data_data_mux1h_5_rmff
      , weight_write_data_data_mux1h_4_rmff , weight_write_data_data_mux1h_3_rmff
      , weight_write_data_data_mux1h_2_rmff , weight_write_data_data_mux1h_1_rmff
      , weight_write_data_data_mux1h_rmff};
  assign weight_mem_banks_bank_array_impl_data13_rsci_radr_d = MUX_v_12_16_2(weight_read_addrs_0_15_4_lpi_1_dfm_5_mx0,
      (weight_read_addrs_1_lpi_1_dfm_2[15:4]), (weight_read_addrs_2_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_3_lpi_1_dfm_2[15:4]), (weight_read_addrs_4_15_2_lpi_1_dfm_2[13:2]),
      (weight_read_addrs_5_lpi_1_dfm_2[15:4]), (weight_read_addrs_6_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_7_lpi_1_dfm_2[15:4]), (weight_read_addrs_8_15_3_lpi_1_dfm_3[12:1]),
      (weight_read_addrs_9_lpi_1_dfm_3[15:4]), (weight_read_addrs_10_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_11_lpi_1_dfm_3[15:4]), (weight_read_addrs_12_15_2_lpi_1_dfm_3[13:2]),
      (weight_read_addrs_13_lpi_1_dfm_3[15:4]), (weight_read_addrs_14_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_15_lpi_1_dfm_3[15:4]), {weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_16_2_sva_1 , weight_mem_read_arbxbar_xbar_for_3_source_local_16_1_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_16_0_sva_1});
  assign weight_mem_banks_bank_array_impl_data13_rsci_we_d_pff = and_2987_cse;
  assign weight_mem_banks_bank_array_impl_data13_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = or_1457_cse;
  assign weight_mem_banks_bank_array_impl_data14_rsci_d_d = {while_while_and_18_itm
      , weight_write_data_data_mux1h_14_rmff , weight_write_data_data_mux1h_13_rmff
      , weight_write_data_data_mux1h_12_rmff , weight_write_data_data_mux1h_11_rmff
      , weight_write_data_data_mux1h_10_rmff , weight_write_data_data_mux1h_9_rmff
      , weight_write_data_data_mux1h_8_rmff , weight_write_data_data_mux1h_7_rmff
      , weight_write_data_data_mux1h_6_rmff , weight_write_data_data_mux1h_5_rmff
      , weight_write_data_data_mux1h_4_rmff , weight_write_data_data_mux1h_3_rmff
      , weight_write_data_data_mux1h_2_rmff , weight_write_data_data_mux1h_1_rmff
      , weight_write_data_data_mux1h_rmff};
  assign weight_mem_banks_bank_array_impl_data14_rsci_radr_d = MUX_v_12_16_2(weight_read_addrs_0_15_4_lpi_1_dfm_5_mx0,
      (weight_read_addrs_1_lpi_1_dfm_2[15:4]), (weight_read_addrs_2_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_3_lpi_1_dfm_2[15:4]), (weight_read_addrs_4_15_2_lpi_1_dfm_2[13:2]),
      (weight_read_addrs_5_lpi_1_dfm_2[15:4]), (weight_read_addrs_6_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_7_lpi_1_dfm_2[15:4]), (weight_read_addrs_8_15_3_lpi_1_dfm_3[12:1]),
      (weight_read_addrs_9_lpi_1_dfm_3[15:4]), (weight_read_addrs_10_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_11_lpi_1_dfm_3[15:4]), (weight_read_addrs_12_15_2_lpi_1_dfm_3[13:2]),
      (weight_read_addrs_13_lpi_1_dfm_3[15:4]), (weight_read_addrs_14_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_15_lpi_1_dfm_3[15:4]), {weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_17_2_sva_1 , weight_mem_read_arbxbar_xbar_for_3_source_local_17_1_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_17_0_sva_1});
  assign weight_mem_banks_bank_array_impl_data14_rsci_we_d_pff = and_2983_cse;
  assign weight_mem_banks_bank_array_impl_data14_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = or_1461_cse;
  assign weight_mem_banks_bank_array_impl_data15_rsci_d_d = {while_while_and_18_itm
      , weight_write_data_data_mux1h_14_rmff , weight_write_data_data_mux1h_13_rmff
      , weight_write_data_data_mux1h_12_rmff , weight_write_data_data_mux1h_11_rmff
      , weight_write_data_data_mux1h_10_rmff , weight_write_data_data_mux1h_9_rmff
      , weight_write_data_data_mux1h_8_rmff , weight_write_data_data_mux1h_7_rmff
      , weight_write_data_data_mux1h_6_rmff , weight_write_data_data_mux1h_5_rmff
      , weight_write_data_data_mux1h_4_rmff , weight_write_data_data_mux1h_3_rmff
      , weight_write_data_data_mux1h_2_rmff , weight_write_data_data_mux1h_1_rmff
      , weight_write_data_data_mux1h_rmff};
  assign weight_mem_banks_bank_array_impl_data15_rsci_radr_d = MUX_v_12_16_2(weight_read_addrs_0_15_4_lpi_1_dfm_5_mx0,
      (weight_read_addrs_1_lpi_1_dfm_2[15:4]), (weight_read_addrs_2_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_3_lpi_1_dfm_2[15:4]), (weight_read_addrs_4_15_2_lpi_1_dfm_2[13:2]),
      (weight_read_addrs_5_lpi_1_dfm_2[15:4]), (weight_read_addrs_6_15_1_lpi_1_dfm_2[14:3]),
      (weight_read_addrs_7_lpi_1_dfm_2[15:4]), (weight_read_addrs_8_15_3_lpi_1_dfm_3[12:1]),
      (weight_read_addrs_9_lpi_1_dfm_3[15:4]), (weight_read_addrs_10_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_11_lpi_1_dfm_3[15:4]), (weight_read_addrs_12_15_2_lpi_1_dfm_3[13:2]),
      (weight_read_addrs_13_lpi_1_dfm_3[15:4]), (weight_read_addrs_14_15_1_lpi_1_dfm_3[14:3]),
      (weight_read_addrs_15_lpi_1_dfm_3[15:4]), {weight_mem_read_arbxbar_xbar_for_3_source_local_2_3_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_2_2_sva_1 , weight_mem_read_arbxbar_xbar_for_3_source_local_2_1_sva_1
      , weight_mem_read_arbxbar_xbar_for_3_source_local_2_0_sva_1});
  assign weight_mem_banks_bank_array_impl_data15_rsci_we_d_pff = and_2979_cse;
  assign weight_mem_banks_bank_array_impl_data15_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = or_1465_cse;
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_36_nl
      = (input_port_PopNB_mioi_idat_mxwt[127:120]) & ({{7{input_port_PopNB_mioi_ivld_mxwt}},
      input_port_PopNB_mioi_ivld_mxwt}) & ({{7{PECore_RunFSM_switch_lp_equal_tmp_3}},
      PECore_RunFSM_switch_lp_equal_tmp_3});
  assign while_mux_111_nl = MUX_v_8_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_36_nl,
      (rva_in_PopNB_mio_mrgout_dat_sva_1[127:120]), while_and_127_cse_1);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_35_nl
      = (input_port_PopNB_mioi_idat_mxwt[119:112]) & ({{7{input_port_PopNB_mioi_ivld_mxwt}},
      input_port_PopNB_mioi_ivld_mxwt}) & ({{7{PECore_RunFSM_switch_lp_equal_tmp_3}},
      PECore_RunFSM_switch_lp_equal_tmp_3});
  assign while_mux_110_nl = MUX_v_8_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_35_nl,
      (rva_in_PopNB_mio_mrgout_dat_sva_1[119:112]), while_and_127_cse_1);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_34_nl
      = (input_port_PopNB_mioi_idat_mxwt[111:104]) & ({{7{input_port_PopNB_mioi_ivld_mxwt}},
      input_port_PopNB_mioi_ivld_mxwt}) & ({{7{PECore_RunFSM_switch_lp_equal_tmp_3}},
      PECore_RunFSM_switch_lp_equal_tmp_3});
  assign while_mux_109_nl = MUX_v_8_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_34_nl,
      (rva_in_PopNB_mio_mrgout_dat_sva_1[111:104]), while_and_127_cse_1);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_33_nl
      = (input_port_PopNB_mioi_idat_mxwt[103:96]) & ({{7{input_port_PopNB_mioi_ivld_mxwt}},
      input_port_PopNB_mioi_ivld_mxwt}) & ({{7{PECore_RunFSM_switch_lp_equal_tmp_3}},
      PECore_RunFSM_switch_lp_equal_tmp_3});
  assign while_mux_108_nl = MUX_v_8_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_33_nl,
      (rva_in_PopNB_mio_mrgout_dat_sva_1[103:96]), while_and_127_cse_1);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_32_nl
      = (input_port_PopNB_mioi_idat_mxwt[95:88]) & ({{7{input_port_PopNB_mioi_ivld_mxwt}},
      input_port_PopNB_mioi_ivld_mxwt}) & ({{7{PECore_RunFSM_switch_lp_equal_tmp_3}},
      PECore_RunFSM_switch_lp_equal_tmp_3});
  assign while_mux_107_nl = MUX_v_8_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_32_nl,
      (rva_in_PopNB_mio_mrgout_dat_sva_1[95:88]), while_and_127_cse_1);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_31_nl
      = (input_port_PopNB_mioi_idat_mxwt[87:80]) & ({{7{input_port_PopNB_mioi_ivld_mxwt}},
      input_port_PopNB_mioi_ivld_mxwt}) & ({{7{PECore_RunFSM_switch_lp_equal_tmp_3}},
      PECore_RunFSM_switch_lp_equal_tmp_3});
  assign while_mux_106_nl = MUX_v_8_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_31_nl,
      (rva_in_PopNB_mio_mrgout_dat_sva_1[87:80]), while_and_127_cse_1);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_30_nl
      = (input_port_PopNB_mioi_idat_mxwt[79:72]) & ({{7{input_port_PopNB_mioi_ivld_mxwt}},
      input_port_PopNB_mioi_ivld_mxwt}) & ({{7{PECore_RunFSM_switch_lp_equal_tmp_3}},
      PECore_RunFSM_switch_lp_equal_tmp_3});
  assign while_mux_105_nl = MUX_v_8_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_30_nl,
      (rva_in_PopNB_mio_mrgout_dat_sva_1[79:72]), while_and_127_cse_1);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_29_nl
      = (input_port_PopNB_mioi_idat_mxwt[71:64]) & ({{7{input_port_PopNB_mioi_ivld_mxwt}},
      input_port_PopNB_mioi_ivld_mxwt}) & ({{7{PECore_RunFSM_switch_lp_equal_tmp_3}},
      PECore_RunFSM_switch_lp_equal_tmp_3});
  assign while_mux_104_nl = MUX_v_8_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_29_nl,
      (rva_in_PopNB_mio_mrgout_dat_sva_1[71:64]), while_and_127_cse_1);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_28_nl
      = (input_port_PopNB_mioi_idat_mxwt[63:56]) & ({{7{input_port_PopNB_mioi_ivld_mxwt}},
      input_port_PopNB_mioi_ivld_mxwt}) & ({{7{PECore_RunFSM_switch_lp_equal_tmp_3}},
      PECore_RunFSM_switch_lp_equal_tmp_3});
  assign while_mux_103_nl = MUX_v_8_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_28_nl,
      (rva_in_PopNB_mio_mrgout_dat_sva_1[63:56]), while_and_127_cse_1);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_27_nl
      = (input_port_PopNB_mioi_idat_mxwt[55:48]) & ({{7{input_port_PopNB_mioi_ivld_mxwt}},
      input_port_PopNB_mioi_ivld_mxwt}) & ({{7{PECore_RunFSM_switch_lp_equal_tmp_3}},
      PECore_RunFSM_switch_lp_equal_tmp_3});
  assign while_mux_102_nl = MUX_v_8_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_27_nl,
      (rva_in_PopNB_mio_mrgout_dat_sva_1[55:48]), while_and_127_cse_1);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_26_nl
      = (input_port_PopNB_mioi_idat_mxwt[47:40]) & ({{7{input_port_PopNB_mioi_ivld_mxwt}},
      input_port_PopNB_mioi_ivld_mxwt}) & ({{7{PECore_RunFSM_switch_lp_equal_tmp_3}},
      PECore_RunFSM_switch_lp_equal_tmp_3});
  assign while_mux_101_nl = MUX_v_8_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_26_nl,
      (rva_in_PopNB_mio_mrgout_dat_sva_1[47:40]), while_and_127_cse_1);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_25_nl
      = (input_port_PopNB_mioi_idat_mxwt[39:32]) & ({{7{input_port_PopNB_mioi_ivld_mxwt}},
      input_port_PopNB_mioi_ivld_mxwt}) & ({{7{PECore_RunFSM_switch_lp_equal_tmp_3}},
      PECore_RunFSM_switch_lp_equal_tmp_3});
  assign while_mux_100_nl = MUX_v_8_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_25_nl,
      (rva_in_PopNB_mio_mrgout_dat_sva_1[39:32]), while_and_127_cse_1);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_24_nl
      = (input_port_PopNB_mioi_idat_mxwt[31:24]) & ({{7{input_port_PopNB_mioi_ivld_mxwt}},
      input_port_PopNB_mioi_ivld_mxwt}) & ({{7{PECore_RunFSM_switch_lp_equal_tmp_3}},
      PECore_RunFSM_switch_lp_equal_tmp_3});
  assign while_mux_99_nl = MUX_v_8_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_24_nl,
      (rva_in_PopNB_mio_mrgout_dat_sva_1[31:24]), while_and_127_cse_1);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_23_nl
      = (input_port_PopNB_mioi_idat_mxwt[23:16]) & ({{7{input_port_PopNB_mioi_ivld_mxwt}},
      input_port_PopNB_mioi_ivld_mxwt}) & ({{7{PECore_RunFSM_switch_lp_equal_tmp_3}},
      PECore_RunFSM_switch_lp_equal_tmp_3});
  assign while_mux_98_nl = MUX_v_8_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_23_nl,
      (rva_in_PopNB_mio_mrgout_dat_sva_1[23:16]), while_and_127_cse_1);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_22_nl
      = (input_port_PopNB_mioi_idat_mxwt[15:8]) & ({{7{input_port_PopNB_mioi_ivld_mxwt}},
      input_port_PopNB_mioi_ivld_mxwt}) & ({{7{PECore_RunFSM_switch_lp_equal_tmp_3}},
      PECore_RunFSM_switch_lp_equal_tmp_3});
  assign while_mux_97_nl = MUX_v_8_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_22_nl,
      (rva_in_PopNB_mio_mrgout_dat_sva_1[15:8]), while_and_127_cse_1);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_21_nl
      = (input_port_PopNB_mioi_idat_mxwt[7:0]) & ({{7{input_port_PopNB_mioi_ivld_mxwt}},
      input_port_PopNB_mioi_ivld_mxwt}) & ({{7{PECore_RunFSM_switch_lp_equal_tmp_3}},
      PECore_RunFSM_switch_lp_equal_tmp_3});
  assign while_mux_96_nl = MUX_v_8_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_21_nl,
      (rva_in_PopNB_mio_mrgout_dat_sva_1[7:0]), while_and_127_cse_1);
  assign input_mem_banks_bank_array_impl_data0_rsci_d_d = {while_mux_111_nl , while_mux_110_nl
      , while_mux_109_nl , while_mux_108_nl , while_mux_107_nl , while_mux_106_nl
      , while_mux_105_nl , while_mux_104_nl , while_mux_103_nl , while_mux_102_nl
      , while_mux_101_nl , while_mux_100_nl , while_mux_99_nl , while_mux_98_nl ,
      while_mux_97_nl , while_mux_96_nl};
  assign or_1593_cse = nand_199_cse | (rva_in_PopNB_mioi_idat_mxwt[151]) | (~ (rva_in_PopNB_mioi_idat_mxwt[149]))
      | (rva_in_PopNB_mioi_idat_mxwt[148]) | is_start_sva;
  assign and_tmp = or_1593_cse & (~(PECore_RunFSM_switch_lp_nor_3_cse_1 & (pe_config_is_bias_sva
      | (~ PECore_RunFSM_switch_lp_equal_tmp_4))));
  assign nl_PEManager_16U_GetInputAddr_1_acc_nl = pe_config_input_counter_sva + z_out_41;
  assign PEManager_16U_GetInputAddr_1_acc_nl = nl_PEManager_16U_GetInputAddr_1_acc_nl[7:0];
  assign nl_PEManager_16U_GetBiasAddr_acc_nl = pe_config_output_counter_sva + z_out_41;
  assign PEManager_16U_GetBiasAddr_acc_nl = nl_PEManager_16U_GetBiasAddr_acc_nl[7:0];
  assign PECore_DecodeAxi_if_and_nl = (~ PECore_RunFSM_switch_lp_equal_tmp_4) & or_1593_cse
      & (~ and_tmp);
  assign PECore_DecodeAxi_if_and_1_nl = PECore_RunFSM_switch_lp_equal_tmp_4 & or_1593_cse
      & (~ and_tmp);
  assign mux1h_7_nl = MUX1HOT_v_8_3_2((rva_in_PopNB_mio_mrgout_dat_sva_1[139:132]),
      PEManager_16U_GetInputAddr_1_acc_nl, PEManager_16U_GetBiasAddr_acc_nl, {(~
      or_1593_cse) , PECore_DecodeAxi_if_and_nl , PECore_DecodeAxi_if_and_1_nl});
  assign not_3760_nl = ~ and_tmp;
  assign input_mem_banks_bank_array_impl_data0_rsci_radr_d = MUX_v_8_2_2(8'b00000000,
      mux1h_7_nl, not_3760_nl);
  assign nl_PEManager_16U_GetInputAddr_acc_nl = (input_port_PopNB_mioi_idat_mxwt[136:129])
      + z_out_41;
  assign PEManager_16U_GetInputAddr_acc_nl = nl_PEManager_16U_GetInputAddr_acc_nl[7:0];
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_35_nl = PEManager_16U_GetInputAddr_acc_nl
      & ({{7{input_port_PopNB_mioi_ivld_mxwt}}, input_port_PopNB_mioi_ivld_mxwt})
      & ({{7{PECore_RunFSM_switch_lp_equal_tmp_3}}, PECore_RunFSM_switch_lp_equal_tmp_3});
  assign or_1589_nl = nand_199_cse | (rva_in_PopNB_mioi_idat_mxwt[151]) | (~ (rva_in_PopNB_mioi_idat_mxwt[149]))
      | or_dcpl_286;
  assign input_mem_banks_bank_array_impl_data0_rsci_wadr_d = MUX_v_8_2_2((rva_in_PopNB_mio_mrgout_dat_sva_1[139:132]),
      PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_35_nl, or_1589_nl);
  assign and_1488_nl = or_55_cse & or_1584_cse;
  assign mux_601_nl = MUX_s_1_2_2(and_1488_nl, or_55_cse, is_start_sva);
  assign input_mem_banks_bank_array_impl_data0_rsci_we_d_pff = (~ mux_601_nl) & (fsm_output[1]);
  assign input_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = and_2973_cse;
  assign or_dcpl_717 = (PECore_PushAxiRsp_if_and_45_cse & PECore_DecodeAxiRead_switch_lp_nor_10_cse_1
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_5) | (or_tmp_545 & PECore_PushAxiRsp_if_asn_70);
  assign or_dcpl_718 = ~((PECore_UpdateFSM_switch_lp_equal_tmp_1 | while_and_30_itm_1)
      & while_stage_0_2);
  assign or_dcpl_724 = or_dcpl_375 | PECore_DecodeAxiWrite_case_4_switch_lp_or_6_cse_1;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2 = (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_1_lpi_1_dfm_mx0)
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_1_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_1_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_1_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_1_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_1_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_1_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_1_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0 = ~(nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_1_lpi_1_dfm_mx0
      | nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_1_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_1_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_1_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_1_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_1_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_1_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_1_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_1_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_1_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_1_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_1_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_1_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_1_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_1_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_1_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_1_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_1_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_1_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_1_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_1_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_1_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_1 = (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_2_lpi_1_dfm_mx0)
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_2_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_1
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_2_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_1
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_2_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_1 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_2_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_2_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_1
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_2_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_1
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_2_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_1 = ~(nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_2_lpi_1_dfm_mx0
      | nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_2_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_1
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_2_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_1
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_2_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_1 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_2_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_1
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_2_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_1
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_2_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_1
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_2_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_1
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_2_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_1
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_2_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_1
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_2_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_1
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_2_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_1
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_2_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_1
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_2_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_1
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_2_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_1
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_2_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_1
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_2_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_1
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_2_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_1
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_2_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_1
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_2_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_1
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_2_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_1 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_1
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_2_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_2 = (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_3_lpi_1_dfm_mx0)
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_2
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_2
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_2 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_3_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_2
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_2
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_2 = ~(nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_3_lpi_1_dfm_mx0
      | nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_2
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_2
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_2 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_2
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_2
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_2
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_2
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_2
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_2
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_2
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_2
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_2
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_2
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_2
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_2
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_2
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_2
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_2
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_2
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_2 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_2
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_3 = (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_4_lpi_1_dfm_mx0)
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_4_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_3
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_4_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_3
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_4_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_3 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_4_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_4_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_3
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_4_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_3
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_4_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_3 = ~(nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_4_lpi_1_dfm_mx0
      | nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_4_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_3
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_4_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_3
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_4_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_3 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_4_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_3
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_4_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_3
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_4_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_3
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_4_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_3
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_4_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_3
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_4_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_3
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_4_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_3
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_4_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_3
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_4_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_3
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_4_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_3
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_4_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_3
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_4_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_3
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_4_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_3
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_4_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_3
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_4_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_3
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_4_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_3
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_4_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_3 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_3
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_4_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_4 = (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_5_lpi_1_dfm_mx0)
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_5_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_4
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_5_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_4
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_5_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_4 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_5_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_5_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_4
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_5_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_4
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_5_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_4 = ~(nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_5_lpi_1_dfm_mx0
      | nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_5_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_4
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_5_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_4
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_5_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_4 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_5_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_4
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_5_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_4
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_5_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_4
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_5_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_4
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_5_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_4
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_5_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_4
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_5_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_4
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_5_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_4
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_5_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_4
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_5_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_4
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_5_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_4
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_5_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_4
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_5_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_4
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_5_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_4
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_5_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_4
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_5_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_4
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_5_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_4 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_4
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_5_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_5 = (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_6_lpi_1_dfm_mx0)
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_6_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_5
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_6_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_5
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_6_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_5 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_6_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_6_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_5
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_6_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_5
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_6_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_5 = ~(nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_6_lpi_1_dfm_mx0
      | nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_6_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_5
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_6_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_5
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_6_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_5 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_6_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_5
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_6_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_5
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_6_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_5
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_6_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_5
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_6_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_5
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_6_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_5
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_6_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_5
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_6_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_5
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_6_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_5
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_6_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_5
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_6_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_5
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_6_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_5
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_6_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_5
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_6_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_5
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_6_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_5
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_6_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_5
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_6_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_5 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_5
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_6_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_6 = (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_7_lpi_1_dfm_mx0)
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_7_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_6
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_7_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_6
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_7_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_6 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_7_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_7_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_6
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_7_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_6
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_7_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_6 = ~(nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_7_lpi_1_dfm_mx0
      | nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_7_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_6
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_7_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_6
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_7_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_6 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_7_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_6
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_7_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_6
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_7_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_6
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_7_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_6
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_7_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_6
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_7_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_6
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_7_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_6
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_7_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_6
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_7_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_6
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_7_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_6
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_7_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_6
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_7_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_6
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_7_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_6
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_7_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_6
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_7_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_6
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_7_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_6
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_7_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_6 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_6
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_7_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_7 = (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_8_lpi_1_dfm_mx0)
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_8_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_7
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_8_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_7
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_8_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_7 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_8_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_8_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_7
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_8_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_7
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_8_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_7 = ~(nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_8_lpi_1_dfm_mx0
      | nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_8_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_7
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_8_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_7
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_8_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_7 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_8_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_8_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_7
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_8_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_7
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_8_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_7
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_8_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_7
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_8_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_7
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_8_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_7
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_8_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_7
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_8_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_7
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_8_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_7
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_8_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_7
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_8_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_7
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_8_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_7
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_8_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_7
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_8_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_7
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_8_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_7
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_8_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_7
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_8_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_7 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_7
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_8_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_8 = (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_9_lpi_1_dfm_mx0)
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_9_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_8
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_9_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_8
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_9_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_8 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_9_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_9_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_8
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_9_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_8
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_9_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_8 = ~(nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_9_lpi_1_dfm_mx0
      | nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_9_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_8
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_9_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_8
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_9_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_8 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_9_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_9_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_8
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_9_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_8
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_9_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_8
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_9_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_8
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_9_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_8
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_9_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_8
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_9_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_8
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_9_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_8
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_9_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_8
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_9_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_8
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_9_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_8
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_9_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_8
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_9_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_8
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_9_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_8
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_9_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_8
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_9_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_8
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_9_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_8 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_8
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_9_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_9 = (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_10_lpi_1_dfm_mx0)
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_10_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_9
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_10_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_9
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_10_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_9 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_10_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_10_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_9
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_10_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_9
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_10_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_9 = ~(nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_10_lpi_1_dfm_mx0
      | nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_10_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_9
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_10_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_9
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_10_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_9 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_10_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_10_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_9
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_10_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_9
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_10_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_9
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_10_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_9
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_10_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_9
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_10_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_9
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_10_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_9
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_10_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_9
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_10_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_9
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_10_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_9
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_10_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_9
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_10_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_9
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_10_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_9
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_10_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_9
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_10_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_9
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_10_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_9
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_10_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_9 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_9
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_10_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_10 = (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_11_lpi_1_dfm_mx0)
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_11_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_10
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_11_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_10
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_11_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_10 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_11_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_11_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_10
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_11_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_10
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_11_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_10 = ~(nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_11_lpi_1_dfm_mx0
      | nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_11_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_10
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_11_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_10
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_11_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_10 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_11_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_11_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_10
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_11_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_10
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_11_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_10
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_11_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_10
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_11_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_10
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_11_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_10
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_11_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_10
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_11_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_10
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_11_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_10
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_11_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_10
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_11_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_10
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_11_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_10
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_11_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_10
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_11_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_10
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_11_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_10
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_11_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_10
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_11_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_10 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_10
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_11_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_11 = (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_12_lpi_1_dfm_mx0)
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_12_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_11
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_12_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_11
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_12_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_11 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_12_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_12_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_11
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_12_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_11
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_12_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_11 = ~(nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_12_lpi_1_dfm_mx0
      | nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_12_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_11
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_12_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_11
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_12_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_11 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_12_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_12_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_11
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_12_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_11
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_12_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_11
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_12_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_11
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_12_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_11
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_12_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_11
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_12_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_11
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_12_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_11
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_12_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_11
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_12_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_11
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_12_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_11
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_12_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_11
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_12_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_11
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_12_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_11
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_12_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_11
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_12_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_11
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_12_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_11 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_11
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_12_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_12 = (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_13_lpi_1_dfm_mx0)
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_13_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_12
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_13_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_12
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_13_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_12 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_13_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_13_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_12
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_13_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_12
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_13_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_12 = ~(nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_13_lpi_1_dfm_mx0
      | nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_13_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_12
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_13_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_12
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_13_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_12 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_13_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_13_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_12
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_13_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_12
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_13_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_12
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_13_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_12
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_13_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_12
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_13_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_12
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_13_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_12
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_13_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_12
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_13_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_12
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_13_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_12
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_13_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_12
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_13_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_12
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_13_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_12
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_13_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_12
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_13_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_12
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_13_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_12
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_13_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_12 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_12
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_13_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_13 = (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_14_lpi_1_dfm_mx0)
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_14_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_13
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_14_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_13
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_14_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_13 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_14_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_14_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_13
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_14_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_13
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_14_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_13 = ~(nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_14_lpi_1_dfm_mx0
      | nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_14_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_13
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_14_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_13
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_14_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_13 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_14_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_14_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_13
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_14_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_13
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_14_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_13
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_14_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_13
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_14_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_13
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_14_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_13
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_14_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_13
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_14_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_13
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_14_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_13
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_14_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_13
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_14_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_13
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_14_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_13
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_14_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_13
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_14_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_13
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_14_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_13
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_14_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_13
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_14_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_13 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_13
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_14_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_14 = (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_15_lpi_1_dfm_mx0)
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_15_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_14
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_15_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_14
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_15_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_14 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_15_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_15_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_14
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_15_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_14
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_15_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_14 = ~(nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_15_lpi_1_dfm_mx0
      | nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_15_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_14
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_15_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_14
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_15_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_14 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_15_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_15_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_14
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_15_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_14
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_15_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_14
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_15_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_14
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_15_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_14
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_15_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_14
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_15_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_14
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_15_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_14
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_15_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_14
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_15_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_14
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_15_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_14
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_15_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_14
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_15_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_14
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_15_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_14
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_15_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_14
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_15_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_14
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_15_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_14 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_14
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_15_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_15 = (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_lpi_1_dfm_mx0)
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_15
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_15
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_15 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_15
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_15
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_15 = ~(nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_lpi_1_dfm_mx0
      | nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_15
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_15
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_15 = nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_lpi_1_dfm_mx0
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_15
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_15
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_15
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_15
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_15
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_15
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_15
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_15
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_15
      & nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_lpi_1_dfm_mx0;
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_15
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_15
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_15
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_15
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_15
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_15
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_15
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_lpi_1_dfm_mx0);
  assign Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_15 = Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_15
      & (~ nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_lpi_1_dfm_mx0);
  assign and_5541_cse = pe_config_is_cluster_sva & (fsm_output[1]);
  assign or_tmp_3038 = state_2_0_sva_0 & (fsm_output[1]);
  assign PECore_RunBias_if_for_or_m1c_5 = (fsm_output[2]) | (fsm_output[4]);
  assign PECore_RunMac_if_or_5_m1c = or_3399_cse | (fsm_output[4]);
  assign PECore_RunMac_if_or_140_m1c = (~ (fsm_output[2])) | or_dcpl_247;
  assign PECore_RunMac_if_and_817_rgt = PECore_RunBias_if_for_and_45_rgt & PECore_RunMac_if_or_140_m1c;
  assign PECore_RunMac_if_and_470_cse = and_dcpl_708 & (fsm_output[2]);
  assign PECore_RunMac_if_and_472_rgt = and_dcpl_706 & (fsm_output[2]);
  assign PECore_RunMac_if_and_444_cse = (~ crossbar_spec_PE_Weight_WordType_16U_16U_for_land_9_lpi_1_dfm)
      & and_dcpl_708 & (fsm_output[2]);
  assign PECore_RunMac_if_and_445_cse = crossbar_spec_PE_Weight_WordType_16U_16U_for_land_9_lpi_1_dfm
      & and_dcpl_708 & (fsm_output[2]);
  assign PECore_RunMac_if_and_398_cse = PECore_RunMac_if_and_12_cse & (fsm_output[2]);
  assign PECore_RunMac_if_and_399_cse = PECore_RunMac_if_and_13_cse & (fsm_output[2]);
  assign PECore_RunMac_if_and_859_cse = PECoreRun_wen & ((~ (fsm_output[2])) | PECore_RunMac_if_and_674_rgt
      | PECore_RunMac_if_and_398_cse | PECore_RunMac_if_and_399_cse);
  assign PECore_RunMac_if_and_390_cse = PECore_RunMac_if_and_10_cse & (fsm_output[2]);
  assign PECore_RunMac_if_and_391_cse = PECore_RunMac_if_and_11_cse & (fsm_output[2]);
  assign PECore_RunMac_if_and_860_cse = PECoreRun_wen & (~ PECore_RunBias_if_for_and_42_cse);
  assign PECore_RunMac_if_and_359_cse = and_dcpl_707 & (~ or_3399_cse);
  assign PECore_RunMac_if_and_360_cse = PECore_RunMac_if_and_10_cse & (~ or_3399_cse);
  assign PECore_RunMac_if_and_361_cse = PECore_RunMac_if_and_11_cse & (~ or_3399_cse);
  assign Datapath_for_and_enex5 = PECore_RunMac_if_and_cse & reg_PECore_RunMac_if_mux_31_enexo;
  assign while_and_74_cse = z_out_12_13 & while_and_46_tmp_1;
  assign while_and_66_cse = z_out_13_13 & while_and_46_tmp_1;
  assign PECore_RunMac_if_and_854_tmp = PECoreRun_wen & (~(PECore_PushAxiRsp_if_asn_66
      & PECore_RunBias_if_for_and_42_cse));
  assign PECore_RunMac_if_and_865_tmp = PECoreRun_wen & (~(PECore_PushAxiRsp_if_asn_66
      & (fsm_output[2]) & PECore_RunMac_if_nand_56_rgt));
  assign operator_16_false_1_mux_10_cse = MUX_v_12_2_2(PEManager_16U_GetWeightAddr_1_else_acc_2_psp_sva_1,
      (PEManager_16U_GetWeightAddr_if_acc_2_psp_sva_1[12:1]), and_5541_cse);
  assign operator_16_false_1_mux_14_cse = MUX_s_1_2_2((PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx1[3]),
      (PEManager_16U_GetWeightAddr_if_acc_2_psp_sva_1[0]), and_5541_cse);
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_input_port_PopNB_mioi_oswt_cse <= 1'b0;
      reg_rva_in_PopNB_mioi_oswt_cse <= 1'b0;
      reg_Datapath_for_1_ProductSum_cmp_cgo_ir_3_cse <= 1'b0;
      reg_input_mem_banks_bank_array_impl_data0_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_array_impl_data15_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_array_impl_data14_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_array_impl_data13_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_array_impl_data12_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_array_impl_data11_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_array_impl_data10_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_array_impl_data9_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_array_impl_data8_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_array_impl_data7_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_array_impl_data6_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_array_impl_data5_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_array_impl_data4_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_array_impl_data3_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_array_impl_data2_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_array_impl_data1_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_array_impl_data0_rsci_cgo_ir_cse <= 1'b0;
      reg_start_PopNB_mioi_iswt0_cse <= 1'b0;
      reg_rva_out_Push_mioi_iswt0_cse <= 1'b0;
      reg_act_port_Push_mioi_iswt0_cse <= 1'b0;
      input_read_req_valid_lpi_1_dfm_5 <= 1'b0;
      weight_mem_write_arbxbar_xbar_for_empty_sva <= 16'b0000000000000000;
      input_write_req_valid_lpi_1_dfm_5 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_lpi_1_dfm <= 1'b0;
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_15_lpi_1_dfm <= 1'b0;
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_14_lpi_1_dfm <= 1'b0;
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_13_lpi_1_dfm <= 1'b0;
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm <= 1'b0;
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_9_lpi_1_dfm <= 1'b0;
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm <= 1'b0;
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm <= 1'b0;
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm <= 1'b0;
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm <= 1'b0;
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm <= 1'b0;
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm <= 1'b0;
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm <= 1'b0;
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_11_lpi_1_dfm <= 1'b0;
      reg_PECore_RunMac_if_mux_1_ftd <= 3'b000;
      reg_PECore_RunMac_if_mux_10_ftd <= 3'b000;
      PECore_RunMac_if_mux_13_itm <= 8'b00000000;
      PECore_RunMac_if_mux_130_itm <= 8'b00000000;
      PECore_RunMac_if_mux_131_itm <= 8'b00000000;
      PECore_RunMac_if_mux_132_itm <= 8'b00000000;
      PECore_RunMac_if_mux_133_itm <= 8'b00000000;
      PECore_RunMac_if_mux_134_itm <= 8'b00000000;
      PECore_RunMac_if_mux_135_itm <= 8'b00000000;
      PECore_RunMac_if_mux_136_itm <= 8'b00000000;
      reg_PECore_RunMac_if_mux_122_ftd <= 4'b0000;
      reg_PECore_RunMac_if_mux_11_ftd <= 4'b0000;
      reg_PECore_RunMac_if_mux_11_ftd_1 <= 4'b0000;
      reg_PECore_RunMac_if_mux_123_ftd <= 4'b0000;
      reg_PECore_RunMac_if_mux_124_ftd <= 4'b0000;
      reg_PECore_RunMac_if_mux_125_ftd <= 4'b0000;
      reg_PECore_RunMac_if_mux_126_ftd <= 4'b0000;
      reg_PECore_RunMac_if_mux_127_ftd <= 4'b0000;
      reg_PECore_RunMac_if_mux_128_ftd <= 4'b0000;
      reg_PECore_RunMac_if_mux_128_ftd_1 <= 4'b0000;
      reg_PECore_RunMac_if_mux_129_ftd <= 4'b0000;
      reg_PECore_RunMac_if_mux_129_ftd_1 <= 4'b0000;
      reg_PECore_RunMac_if_mux_137_ftd <= 6'b000000;
      reg_PECore_RunMac_if_mux_138_ftd <= 3'b000;
      reg_PECore_RunMac_if_mux_139_ftd <= 6'b000000;
      reg_PECore_RunMac_if_mux_14_ftd <= 3'b000;
      reg_PECore_RunMac_if_mux_140_ftd <= 6'b000000;
      reg_PECore_RunMac_if_mux_141_ftd <= 3'b000;
      reg_PECore_RunMac_if_mux_142_ftd <= 4'b0000;
      reg_PECore_RunMac_if_mux_143_ftd <= 1'b0;
    end
    else if ( PECoreRun_wen ) begin
      reg_input_port_PopNB_mioi_oswt_cse <= ~(and_2164_cse | (((~((~(and_5345_cse
          | (pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_pe_config_UpdateInputCounter_if_nor_svs
          & PECore_RunFSM_switch_lp_equal_tmp_1) | (PECore_UpdateFSM_switch_lp_equal_tmp_1
          & PECore_RunMac_nor_tmp) | (~ PECore_RunFSM_switch_lp_equal_tmp) | is_start_sva))
          | state_2_0_sva_2)) | PECore_RunFSM_switch_lp_equal_tmp_2) & (fsm_output[4])));
      reg_rva_in_PopNB_mioi_oswt_cse <= ~(and_2164_cse | (or_1521_cse & (PECore_UpdateFSM_case_4_is_output_end_pe_config_UpdateManagerCounter_nand_itm
          | PECore_UpdateFSM_switch_lp_unequal_tmp | (~ state_2_0_sva_2)) & (fsm_output[4])));
      reg_Datapath_for_1_ProductSum_cmp_cgo_ir_3_cse <= or_2421_rmff;
      reg_input_mem_banks_bank_array_impl_data0_rsci_cgo_ir_cse <= or_2422_rmff;
      reg_weight_mem_banks_bank_array_impl_data15_rsci_cgo_ir_cse <= or_2423_rmff;
      reg_weight_mem_banks_bank_array_impl_data14_rsci_cgo_ir_cse <= or_2424_rmff;
      reg_weight_mem_banks_bank_array_impl_data13_rsci_cgo_ir_cse <= or_2425_rmff;
      reg_weight_mem_banks_bank_array_impl_data12_rsci_cgo_ir_cse <= or_2426_rmff;
      reg_weight_mem_banks_bank_array_impl_data11_rsci_cgo_ir_cse <= or_2427_rmff;
      reg_weight_mem_banks_bank_array_impl_data10_rsci_cgo_ir_cse <= or_2428_rmff;
      reg_weight_mem_banks_bank_array_impl_data9_rsci_cgo_ir_cse <= or_2429_rmff;
      reg_weight_mem_banks_bank_array_impl_data8_rsci_cgo_ir_cse <= or_2430_rmff;
      reg_weight_mem_banks_bank_array_impl_data7_rsci_cgo_ir_cse <= or_2431_rmff;
      reg_weight_mem_banks_bank_array_impl_data6_rsci_cgo_ir_cse <= or_2432_rmff;
      reg_weight_mem_banks_bank_array_impl_data5_rsci_cgo_ir_cse <= or_2433_rmff;
      reg_weight_mem_banks_bank_array_impl_data4_rsci_cgo_ir_cse <= or_2434_rmff;
      reg_weight_mem_banks_bank_array_impl_data3_rsci_cgo_ir_cse <= or_2435_rmff;
      reg_weight_mem_banks_bank_array_impl_data2_rsci_cgo_ir_cse <= or_2436_rmff;
      reg_weight_mem_banks_bank_array_impl_data1_rsci_cgo_ir_cse <= or_2437_rmff;
      reg_weight_mem_banks_bank_array_impl_data0_rsci_cgo_ir_cse <= or_2438_rmff;
      reg_start_PopNB_mioi_iswt0_cse <= and_2966_cse;
      reg_rva_out_Push_mioi_iswt0_cse <= w_axi_rsp_lpi_1_dfm_1 & (~ is_start_sva)
          & (fsm_output[3]);
      reg_act_port_Push_mioi_iswt0_cse <= state_2_0_sva_2 & (~ state_2_0_sva_1) &
          and_dcpl_210 & (fsm_output[3]);
      input_read_req_valid_lpi_1_dfm_5 <= MUX_s_1_2_2(PECore_DecodeAxi_mux_133_nl,
          input_read_req_valid_lpi_1_dfm_6, is_start_sva);
      weight_mem_write_arbxbar_xbar_for_empty_sva <= weight_mem_write_arbxbar_xbar_for_lshift_tmp;
      input_write_req_valid_lpi_1_dfm_5 <= MUX_s_1_2_2(PECore_DecodeAxi_mux_138_nl,
          input_write_req_valid_lpi_1_dfm_6, is_start_sva);
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_lpi_1_dfm <= ~(crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_258_nl
          | (~ weight_read_ack_15_lpi_1_dfm_15_mx0));
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_15_lpi_1_dfm <= ~(crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_257_nl
          | (~ weight_read_ack_14_lpi_1_dfm_15_mx0));
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_14_lpi_1_dfm <= ~(crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_256_nl
          | (~ weight_read_ack_13_lpi_1_dfm_15_mx0));
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_13_lpi_1_dfm <= ~(crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_255_nl
          | (~ weight_read_ack_12_lpi_1_dfm_15_mx0));
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm <= ~(crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_254_nl
          | (~ weight_read_ack_11_lpi_1_dfm_15_mx0));
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_9_lpi_1_dfm <= ~(crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_251_nl
          | (~ weight_read_ack_8_lpi_1_dfm_15_mx0));
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm <= ~(crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_250_nl
          | (~ weight_read_ack_7_lpi_1_dfm_15_mx0));
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm <= ~(crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_249_nl
          | (~ weight_read_ack_6_lpi_1_dfm_15_mx0));
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm <= ~(crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_248_nl
          | (~ weight_read_ack_5_lpi_1_dfm_15_mx0));
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm <= ~(crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_247_nl
          | (~ weight_read_ack_4_lpi_1_dfm_15_mx0));
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm <= ~(crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_246_nl
          | (~ weight_read_ack_3_lpi_1_dfm_15_mx0));
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm <= ~(crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_245_nl
          | (~ weight_read_ack_2_lpi_1_dfm_15_mx0));
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm <= ~(crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_244_nl
          | (~ weight_read_ack_1_lpi_1_dfm_15_mx0));
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_11_lpi_1_dfm <= ~(crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_253_nl
          | (~ weight_read_ack_10_lpi_1_dfm_15_mx0));
      reg_PECore_RunMac_if_mux_1_ftd <= MUX1HOT_v_3_3_2(PEManager_16U_ClusterLookup_for_mux_15_nl,
          (weight_port_read_out_data_0_1_sva_dfm_mx1[7:5]), (crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_12_mx1w2[7:5]),
          {PECore_RunMac_if_and_569_rgt , PECore_RunMac_if_and_570_rgt , PECore_RunBias_if_for_and_42_cse});
      reg_PECore_RunMac_if_mux_10_ftd <= MUX1HOT_v_3_3_2(PEManager_16U_ClusterLookup_for_mux_6_nl,
          (weight_port_read_out_data_0_10_sva_dfm_mx1[7:5]), (crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_11_mx1w2[7:5]),
          {PECore_RunMac_if_and_569_rgt , PECore_RunMac_if_and_570_rgt , PECore_RunBias_if_for_and_42_cse});
      PECore_RunMac_if_mux_13_itm <= MUX1HOT_v_8_3_2(({6'b000000 , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_13_3_2_lpi_1_dfm_1}),
          weight_port_read_out_data_0_13_sva_dfm_mx1, PEManager_16U_ClusterLookup_for_mux_3_nl,
          {(~ (fsm_output[2])) , PECore_RunMac_if_and_433_cse , PECore_RunMac_if_and_434_cse});
      PECore_RunMac_if_mux_130_itm <= MUX1HOT_v_8_4_2(({5'b00000 , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_3_1_lpi_1_dfm_1}),
          weight_port_read_out_data_8_2_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1,
          PEManager_16U_ClusterLookup_for_mux_74_nl, {(~ (fsm_output[2])) , PECore_RunMac_if_and_430_cse
          , PECore_RunMac_if_and_431_cse , PECore_RunMac_if_and_434_cse});
      PECore_RunMac_if_mux_131_itm <= MUX1HOT_v_8_4_2(({6'b000000 , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_5_1_0_lpi_1_dfm_1}),
          weight_port_read_out_data_8_3_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1,
          PEManager_16U_ClusterLookup_for_mux_72_nl, {(~ (fsm_output[2])) , PECore_RunMac_if_and_430_cse
          , PECore_RunMac_if_and_431_cse , PECore_RunMac_if_and_434_cse});
      PECore_RunMac_if_mux_132_itm <= MUX1HOT_v_8_4_2(({6'b000000 , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_5_3_2_lpi_1_dfm_1}),
          weight_port_read_out_data_8_4_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1,
          PEManager_16U_ClusterLookup_for_mux_70_nl, {(~ (fsm_output[2])) , PECore_RunMac_if_and_430_cse
          , PECore_RunMac_if_and_431_cse , PECore_RunMac_if_and_434_cse});
      PECore_RunMac_if_mux_133_itm <= MUX1HOT_v_8_4_2(({5'b00000 , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_3_1_lpi_1_dfm_1}),
          weight_port_read_out_data_8_5_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1,
          PEManager_16U_ClusterLookup_for_mux_68_nl, {(~ (fsm_output[2])) , PECore_RunMac_if_and_430_cse
          , PECore_RunMac_if_and_431_cse , PECore_RunMac_if_and_434_cse});
      PECore_RunMac_if_mux_134_itm <= MUX1HOT_v_8_4_2(({4'b0000 , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_8_lpi_1_dfm_1}),
          weight_port_read_out_data_8_6_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1,
          PEManager_16U_ClusterLookup_for_mux_66_nl, {(~ (fsm_output[2])) , PECore_RunMac_if_and_430_cse
          , PECore_RunMac_if_and_431_cse , PECore_RunMac_if_and_434_cse});
      PECore_RunMac_if_mux_135_itm <= MUX1HOT_v_8_4_2(({5'b00000 , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_2_0_lpi_1_dfm_1}),
          weight_port_read_out_data_8_7_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1,
          PEManager_16U_ClusterLookup_for_mux_64_nl, {(~ (fsm_output[2])) , PECore_RunMac_if_and_430_cse
          , PECore_RunMac_if_and_431_cse , PECore_RunMac_if_and_434_cse});
      PECore_RunMac_if_mux_136_itm <= MUX1HOT_v_8_4_2(({4'b0000 , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_lpi_1_dfm_1}),
          weight_port_read_out_data_8_8_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1,
          PEManager_16U_ClusterLookup_for_mux_65_nl, {(~ (fsm_output[2])) , PECore_RunMac_if_and_430_cse
          , PECore_RunMac_if_and_431_cse , PECore_RunMac_if_and_434_cse});
      reg_PECore_RunMac_if_mux_122_ftd <= MUX_v_4_2_2(PEManager_16U_ClusterLookup_1_for_mux_53_nl,
          (weight_port_read_out_data_7_10_sva_dfm_mx1[7:4]), PECore_RunMac_if_and_570_rgt);
      reg_PECore_RunMac_if_mux_11_ftd <= MUX1HOT_v_4_3_2(PEManager_16U_ClusterLookup_for_mux_5_nl,
          (weight_port_read_out_data_0_11_sva_dfm_mx1[7:4]), (crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_13_mx1w2[7:4]),
          {PECore_RunMac_if_and_569_rgt , PECore_RunMac_if_and_570_rgt , PECore_RunBias_if_for_and_42_cse});
      reg_PECore_RunMac_if_mux_11_ftd_1 <= MUX1HOT_v_4_5_2(crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_10_lpi_1_dfm_1,
          adpfloat_tmp_to_fixed_20U_14U_acc_sdt_12_sva_mx0w1, PEManager_16U_ClusterLookup_for_mux_138_nl,
          (weight_port_read_out_data_0_11_sva_dfm_mx1[3:0]), (crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_13_mx1w2[3:0]),
          {(~ (fsm_output[2])) , PECore_RunMac_if_and_820_rgt , PECore_RunMac_if_and_569_rgt
          , PECore_RunMac_if_and_570_rgt , PECore_RunBias_if_for_and_42_cse});
      reg_PECore_RunMac_if_mux_123_ftd <= MUX_v_4_2_2(PEManager_16U_ClusterLookup_1_for_mux_55_nl,
          (weight_port_read_out_data_7_11_sva_dfm_mx1[7:4]), PECore_RunMac_if_and_570_rgt);
      reg_PECore_RunMac_if_mux_124_ftd <= MUX_v_4_2_2(PEManager_16U_ClusterLookup_1_for_mux_57_nl,
          (weight_port_read_out_data_7_12_sva_dfm_mx1[7:4]), PECore_RunMac_if_and_470_cse);
      reg_PECore_RunMac_if_mux_125_ftd <= MUX_v_4_2_2(PEManager_16U_ClusterLookup_1_for_mux_59_nl,
          (weight_port_read_out_data_7_13_sva_dfm_mx1[7:4]), PECore_RunMac_if_and_470_cse);
      reg_PECore_RunMac_if_mux_126_ftd <= MUX_v_4_2_2(PEManager_16U_ClusterLookup_1_for_mux_61_nl,
          (weight_port_read_out_data_7_14_sva_dfm_mx1[7:4]), PECore_RunMac_if_and_470_cse);
      reg_PECore_RunMac_if_mux_127_ftd <= MUX_v_4_2_2(PEManager_16U_ClusterLookup_1_for_mux_63_nl,
          (weight_port_read_out_data_7_15_sva_dfm_mx1[7:4]), PECore_RunMac_if_and_470_cse);
      reg_PECore_RunMac_if_mux_128_ftd <= MUX1HOT_v_4_3_2(PEManager_16U_ClusterLookup_for_mux_78_nl,
          (weight_port_read_out_data_8_0_sva_dfm[7:4]), (crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1[7:4]),
          {PECore_RunMac_if_and_472_rgt , PECore_RunMac_if_and_444_cse , PECore_RunMac_if_and_445_cse});
      reg_PECore_RunMac_if_mux_128_ftd_1 <= MUX1HOT_v_4_5_2(crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_4_lpi_1_dfm_1,
          adpfloat_tmp_to_fixed_20U_14U_acc_sdt_8_sva_mx0w1, PEManager_16U_ClusterLookup_for_mux_137_nl,
          (weight_port_read_out_data_8_0_sva_dfm[3:0]), (crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1[3:0]),
          {(~ (fsm_output[2])) , PECore_RunMac_if_and_571_rgt , PECore_RunMac_if_and_472_rgt
          , PECore_RunMac_if_and_444_cse , PECore_RunMac_if_and_445_cse});
      reg_PECore_RunMac_if_mux_129_ftd <= MUX1HOT_v_4_3_2(PEManager_16U_ClusterLookup_for_mux_76_nl,
          (weight_port_read_out_data_8_1_sva_dfm[7:4]), (crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1[7:4]),
          {PECore_RunMac_if_and_472_rgt , PECore_RunMac_if_and_444_cse , PECore_RunMac_if_and_445_cse});
      reg_PECore_RunMac_if_mux_129_ftd_1 <= MUX1HOT_v_4_5_2(crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_6_lpi_1_dfm_1,
          adpfloat_tmp_to_fixed_20U_14U_acc_sdt_9_sva_mx0w1, PEManager_16U_ClusterLookup_for_mux_136_nl,
          (weight_port_read_out_data_8_1_sva_dfm[3:0]), (crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1[3:0]),
          {(~ (fsm_output[2])) , PECore_RunMac_if_and_571_rgt , PECore_RunMac_if_and_472_rgt
          , PECore_RunMac_if_and_444_cse , PECore_RunMac_if_and_445_cse});
      reg_PECore_RunMac_if_mux_137_ftd <= MUX1HOT_v_6_3_2(PEManager_16U_ClusterLookup_for_mux_67_nl,
          (weight_port_read_out_data_8_9_sva_dfm[7:2]), (crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1[7:2]),
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_398_cse , PECore_RunMac_if_and_399_cse});
      reg_PECore_RunMac_if_mux_138_ftd <= MUX1HOT_v_3_3_2(PEManager_16U_ClusterLookup_for_mux_69_nl,
          (weight_port_read_out_data_8_10_sva_dfm[7:5]), (crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1[7:5]),
          {PECore_RunMac_if_and_569_rgt , PECore_RunMac_if_and_390_cse , PECore_RunMac_if_and_391_cse});
      reg_PECore_RunMac_if_mux_139_ftd <= MUX1HOT_v_6_3_2(PEManager_16U_ClusterLookup_for_mux_71_nl,
          (weight_port_read_out_data_8_11_sva_dfm[7:2]), (crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1[7:2]),
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_398_cse , PECore_RunMac_if_and_399_cse});
      reg_PECore_RunMac_if_mux_14_ftd <= MUX_v_3_2_2(PEManager_16U_ClusterLookup_for_mux_2_nl,
          (weight_port_read_out_data_0_14_sva_dfm_mx1[7:5]), PECore_RunMac_if_and_570_rgt);
      reg_PECore_RunMac_if_mux_140_ftd <= MUX1HOT_v_6_3_2(PEManager_16U_ClusterLookup_for_mux_73_nl,
          (weight_port_read_out_data_8_12_sva_dfm[7:2]), (crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1[7:2]),
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_398_cse , PECore_RunMac_if_and_399_cse});
      reg_PECore_RunMac_if_mux_141_ftd <= MUX1HOT_v_3_3_2(PEManager_16U_ClusterLookup_for_mux_75_nl,
          (weight_port_read_out_data_8_13_sva_dfm[7:5]), (crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1[7:5]),
          {PECore_RunMac_if_and_359_cse , PECore_RunMac_if_and_360_cse , PECore_RunMac_if_and_361_cse});
      reg_PECore_RunMac_if_mux_142_ftd <= MUX1HOT_v_4_3_2(PEManager_16U_ClusterLookup_for_mux_77_nl,
          (weight_port_read_out_data_8_14_sva_dfm[7:4]), (crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1[7:4]),
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_398_cse , PECore_RunMac_if_and_399_cse});
      reg_PECore_RunMac_if_mux_143_ftd <= MUX1HOT_s_1_3_2(PEManager_16U_ClusterLookup_for_mux_79_nl,
          (weight_port_read_out_data_8_15_sva_dfm[7]), (crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1[7]),
          {and_dcpl_704 , PECore_RunMac_if_and_12_cse , PECore_RunMac_if_and_13_cse});
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_idat_0 <= 1'b0;
      rva_out_Push_mioi_idat_8 <= 1'b0;
      rva_out_Push_mioi_idat_16 <= 1'b0;
      rva_out_Push_mioi_idat_24 <= 1'b0;
    end
    else if ( PECore_PushAxiRsp_if_and_cse ) begin
      rva_out_Push_mioi_idat_0 <= MUX_s_1_2_2((weight_port_read_out_data_0_0_sva_dfm[0]),
          PECore_PushAxiRsp_if_else_mux_14_nl, or_tmp_1655);
      rva_out_Push_mioi_idat_8 <= MUX_s_1_2_2((reg_PECore_RunMac_if_mux_11_ftd_1[0]),
          PECore_PushAxiRsp_if_else_mux_15_nl, or_tmp_1655);
      rva_out_Push_mioi_idat_16 <= MUX_s_1_2_2((reg_PECore_RunMac_if_mux_1_ftd_1[0]),
          PECore_PushAxiRsp_if_else_mux_16_nl, or_tmp_1655);
      rva_out_Push_mioi_idat_24 <= MUX_s_1_2_2((reg_PECore_RunMac_if_mux_10_ftd_1[0]),
          PECore_PushAxiRsp_if_else_mux_17_nl, or_tmp_1655);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_idat_7_1 <= 7'b0000000;
      rva_out_Push_mioi_idat_10_9 <= 2'b00;
      rva_out_Push_mioi_idat_15_11 <= 5'b00000;
      rva_out_Push_mioi_idat_18_17 <= 2'b00;
      rva_out_Push_mioi_idat_23_19 <= 5'b00000;
      rva_out_Push_mioi_idat_26_25 <= 2'b00;
      rva_out_Push_mioi_idat_31_27 <= 5'b00000;
    end
    else if ( PECore_PushAxiRsp_if_and_10_cse ) begin
      rva_out_Push_mioi_idat_7_1 <= MUX1HOT_v_7_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_18_nl,
          (input_mem_banks_read_read_data_lpi_1[7:1]), (weight_port_read_out_data_0_0_sva_dfm[7:1]),
          reg_PECore_RunMac_if_mux_143_ftd_1, {and_5501_cse , and_5502_cse , crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm
          , or_dcpl_717});
      rva_out_Push_mioi_idat_10_9 <= MUX1HOT_v_2_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl,
          (input_mem_banks_read_read_data_lpi_1[10:9]), (reg_PECore_RunMac_if_mux_11_ftd_1[2:1]),
          reg_PECore_RunMac_if_mux_137_ftd_1, {and_5501_cse , and_5502_cse , crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm
          , or_dcpl_717});
      rva_out_Push_mioi_idat_15_11 <= MUX1HOT_v_5_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_15_nl,
          (input_mem_banks_read_read_data_lpi_1[15:11]), ({reg_PECore_RunMac_if_mux_11_ftd
          , (reg_PECore_RunMac_if_mux_11_ftd_1[3])}), reg_PECore_RunMac_if_mux_138_ftd_1,
          {and_5501_cse , and_5502_cse , crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm
          , or_dcpl_717});
      rva_out_Push_mioi_idat_18_17 <= MUX1HOT_v_2_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_12_nl,
          (input_mem_banks_read_read_data_lpi_1[18:17]), (reg_PECore_RunMac_if_mux_1_ftd_1[2:1]),
          reg_PECore_RunMac_if_mux_139_ftd_1, {and_5501_cse , and_5502_cse , crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm
          , or_dcpl_717});
      rva_out_Push_mioi_idat_23_19 <= MUX1HOT_v_5_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_10_nl,
          (input_mem_banks_read_read_data_lpi_1[23:19]), ({reg_PECore_RunMac_if_mux_1_ftd
          , (reg_PECore_RunMac_if_mux_1_ftd_1[4:3])}), reg_PECore_RunMac_if_mux_14_ftd_1,
          {and_5501_cse , and_5502_cse , crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm
          , or_dcpl_717});
      rva_out_Push_mioi_idat_26_25 <= MUX1HOT_v_2_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_9_nl,
          (input_mem_banks_read_read_data_lpi_1[26:25]), (reg_PECore_RunMac_if_mux_10_ftd_1[2:1]),
          reg_PECore_RunMac_if_mux_140_ftd_1, {and_5501_cse , and_5502_cse , crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm
          , or_dcpl_717});
      rva_out_Push_mioi_idat_31_27 <= MUX1HOT_v_5_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl,
          (input_mem_banks_read_read_data_lpi_1[31:27]), ({reg_PECore_RunMac_if_mux_10_ftd
          , (reg_PECore_RunMac_if_mux_10_ftd_1[4:3])}), reg_PECore_RunMac_if_mux_141_ftd_1,
          {and_5501_cse , and_5502_cse , crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm
          , or_dcpl_717});
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_idat_35_32 <= 4'b0000;
    end
    else if ( PECore_PushAxiRsp_if_and_47_enex5 ) begin
      rva_out_Push_mioi_idat_35_32 <= reg_PECore_RunMac_if_mux_123_ftd_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_idat_39_36 <= 4'b0000;
    end
    else if ( PECore_PushAxiRsp_if_and_48_enex5 ) begin
      rva_out_Push_mioi_idat_39_36 <= reg_PECore_RunMac_if_mux_142_ftd_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_idat_47_40 <= 8'b00000000;
    end
    else if ( PECore_PushAxiRsp_if_and_49_enex5 ) begin
      rva_out_Push_mioi_idat_47_40 <= rva_out_reg_data_47_40_sva_dfm_4;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_idat_55_48 <= 8'b00000000;
    end
    else if ( PECore_PushAxiRsp_if_and_50_enex5 ) begin
      rva_out_Push_mioi_idat_55_48 <= rva_out_reg_data_55_48_sva_dfm_4;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_idat_63_56 <= 8'b00000000;
    end
    else if ( PECore_PushAxiRsp_if_and_51_enex5 ) begin
      rva_out_Push_mioi_idat_63_56 <= rva_out_reg_data_63_56_sva_dfm_4;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_idat_71_64 <= 8'b00000000;
    end
    else if ( PECore_PushAxiRsp_if_and_52_enex5 ) begin
      rva_out_Push_mioi_idat_71_64 <= rva_out_reg_data_71_64_sva_dfm_4;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_idat_79_72 <= 8'b00000000;
    end
    else if ( PECore_PushAxiRsp_if_and_53_enex5 ) begin
      rva_out_Push_mioi_idat_79_72 <= rva_out_reg_data_79_72_sva_dfm_4;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_idat_87_80 <= 8'b00000000;
    end
    else if ( PECore_PushAxiRsp_if_and_54_enex5 ) begin
      rva_out_Push_mioi_idat_87_80 <= rva_out_reg_data_87_80_sva_dfm_4;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_idat_95_88 <= 8'b00000000;
    end
    else if ( PECore_PushAxiRsp_if_and_55_enex5 ) begin
      rva_out_Push_mioi_idat_95_88 <= rva_out_reg_data_95_88_sva_dfm_4;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_idat_103_96 <= 8'b00000000;
    end
    else if ( PECore_PushAxiRsp_if_and_56_enex5 ) begin
      rva_out_Push_mioi_idat_103_96 <= rva_out_reg_data_103_96_sva_dfm_4;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_idat_111_104 <= 8'b00000000;
    end
    else if ( PECore_PushAxiRsp_if_and_57_enex5 ) begin
      rva_out_Push_mioi_idat_111_104 <= rva_out_reg_data_111_104_sva_dfm_4;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_idat_119_112 <= 8'b00000000;
    end
    else if ( PECore_PushAxiRsp_if_and_58_enex5 ) begin
      rva_out_Push_mioi_idat_119_112 <= rva_out_reg_data_119_112_sva_dfm_4;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_idat_127_120 <= 8'b00000000;
    end
    else if ( PECore_PushAxiRsp_if_and_59_enex5 ) begin
      rva_out_Push_mioi_idat_127_120 <= rva_out_reg_data_127_120_sva_dfm_4;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_Push_mioi_idat_19_0 <= 20'b00000000000000000000;
      act_port_Push_mioi_idat_159_140 <= 20'b00000000000000000000;
      act_port_Push_mioi_idat_179_160 <= 20'b00000000000000000000;
      act_port_Push_mioi_idat_239_220 <= 20'b00000000000000000000;
    end
    else if ( PECore_PushOutput_if_and_16_enex5 ) begin
      act_port_Push_mioi_idat_19_0 <= act_port_reg_data_0_sva;
      act_port_Push_mioi_idat_159_140 <= act_port_reg_data_7_sva;
      act_port_Push_mioi_idat_179_160 <= act_port_reg_data_8_sva;
      act_port_Push_mioi_idat_239_220 <= act_port_reg_data_11_sva;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_Push_mioi_idat_39_20 <= 20'b00000000000000000000;
    end
    else if ( PECore_PushOutput_if_and_17_enex5 ) begin
      act_port_Push_mioi_idat_39_20 <= act_port_reg_data_1_sva;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_Push_mioi_idat_59_40 <= 20'b00000000000000000000;
    end
    else if ( PECore_PushOutput_if_and_18_enex5 ) begin
      act_port_Push_mioi_idat_59_40 <= act_port_reg_data_2_sva;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_Push_mioi_idat_79_60 <= 20'b00000000000000000000;
    end
    else if ( PECore_PushOutput_if_and_19_enex5 ) begin
      act_port_Push_mioi_idat_79_60 <= act_port_reg_data_3_sva;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_Push_mioi_idat_99_80 <= 20'b00000000000000000000;
    end
    else if ( PECore_PushOutput_if_and_20_enex5 ) begin
      act_port_Push_mioi_idat_99_80 <= act_port_reg_data_4_sva;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_Push_mioi_idat_119_100 <= 20'b00000000000000000000;
    end
    else if ( PECore_PushOutput_if_and_21_enex5 ) begin
      act_port_Push_mioi_idat_119_100 <= act_port_reg_data_5_sva;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_Push_mioi_idat_139_120 <= 20'b00000000000000000000;
    end
    else if ( PECore_PushOutput_if_and_22_enex5 ) begin
      act_port_Push_mioi_idat_139_120 <= act_port_reg_data_6_sva;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_Push_mioi_idat_199_180 <= 20'b00000000000000000000;
    end
    else if ( PECore_PushOutput_if_and_25_enex5 ) begin
      act_port_Push_mioi_idat_199_180 <= act_port_reg_data_9_sva;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_Push_mioi_idat_219_200 <= 20'b00000000000000000000;
    end
    else if ( PECore_PushOutput_if_and_26_enex5 ) begin
      act_port_Push_mioi_idat_219_200 <= act_port_reg_data_10_sva;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_Push_mioi_idat_259_240 <= 20'b00000000000000000000;
    end
    else if ( PECore_PushOutput_if_and_28_enex5 ) begin
      act_port_Push_mioi_idat_259_240 <= act_port_reg_data_asn_3_itm;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_Push_mioi_idat_279_260 <= 20'b00000000000000000000;
    end
    else if ( PECore_PushOutput_if_and_29_enex5 ) begin
      act_port_Push_mioi_idat_279_260 <= act_port_reg_data_asn_2_itm;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_Push_mioi_idat_299_280 <= 20'b00000000000000000000;
    end
    else if ( PECore_PushOutput_if_and_30_enex5 ) begin
      act_port_Push_mioi_idat_299_280 <= act_port_reg_data_asn_1_itm;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_Push_mioi_idat_319_300 <= 20'b00000000000000000000;
    end
    else if ( PECore_PushOutput_if_and_31_enex5 ) begin
      act_port_Push_mioi_idat_319_300 <= act_port_reg_data_asn_itm;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      is_start_sva <= 1'b0;
      state_2_0_sva_2 <= 1'b0;
      state_2_0_sva_1 <= 1'b0;
      state_2_0_sva_0 <= 1'b0;
      accum_vector_data_8_sva <= 32'b00000000000000000000000000000000;
      accum_vector_data_7_sva <= 32'b00000000000000000000000000000000;
      act_port_reg_data_1_sva <= 20'b00000000000000000000;
      act_port_reg_data_2_sva <= 20'b00000000000000000000;
      act_port_reg_data_3_sva <= 20'b00000000000000000000;
      act_port_reg_data_4_sva <= 20'b00000000000000000000;
      reg_PECore_RunMac_asn_15_itm_1_ftd <= 1'b0;
      reg_PECore_RunMac_asn_15_itm_1_ftd_1 <= 1'b0;
      reg_PECore_RunMac_asn_15_itm_1_ftd_2 <= 1'b0;
      while_asn_41_itm_1 <= 1'b0;
      while_stage_0_2 <= 1'b0;
      while_and_29_itm_1 <= 1'b0;
      PECore_RunBias_if_accum_vector_out_data_13_lpi_1_dfm <= 32'b00000000000000000000000000000000;
      PECore_RunBias_if_accum_vector_out_data_lpi_1_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( is_start_and_cse ) begin
      is_start_sva <= MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_mux_6_nl, or_1521_cse,
          and_3383_nl);
      state_2_0_sva_2 <= PECore_RunFSM_switch_lp_equal_tmp_2;
      state_2_0_sva_1 <= ~(PECore_RunFSM_switch_lp_equal_tmp | PECore_RunFSM_switch_lp_equal_tmp_2
          | state_2_0_sva_2);
      state_2_0_sva_0 <= ~((~(PECore_UpdateFSM_switch_lp_mux1h_42_nl & (~ PECore_RunFSM_switch_lp_equal_tmp_2)))
          | state_2_0_sva_2);
      accum_vector_data_8_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_15_cse;
      accum_vector_data_7_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_14_cse;
      act_port_reg_data_1_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_25_cse;
      act_port_reg_data_2_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_26_cse;
      act_port_reg_data_3_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_21_cse;
      act_port_reg_data_4_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_22_cse;
      reg_PECore_RunMac_asn_15_itm_1_ftd <= state_2_0_sva_2;
      reg_PECore_RunMac_asn_15_itm_1_ftd_1 <= state_2_0_sva_1;
      reg_PECore_RunMac_asn_15_itm_1_ftd_2 <= state_2_0_sva_0;
      while_asn_41_itm_1 <= is_start_sva;
      while_stage_0_2 <= 1'b1;
      while_and_29_itm_1 <= while_and_30_itm_1;
      PECore_RunBias_if_accum_vector_out_data_13_lpi_1_dfm <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_12_cse;
      PECore_RunBias_if_accum_vector_out_data_lpi_1_dfm <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_13_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      accum_vector_data_4_sva <= 32'b00000000000000000000000000000000;
      accum_vector_data_3_sva <= 32'b00000000000000000000000000000000;
      accum_vector_data_2_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( accum_vector_data_and_6_cse ) begin
      accum_vector_data_4_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_4_cse;
      accum_vector_data_3_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_3_cse;
      accum_vector_data_2_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_2_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_reg_data_10_sva <= 20'b00000000000000000000;
      act_port_reg_data_9_sva <= 20'b00000000000000000000;
      act_port_reg_data_6_sva <= 20'b00000000000000000000;
      act_port_reg_data_5_sva <= 20'b00000000000000000000;
    end
    else if ( act_port_reg_data_and_8_cse ) begin
      act_port_reg_data_10_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_26_cse;
      act_port_reg_data_9_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_25_cse;
      act_port_reg_data_6_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_22_cse;
      act_port_reg_data_5_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_21_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_lpi_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & input_read_req_valid_lpi_1_dfm_5 & (~ input_write_req_valid_lpi_1_dfm_5)
        & (fsm_output[2]) ) begin
      input_mem_banks_read_read_data_lpi_1 <= input_mem_banks_bank_array_impl_data0_rsci_q_d;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      while_and_46_tmp_1 <= 1'b0;
      pe_manager_cluster_lut_data_1_0_sva_0 <= 1'b0;
      pe_manager_cluster_lut_data_1_1_sva_0 <= 1'b0;
      pe_manager_cluster_lut_data_1_2_sva_0 <= 1'b0;
      pe_manager_cluster_lut_data_1_3_sva_0 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm <= 1'b0;
      crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm <= 1'b0;
      crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm <= 1'b0;
      crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm <= 1'b0;
    end
    else if ( while_and_cse ) begin
      while_and_46_tmp_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_16U_16U_for_if_1_crossbar_spec_PE_Weight_WordType_16U_16U_for_if_1_crossbar_spec_PE_Weight_WordType_16U_16U_for_if_1_nor_5_nl,
          while_and_48_tmp_1, fsm_output[2]);
      pe_manager_cluster_lut_data_1_0_sva_0 <= pe_manager_cluster_lut_data_1_0_sva_dfm_4[0];
      pe_manager_cluster_lut_data_1_1_sva_0 <= pe_manager_cluster_lut_data_1_1_sva_dfm_4[0];
      pe_manager_cluster_lut_data_1_2_sva_0 <= pe_manager_cluster_lut_data_1_2_sva_dfm_4[0];
      pe_manager_cluster_lut_data_1_3_sva_0 <= pe_manager_cluster_lut_data_1_3_sva_dfm_4[0];
      crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm_1,
          (pe_manager_cluster_lut_data_0_0_sva_dfm_4[0]), fsm_output[2]);
      crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm_1,
          (pe_manager_cluster_lut_data_0_1_sva_dfm_4[0]), fsm_output[2]);
      crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm_1,
          (pe_manager_cluster_lut_data_0_2_sva_dfm_4[0]), fsm_output[2]);
      crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm_1,
          (pe_manager_cluster_lut_data_0_3_sva_dfm_4[0]), fsm_output[2]);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      pe_manager_adplfloat_bias_weight_0_sva <= 3'b000;
      pe_manager_adplfloat_bias_bias_0_sva <= 3'b000;
      pe_manager_adplfloat_bias_input_0_sva <= 3'b000;
      pe_manager_base_input_0_sva <= 16'b0000000000000000;
      pe_manager_num_input_0_sva <= 8'b00000001;
      pe_manager_base_bias_0_sva <= 16'b0000000000000000;
      pe_manager_base_weight_0_sva <= 16'b0000000000000000;
    end
    else if ( pe_manager_adplfloat_bias_weight_and_cse ) begin
      pe_manager_adplfloat_bias_weight_0_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[10:8];
      pe_manager_adplfloat_bias_bias_0_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[18:16];
      pe_manager_adplfloat_bias_input_0_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[26:24];
      pe_manager_base_input_0_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[95:80];
      pe_manager_num_input_0_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[39:32];
      pe_manager_base_bias_0_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[79:64];
      pe_manager_base_weight_0_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[63:48];
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      pe_manager_adplfloat_bias_weight_1_sva <= 3'b000;
      pe_manager_adplfloat_bias_bias_1_sva <= 3'b000;
      pe_manager_adplfloat_bias_input_1_sva <= 3'b000;
      pe_manager_base_input_1_sva <= 16'b0000000000000000;
      pe_manager_num_input_1_sva <= 8'b00000001;
      pe_manager_base_bias_1_sva <= 16'b0000000000000000;
      pe_manager_base_weight_1_sva <= 16'b0000000000000000;
    end
    else if ( pe_manager_adplfloat_bias_weight_and_1_cse ) begin
      pe_manager_adplfloat_bias_weight_1_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[10:8];
      pe_manager_adplfloat_bias_bias_1_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[18:16];
      pe_manager_adplfloat_bias_input_1_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[26:24];
      pe_manager_base_input_1_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[95:80];
      pe_manager_num_input_1_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[39:32];
      pe_manager_base_bias_1_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[79:64];
      pe_manager_base_weight_1_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[63:48];
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      pe_manager_cluster_lut_data_0_4_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_0_5_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_0_12_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_0_13_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_0_14_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_0_15_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_0_10_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_0_11_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_0_8_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_0_9_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_0_6_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_0_7_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_0_0_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_0_1_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_0_2_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_0_3_sva_dfm_4 <= 8'b00000000;
    end
    else if ( pe_manager_cluster_lut_data_and_cse ) begin
      pe_manager_cluster_lut_data_0_4_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[39:32];
      pe_manager_cluster_lut_data_0_5_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[47:40];
      pe_manager_cluster_lut_data_0_12_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[103:96];
      pe_manager_cluster_lut_data_0_13_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[111:104];
      pe_manager_cluster_lut_data_0_14_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[119:112];
      pe_manager_cluster_lut_data_0_15_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[127:120];
      pe_manager_cluster_lut_data_0_10_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[87:80];
      pe_manager_cluster_lut_data_0_11_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[95:88];
      pe_manager_cluster_lut_data_0_8_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[71:64];
      pe_manager_cluster_lut_data_0_9_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[79:72];
      pe_manager_cluster_lut_data_0_6_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[55:48];
      pe_manager_cluster_lut_data_0_7_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[63:56];
      pe_manager_cluster_lut_data_0_0_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[7:0];
      pe_manager_cluster_lut_data_0_1_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[15:8];
      pe_manager_cluster_lut_data_0_2_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[23:16];
      pe_manager_cluster_lut_data_0_3_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[31:24];
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      pe_manager_cluster_lut_data_1_4_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_1_5_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_1_12_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_1_13_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_1_14_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_1_15_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_1_10_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_1_11_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_1_8_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_1_9_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_1_6_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_1_7_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_1_0_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_1_1_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_1_2_sva_dfm_4 <= 8'b00000000;
      pe_manager_cluster_lut_data_1_3_sva_dfm_4 <= 8'b00000000;
    end
    else if ( pe_manager_cluster_lut_data_and_1_cse ) begin
      pe_manager_cluster_lut_data_1_4_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[39:32];
      pe_manager_cluster_lut_data_1_5_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[47:40];
      pe_manager_cluster_lut_data_1_12_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[103:96];
      pe_manager_cluster_lut_data_1_13_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[111:104];
      pe_manager_cluster_lut_data_1_14_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[119:112];
      pe_manager_cluster_lut_data_1_15_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[127:120];
      pe_manager_cluster_lut_data_1_10_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[87:80];
      pe_manager_cluster_lut_data_1_11_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[95:88];
      pe_manager_cluster_lut_data_1_8_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[71:64];
      pe_manager_cluster_lut_data_1_9_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[79:72];
      pe_manager_cluster_lut_data_1_6_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[55:48];
      pe_manager_cluster_lut_data_1_7_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[63:56];
      pe_manager_cluster_lut_data_1_0_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[7:0];
      pe_manager_cluster_lut_data_1_1_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[15:8];
      pe_manager_cluster_lut_data_1_2_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[23:16];
      pe_manager_cluster_lut_data_1_3_sva_dfm_4 <= rva_in_PopNB_mio_mrgout_dat_sva_1[31:24];
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      pe_config_manager_counter_sva <= 4'b0000;
    end
    else if ( (((~((rva_in_PopNB_mioi_idat_mxwt[137:135]!=3'b000))) & (~((rva_in_PopNB_mioi_idat_mxwt[140:138]!=3'b000)))
        & (~((rva_in_PopNB_mioi_idat_mxwt[143:141]!=3'b000))) & (~((rva_in_PopNB_mioi_idat_mxwt[146:144]!=3'b000)))
        & (~((rva_in_PopNB_mioi_idat_mxwt[147]) | (rva_in_PopNB_mioi_idat_mxwt[134])
        | (rva_in_PopNB_mioi_idat_mxwt[133]))) & (rva_in_PopNB_mioi_idat_mxwt[132])
        & (rva_in_PopNB_mioi_idat_mxwt[168]) & (~ (rva_in_PopNB_mioi_idat_mxwt[148]))
        & (~(is_start_sva | (rva_in_PopNB_mioi_idat_mxwt[149]) | (rva_in_PopNB_mioi_idat_mxwt[151])))
        & rva_in_PopNB_mioi_ivld_mxwt & (rva_in_PopNB_mioi_idat_mxwt[150])) | and_5844_cse)
        & (fsm_output[1]) & PECoreRun_wen ) begin
      pe_config_manager_counter_sva <= MUX_v_4_2_2(pe_config_manager_counter_sva_dfm_4_mx1,
          pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_and_1_nl,
          and_3501_nl);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_15_15_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_15_0_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_15_14_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_15_1_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_15_13_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_15_2_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_15_12_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_15_3_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_15_11_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_15_4_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_15_10_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_15_5_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_15_9_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_15_6_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_15_8_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_15_7_sva_dfm <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_cse ) begin
      weight_port_read_out_data_15_15_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_15_0_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_1_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_15_14_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_15_1_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_2_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_15_13_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_15_2_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_3_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_15_12_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_13_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_15_3_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_4_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_15_11_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_12_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_15_4_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_5_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_15_10_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_11_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_15_5_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_6_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_15_9_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_10_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_15_6_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_7_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_15_8_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_9_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_15_7_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_8_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_14_15_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_14_0_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_14_14_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_14_1_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_14_13_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_14_2_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_14_12_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_14_3_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_14_11_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_14_4_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_14_10_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_14_5_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_14_9_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_14_6_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_14_8_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_14_7_sva_dfm <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_16_cse ) begin
      weight_port_read_out_data_14_15_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_14_0_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_1_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_14_14_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_14_1_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_2_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_14_13_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_14_2_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_3_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_14_12_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_13_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_14_3_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_4_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_14_11_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_12_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_14_4_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_5_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_14_10_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_11_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_14_5_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_6_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_14_9_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_10_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_14_6_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_7_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_14_8_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_9_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_14_7_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_8_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_13_15_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_13_0_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_13_14_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_13_1_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_13_13_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_13_2_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_13_12_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_13_3_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_13_11_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_13_4_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_13_10_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_13_5_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_13_9_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_13_6_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_13_8_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_13_7_sva_dfm <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_32_cse ) begin
      weight_port_read_out_data_13_15_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_13_0_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_41;
      weight_port_read_out_data_13_14_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_13_1_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_39;
      weight_port_read_out_data_13_13_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_15;
      weight_port_read_out_data_13_2_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_37;
      weight_port_read_out_data_13_12_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_17;
      weight_port_read_out_data_13_3_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_35;
      weight_port_read_out_data_13_11_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_19;
      weight_port_read_out_data_13_4_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_33;
      weight_port_read_out_data_13_10_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_21;
      weight_port_read_out_data_13_5_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_31;
      weight_port_read_out_data_13_9_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_23;
      weight_port_read_out_data_13_6_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_29;
      weight_port_read_out_data_13_8_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_25;
      weight_port_read_out_data_13_7_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_27;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_12_15_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_12_0_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_12_14_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_12_1_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_12_13_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_12_2_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_12_12_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_12_3_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_12_11_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_12_4_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_12_10_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_12_5_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_12_9_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_12_6_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_12_8_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_12_7_sva_dfm <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_48_cse ) begin
      weight_port_read_out_data_12_15_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1;
      weight_port_read_out_data_12_0_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1;
      weight_port_read_out_data_12_14_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1;
      weight_port_read_out_data_12_1_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1;
      weight_port_read_out_data_12_13_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1;
      weight_port_read_out_data_12_2_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1;
      weight_port_read_out_data_12_12_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1;
      weight_port_read_out_data_12_3_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1;
      weight_port_read_out_data_12_11_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1;
      weight_port_read_out_data_12_4_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1;
      weight_port_read_out_data_12_10_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1;
      weight_port_read_out_data_12_5_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1;
      weight_port_read_out_data_12_9_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1;
      weight_port_read_out_data_12_6_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1;
      weight_port_read_out_data_12_8_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1;
      weight_port_read_out_data_12_7_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_11_0_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_11_1_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_11_2_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_11_3_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_11_4_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_11_5_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_11_6_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_11_7_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_11_8_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_11_9_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_11_10_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_11_11_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_11_12_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_11_13_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_11_14_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_11_15_sva_dfm <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_64_cse ) begin
      weight_port_read_out_data_11_0_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44;
      weight_port_read_out_data_11_1_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42;
      weight_port_read_out_data_11_2_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40;
      weight_port_read_out_data_11_3_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
      weight_port_read_out_data_11_4_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
      weight_port_read_out_data_11_5_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
      weight_port_read_out_data_11_6_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
      weight_port_read_out_data_11_7_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
      weight_port_read_out_data_11_8_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
      weight_port_read_out_data_11_9_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
      weight_port_read_out_data_11_10_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
      weight_port_read_out_data_11_11_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
      weight_port_read_out_data_11_12_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
      weight_port_read_out_data_11_13_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
      weight_port_read_out_data_11_14_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16;
      weight_port_read_out_data_11_15_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_8_0_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_8_1_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_8_2_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_8_3_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_8_4_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_8_5_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_8_6_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_8_7_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_8_8_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_8_9_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_8_10_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_8_11_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_8_12_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_8_13_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_8_14_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_8_15_sva_dfm <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_80_cse ) begin
      weight_port_read_out_data_8_0_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1;
      weight_port_read_out_data_8_1_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1;
      weight_port_read_out_data_8_2_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1;
      weight_port_read_out_data_8_3_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1;
      weight_port_read_out_data_8_4_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1;
      weight_port_read_out_data_8_5_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1;
      weight_port_read_out_data_8_6_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1;
      weight_port_read_out_data_8_7_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1;
      weight_port_read_out_data_8_8_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1;
      weight_port_read_out_data_8_9_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1;
      weight_port_read_out_data_8_10_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1;
      weight_port_read_out_data_8_11_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1;
      weight_port_read_out_data_8_12_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1;
      weight_port_read_out_data_8_13_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1;
      weight_port_read_out_data_8_14_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1;
      weight_port_read_out_data_8_15_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_15_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_7_8_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_7_14_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_7_9_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_7_13_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_7_10_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_7_12_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_7_11_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_7_7_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_7_0_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_7_6_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_7_1_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_7_5_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_7_2_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_7_4_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_7_3_sva_dfm <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_96_cse ) begin
      weight_port_read_out_data_7_15_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_7_8_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
      weight_port_read_out_data_7_14_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16;
      weight_port_read_out_data_7_9_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
      weight_port_read_out_data_7_13_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
      weight_port_read_out_data_7_10_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
      weight_port_read_out_data_7_12_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
      weight_port_read_out_data_7_11_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
      weight_port_read_out_data_7_7_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
      weight_port_read_out_data_7_0_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44;
      weight_port_read_out_data_7_6_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
      weight_port_read_out_data_7_1_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42;
      weight_port_read_out_data_7_5_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
      weight_port_read_out_data_7_2_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40;
      weight_port_read_out_data_7_4_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
      weight_port_read_out_data_7_3_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_6_7_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_6_0_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_6_6_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_6_1_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_6_5_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_6_2_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_6_4_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_6_3_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_6_15_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_6_8_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_6_14_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_6_9_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_6_13_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_6_10_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_6_12_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_6_11_sva_dfm <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_112_cse ) begin
      weight_port_read_out_data_6_7_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1;
      weight_port_read_out_data_6_0_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1;
      weight_port_read_out_data_6_6_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1;
      weight_port_read_out_data_6_1_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1;
      weight_port_read_out_data_6_5_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1;
      weight_port_read_out_data_6_2_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1;
      weight_port_read_out_data_6_4_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1;
      weight_port_read_out_data_6_3_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1;
      weight_port_read_out_data_6_15_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1;
      weight_port_read_out_data_6_8_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1;
      weight_port_read_out_data_6_14_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1;
      weight_port_read_out_data_6_9_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1;
      weight_port_read_out_data_6_13_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1;
      weight_port_read_out_data_6_10_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1;
      weight_port_read_out_data_6_12_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1;
      weight_port_read_out_data_6_11_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_8_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_5_9_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_5_10_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_5_11_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_5_12_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_5_13_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_5_14_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_5_15_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_5_0_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_5_1_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_5_2_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_5_3_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_5_4_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_5_5_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_5_6_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_5_7_sva_dfm <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_128_cse ) begin
      weight_port_read_out_data_5_8_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
      weight_port_read_out_data_5_9_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
      weight_port_read_out_data_5_10_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
      weight_port_read_out_data_5_11_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
      weight_port_read_out_data_5_12_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
      weight_port_read_out_data_5_13_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
      weight_port_read_out_data_5_14_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16;
      weight_port_read_out_data_5_15_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_5_0_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44;
      weight_port_read_out_data_5_1_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42;
      weight_port_read_out_data_5_2_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40;
      weight_port_read_out_data_5_3_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
      weight_port_read_out_data_5_4_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
      weight_port_read_out_data_5_5_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
      weight_port_read_out_data_5_6_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
      weight_port_read_out_data_5_7_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_0_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_4_1_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_4_2_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_4_3_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_4_4_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_4_5_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_4_6_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_4_7_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_4_8_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_4_9_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_4_10_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_4_11_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_4_12_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_4_13_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_4_14_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_4_15_sva_dfm <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_136_cse ) begin
      weight_port_read_out_data_4_0_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1;
      weight_port_read_out_data_4_1_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1;
      weight_port_read_out_data_4_2_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1;
      weight_port_read_out_data_4_3_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1;
      weight_port_read_out_data_4_4_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1;
      weight_port_read_out_data_4_5_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1;
      weight_port_read_out_data_4_6_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1;
      weight_port_read_out_data_4_7_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1;
      weight_port_read_out_data_4_8_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1;
      weight_port_read_out_data_4_9_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1;
      weight_port_read_out_data_4_10_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1;
      weight_port_read_out_data_4_11_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1;
      weight_port_read_out_data_4_12_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1;
      weight_port_read_out_data_4_13_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1;
      weight_port_read_out_data_4_14_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1;
      weight_port_read_out_data_4_15_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_8_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_3_9_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_3_10_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_3_11_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_3_12_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_3_13_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_3_14_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_3_15_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_3_0_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_3_1_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_3_2_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_3_3_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_3_4_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_3_5_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_3_6_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_3_7_sva_dfm <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_152_cse ) begin
      weight_port_read_out_data_3_8_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
      weight_port_read_out_data_3_9_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
      weight_port_read_out_data_3_10_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
      weight_port_read_out_data_3_11_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
      weight_port_read_out_data_3_12_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
      weight_port_read_out_data_3_13_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
      weight_port_read_out_data_3_14_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16;
      weight_port_read_out_data_3_15_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_3_0_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44;
      weight_port_read_out_data_3_1_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42;
      weight_port_read_out_data_3_2_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40;
      weight_port_read_out_data_3_3_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
      weight_port_read_out_data_3_4_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
      weight_port_read_out_data_3_5_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
      weight_port_read_out_data_3_6_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
      weight_port_read_out_data_3_7_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_0_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_2_1_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_2_2_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_2_3_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_2_4_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_2_5_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_2_6_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_2_7_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_2_8_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_2_9_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_2_10_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_2_11_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_2_12_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_2_13_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_2_14_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_2_15_sva_dfm <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_168_cse ) begin
      weight_port_read_out_data_2_0_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1;
      weight_port_read_out_data_2_1_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1;
      weight_port_read_out_data_2_2_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1;
      weight_port_read_out_data_2_3_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1;
      weight_port_read_out_data_2_4_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1;
      weight_port_read_out_data_2_5_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1;
      weight_port_read_out_data_2_6_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1;
      weight_port_read_out_data_2_7_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1;
      weight_port_read_out_data_2_8_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1;
      weight_port_read_out_data_2_9_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1;
      weight_port_read_out_data_2_10_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1;
      weight_port_read_out_data_2_11_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1;
      weight_port_read_out_data_2_12_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1;
      weight_port_read_out_data_2_13_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1;
      weight_port_read_out_data_2_14_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1;
      weight_port_read_out_data_2_15_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_1_8_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_1_9_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_1_10_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_1_11_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_1_12_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_1_13_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_1_14_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_1_15_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_1_0_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_1_1_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_1_2_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_1_3_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_1_4_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_1_5_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_1_6_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_1_7_sva_dfm <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_184_cse ) begin
      weight_port_read_out_data_1_8_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
      weight_port_read_out_data_1_9_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
      weight_port_read_out_data_1_10_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
      weight_port_read_out_data_1_11_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
      weight_port_read_out_data_1_12_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
      weight_port_read_out_data_1_13_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
      weight_port_read_out_data_1_14_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16;
      weight_port_read_out_data_1_15_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_1_0_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44;
      weight_port_read_out_data_1_1_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42;
      weight_port_read_out_data_1_2_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40;
      weight_port_read_out_data_1_3_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
      weight_port_read_out_data_1_4_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
      weight_port_read_out_data_1_5_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
      weight_port_read_out_data_1_6_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
      weight_port_read_out_data_1_7_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_8_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_0_9_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_0_10_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_0_11_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_0_12_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_0_13_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_0_14_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_0_15_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_0_0_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_0_1_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_0_2_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_0_3_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_0_4_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_0_5_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_0_6_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_0_7_sva_dfm <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_200_cse ) begin
      weight_port_read_out_data_0_8_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
      weight_port_read_out_data_0_9_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
      weight_port_read_out_data_0_10_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
      weight_port_read_out_data_0_11_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
      weight_port_read_out_data_0_12_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
      weight_port_read_out_data_0_13_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
      weight_port_read_out_data_0_14_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
      weight_port_read_out_data_0_15_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_2;
      weight_port_read_out_data_0_0_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_1_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
      weight_port_read_out_data_0_1_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_13_mx1w2;
      weight_port_read_out_data_0_2_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_12_mx1w2;
      weight_port_read_out_data_0_3_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_11_mx1w2;
      weight_port_read_out_data_0_4_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
      weight_port_read_out_data_0_5_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
      weight_port_read_out_data_0_6_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
      weight_port_read_out_data_0_7_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      accum_vector_data_15_sva <= 32'b00000000000000000000000000000000;
      accum_vector_data_14_sva <= 32'b00000000000000000000000000000000;
      accum_vector_data_13_sva <= 32'b00000000000000000000000000000000;
      accum_vector_data_12_sva <= 32'b00000000000000000000000000000000;
      act_port_reg_data_0_sva <= 20'b00000000000000000000;
      act_port_reg_data_11_sva <= 20'b00000000000000000000;
      act_port_reg_data_8_sva <= 20'b00000000000000000000;
      act_port_reg_data_7_sva <= 20'b00000000000000000000;
      while_and_30_itm_1 <= 1'b0;
    end
    else if ( accum_vector_data_and_9_cse ) begin
      accum_vector_data_15_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_15_cse;
      accum_vector_data_14_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_14_cse;
      accum_vector_data_13_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_13_cse;
      accum_vector_data_12_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_12_cse;
      act_port_reg_data_0_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_25_cse;
      act_port_reg_data_11_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_26_cse;
      act_port_reg_data_8_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_22_cse;
      act_port_reg_data_7_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_21_cse;
      while_and_30_itm_1 <= while_and_32_cse_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_reg_data_12_sva <= 20'b00000000000000000000;
      act_port_reg_data_13_sva <= 20'b00000000000000000000;
      act_port_reg_data_14_sva <= 20'b00000000000000000000;
      act_port_reg_data_15_sva <= 20'b00000000000000000000;
    end
    else if ( and_5872_cse ) begin
      act_port_reg_data_12_sva <= MUX_v_20_2_2(20'b00000000000000000000, while_while_mux1h_12_nl,
          PECore_UpdateFSM_switch_lp_not_36_nl);
      act_port_reg_data_13_sva <= MUX_v_20_2_2(20'b00000000000000000000, while_while_mux1h_13_nl,
          PECore_UpdateFSM_switch_lp_not_64_nl);
      act_port_reg_data_14_sva <= MUX_v_20_2_2(20'b00000000000000000000, while_while_mux1h_14_nl,
          PECore_UpdateFSM_switch_lp_not_63_nl);
      act_port_reg_data_15_sva <= MUX_v_20_2_2(20'b00000000000000000000, while_while_mux1h_15_nl,
          PECore_UpdateFSM_switch_lp_not_62_nl);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(or_dcpl | nor_499_cse)) ) begin
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva
          <= input_port_PopNB_mioi_ivld_mxwt;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mio_mrgout_dat_sva <= 169'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      PECore_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva
          <= 1'b0;
    end
    else if ( PECore_DecodeAxi_if_and_3_cse ) begin
      rva_in_PopNB_mio_mrgout_dat_sva <= rva_in_PopNB_mioi_idat_mxwt;
      PECore_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva
          <= rva_in_PopNB_mioi_ivld_mxwt;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      pe_config_is_valid_sva <= 1'b0;
      pe_config_is_cluster_sva <= 1'b0;
      pe_config_is_bias_sva <= 1'b0;
    end
    else if ( pe_config_is_valid_and_cse ) begin
      pe_config_is_valid_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[0];
      pe_config_is_cluster_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[16];
      pe_config_is_bias_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[24];
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      pe_config_is_zero_first_sva <= 1'b0;
      PECore_RunFSM_switch_lp_equal_tmp <= 1'b0;
      PECore_RunFSM_switch_lp_equal_tmp_2 <= 1'b0;
      PECore_RunFSM_switch_lp_equal_tmp_1 <= 1'b0;
    end
    else if ( pe_config_manager_counter_and_cse ) begin
      pe_config_is_zero_first_sva <= MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_mux_7_nl,
          pe_config_is_zero_first_sva_dfm_4_mx0, and_3991_nl);
      PECore_RunFSM_switch_lp_equal_tmp <= PECore_RunFSM_switch_lp_equal_tmp_3;
      PECore_RunFSM_switch_lp_equal_tmp_2 <= PECore_RunFSM_switch_lp_equal_tmp_4;
      PECore_RunFSM_switch_lp_equal_tmp_1 <= PECore_RunFSM_switch_lp_equal_tmp_5;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      pe_config_num_output_sva <= 8'b00000001;
      pe_config_num_manager_sva <= 4'b0001;
    end
    else if ( pe_config_num_output_and_cse ) begin
      pe_config_num_output_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[47:40];
      pe_config_num_manager_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[35:32];
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      pe_manager_zero_active_1_sva <= 1'b0;
    end
    else if ( PECoreRun_wen & PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8
        & PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_31 &
        (rva_in_PopNB_mio_mrgout_dat_sva_1[168]) & rva_in_PopNB_mioi_ivld_mxwt &
        (~ or_tmp_2232) ) begin
      pe_manager_zero_active_1_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[0];
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      pe_manager_zero_active_0_sva <= 1'b0;
    end
    else if ( PECoreRun_wen & PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6
        & PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_31 &
        (rva_in_PopNB_mio_mrgout_dat_sva_1[168]) & rva_in_PopNB_mioi_ivld_mxwt &
        (~ or_tmp_2232) ) begin
      pe_manager_zero_active_0_sva <= rva_in_PopNB_mio_mrgout_dat_sva_1[0];
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      pe_config_input_counter_sva <= 8'b00000000;
    end
    else if ( PECoreRun_wen & (~((or_dcpl_724 & and_4031_m1c) | nor_499_cse)) ) begin
      pe_config_input_counter_sva <= MUX_v_8_2_2(pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl,
          ({{7{PECore_DecodeAxiWrite_case_4_switch_lp_or_6_cse_1}}, PECore_DecodeAxiWrite_case_4_switch_lp_or_6_cse_1}),
          PECore_UpdateFSM_switch_lp_and_nl);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      pe_config_output_counter_sva <= 8'b00000000;
    end
    else if ( (~((state_2_0_sva_0 | state_2_0_sva_1 | pe_config_UpdateManagerCounter_if_unequal_tmp
        | (~ state_2_0_sva_2) | (operator_4_false_acc_tmp[4])) & ((~ (rva_in_PopNB_mioi_idat_mxwt[150]))
        | (~ rva_in_PopNB_mioi_ivld_mxwt) | (rva_in_PopNB_mioi_idat_mxwt[151]) |
        (rva_in_PopNB_mioi_idat_mxwt[149]) | is_start_sva | (rva_in_PopNB_mioi_idat_mxwt[148])
        | (~ (rva_in_PopNB_mioi_idat_mxwt[168])) | (~ (rva_in_PopNB_mioi_idat_mxwt[132]))
        | (rva_in_PopNB_mioi_idat_mxwt[133]) | (rva_in_PopNB_mioi_idat_mxwt[134])
        | (rva_in_PopNB_mioi_idat_mxwt[147]) | (rva_in_PopNB_mioi_idat_mxwt[146])
        | (rva_in_PopNB_mioi_idat_mxwt[145]) | (rva_in_PopNB_mioi_idat_mxwt[144])
        | (rva_in_PopNB_mioi_idat_mxwt[143]) | (rva_in_PopNB_mioi_idat_mxwt[142])
        | (rva_in_PopNB_mioi_idat_mxwt[141]) | (rva_in_PopNB_mioi_idat_mxwt[140])
        | (rva_in_PopNB_mioi_idat_mxwt[139]) | (rva_in_PopNB_mioi_idat_mxwt[138])
        | (rva_in_PopNB_mioi_idat_mxwt[137]) | (rva_in_PopNB_mioi_idat_mxwt[136])
        | (rva_in_PopNB_mioi_idat_mxwt[135])))) & (fsm_output[1]) & PECoreRun_wen
        ) begin
      pe_config_output_counter_sva <= MUX_v_8_2_2(pe_config_output_counter_sva_dfm_4_mx0,
          pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl,
          and_4037_nl);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm <= 1'b0;
    end
    else if ( PECoreRun_wen & (fsm_output[1]) & weight_mem_read_arbxbar_xbar_for_3_1_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm <= weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm <= 1'b0;
    end
    else if ( PECoreRun_wen & (fsm_output[1]) & weight_mem_read_arbxbar_xbar_for_3_2_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm <= weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm <= 1'b0;
    end
    else if ( PECoreRun_wen & (fsm_output[1]) & weight_mem_read_arbxbar_xbar_for_3_3_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm <= weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm <= 1'b0;
    end
    else if ( PECoreRun_wen & (fsm_output[1]) & weight_mem_read_arbxbar_xbar_for_3_4_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm <= weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm <= 1'b0;
    end
    else if ( PECoreRun_wen & (fsm_output[1]) & weight_mem_read_arbxbar_xbar_for_3_5_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm <= weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm <= 1'b0;
    end
    else if ( PECoreRun_wen & (fsm_output[1]) & weight_mem_read_arbxbar_xbar_for_3_6_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm <= weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm <= 1'b0;
    end
    else if ( PECoreRun_wen & (fsm_output[1]) & weight_mem_read_arbxbar_xbar_for_3_7_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm <= weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm <= 1'b0;
    end
    else if ( PECoreRun_wen & (fsm_output[1]) & weight_mem_read_arbxbar_xbar_for_3_8_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm <= weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm <= 1'b0;
    end
    else if ( PECoreRun_wen & (fsm_output[1]) & weight_mem_read_arbxbar_xbar_for_3_9_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm <= weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm <= 1'b0;
    end
    else if ( PECoreRun_wen & (fsm_output[1]) & weight_mem_read_arbxbar_xbar_for_3_10_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm <= weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm <= 1'b0;
    end
    else if ( PECoreRun_wen & (fsm_output[1]) & weight_mem_read_arbxbar_xbar_for_3_11_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm <= weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm <= 1'b0;
    end
    else if ( PECoreRun_wen & (fsm_output[1]) & weight_mem_read_arbxbar_xbar_for_3_12_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm <= weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm <= 1'b0;
    end
    else if ( PECoreRun_wen & (fsm_output[1]) & weight_mem_read_arbxbar_xbar_for_3_13_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm <= weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm <= 1'b0;
    end
    else if ( PECoreRun_wen & (fsm_output[1]) & weight_mem_read_arbxbar_xbar_for_3_14_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm <= weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm <= 1'b0;
    end
    else if ( PECoreRun_wen & (fsm_output[1]) & weight_mem_read_arbxbar_xbar_for_3_15_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm <= weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_14
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_13
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_12
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_11
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_10
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_9
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_8
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_7
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_0
          <= 1'b0;
      weight_mem_read_arbxbar_arbiters_next_0_15_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_14_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_13_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_12_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_11_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_10_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_9_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_6_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_8_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_7_sva <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_ssc
        ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_14
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_14;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_13
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_13;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_12
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_12;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_11
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_11;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_10
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_10;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_9
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_9;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_8
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_8;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_7
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_7;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_6
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_6;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_5
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_5;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_4
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_4;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_3
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_3;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_2
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_2;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_1
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_1;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_0
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_0;
      weight_mem_read_arbxbar_arbiters_next_0_15_sva <= Arbiter_16U_Roundrobin_pick_if_1_not_251;
      weight_mem_read_arbxbar_arbiters_next_0_14_sva <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_14
          | Arbiter_16U_Roundrobin_pick_if_1_not_251;
      weight_mem_read_arbxbar_arbiters_next_0_1_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
          | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_251;
      weight_mem_read_arbxbar_arbiters_next_0_13_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_251;
      weight_mem_read_arbxbar_arbiters_next_0_2_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_251;
      weight_mem_read_arbxbar_arbiters_next_0_12_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_251;
      weight_mem_read_arbxbar_arbiters_next_0_3_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_251;
      weight_mem_read_arbxbar_arbiters_next_0_11_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_251;
      weight_mem_read_arbxbar_arbiters_next_0_4_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_251;
      weight_mem_read_arbxbar_arbiters_next_0_10_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_251;
      weight_mem_read_arbxbar_arbiters_next_0_5_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_251;
      weight_mem_read_arbxbar_arbiters_next_0_9_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_251;
      weight_mem_read_arbxbar_arbiters_next_0_6_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_251;
      weight_mem_read_arbxbar_arbiters_next_0_8_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_251;
      weight_mem_read_arbxbar_arbiters_next_0_7_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_251;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_14
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_13
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_12
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_11
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_10
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_9
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_8
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_7
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_0
          <= 1'b0;
      weight_mem_read_arbxbar_arbiters_next_1_15_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_14_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_13_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_12_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_11_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_10_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_9_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_6_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_8_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_7_sva <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_1_ssc
        ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_14
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_14;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_13
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_13;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_12
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_12;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_11
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_11;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_10
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_10;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_9
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_9;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_8
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_8;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_7
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_7;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_6
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_6;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_5
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_5;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_4
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_4;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_3
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_3;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_2
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_2;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_1
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_1;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_0
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_0;
      weight_mem_read_arbxbar_arbiters_next_1_15_sva <= Arbiter_16U_Roundrobin_pick_if_1_not_249;
      weight_mem_read_arbxbar_arbiters_next_1_14_sva <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_14
          | Arbiter_16U_Roundrobin_pick_if_1_not_249;
      weight_mem_read_arbxbar_arbiters_next_1_1_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
          | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_249;
      weight_mem_read_arbxbar_arbiters_next_1_13_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_249;
      weight_mem_read_arbxbar_arbiters_next_1_2_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_249;
      weight_mem_read_arbxbar_arbiters_next_1_12_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_249;
      weight_mem_read_arbxbar_arbiters_next_1_3_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_249;
      weight_mem_read_arbxbar_arbiters_next_1_11_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_249;
      weight_mem_read_arbxbar_arbiters_next_1_4_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_249;
      weight_mem_read_arbxbar_arbiters_next_1_10_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_249;
      weight_mem_read_arbxbar_arbiters_next_1_5_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_249;
      weight_mem_read_arbxbar_arbiters_next_1_9_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_249;
      weight_mem_read_arbxbar_arbiters_next_1_6_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_249;
      weight_mem_read_arbxbar_arbiters_next_1_8_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_249;
      weight_mem_read_arbxbar_arbiters_next_1_7_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_249;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_14
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_13
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_12
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_11
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_10
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_9
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_8
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_7
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_0
          <= 1'b0;
      weight_mem_read_arbxbar_arbiters_next_2_15_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_14_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_13_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_12_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_11_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_10_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_9_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_6_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_8_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_7_sva <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_2_ssc
        ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_14
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_14;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_13
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_13;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_12
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_12;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_11
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_11;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_10
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_10;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_9
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_9;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_8
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_8;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_7
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_7;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_6
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_6;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_5
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_5;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_4
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_4;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_3
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_3;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_2
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_2;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_1
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_1;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_0
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_0;
      weight_mem_read_arbxbar_arbiters_next_2_15_sva <= Arbiter_16U_Roundrobin_pick_if_1_not_247;
      weight_mem_read_arbxbar_arbiters_next_2_14_sva <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_14
          | Arbiter_16U_Roundrobin_pick_if_1_not_247;
      weight_mem_read_arbxbar_arbiters_next_2_1_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
          | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_247;
      weight_mem_read_arbxbar_arbiters_next_2_13_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_247;
      weight_mem_read_arbxbar_arbiters_next_2_2_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_247;
      weight_mem_read_arbxbar_arbiters_next_2_12_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_247;
      weight_mem_read_arbxbar_arbiters_next_2_3_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_247;
      weight_mem_read_arbxbar_arbiters_next_2_11_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_247;
      weight_mem_read_arbxbar_arbiters_next_2_4_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_247;
      weight_mem_read_arbxbar_arbiters_next_2_10_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_247;
      weight_mem_read_arbxbar_arbiters_next_2_5_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_247;
      weight_mem_read_arbxbar_arbiters_next_2_9_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_247;
      weight_mem_read_arbxbar_arbiters_next_2_6_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_247;
      weight_mem_read_arbxbar_arbiters_next_2_8_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_247;
      weight_mem_read_arbxbar_arbiters_next_2_7_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_247;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_14
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_13
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_12
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_11
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_10
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_9
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_8
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_7
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_0
          <= 1'b0;
      weight_mem_read_arbxbar_arbiters_next_3_15_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_14_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_13_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_12_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_11_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_10_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_9_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_6_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_8_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_7_sva <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_3_ssc
        ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_14
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_14;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_13
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_13;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_12
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_12;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_11
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_11;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_10
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_10;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_9
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_9;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_8
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_8;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_7
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_7;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_6
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_6;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_5
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_5;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_4
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_4;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_3
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_3;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_2
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_2;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_1
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_1;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_0
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_0;
      weight_mem_read_arbxbar_arbiters_next_3_15_sva <= Arbiter_16U_Roundrobin_pick_if_1_not_259;
      weight_mem_read_arbxbar_arbiters_next_3_14_sva <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_14
          | Arbiter_16U_Roundrobin_pick_if_1_not_259;
      weight_mem_read_arbxbar_arbiters_next_3_1_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
          | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_259;
      weight_mem_read_arbxbar_arbiters_next_3_13_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_259;
      weight_mem_read_arbxbar_arbiters_next_3_2_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_259;
      weight_mem_read_arbxbar_arbiters_next_3_12_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_259;
      weight_mem_read_arbxbar_arbiters_next_3_3_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_259;
      weight_mem_read_arbxbar_arbiters_next_3_11_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_259;
      weight_mem_read_arbxbar_arbiters_next_3_4_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_259;
      weight_mem_read_arbxbar_arbiters_next_3_10_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_259;
      weight_mem_read_arbxbar_arbiters_next_3_5_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_259;
      weight_mem_read_arbxbar_arbiters_next_3_9_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_259;
      weight_mem_read_arbxbar_arbiters_next_3_6_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_259;
      weight_mem_read_arbxbar_arbiters_next_3_8_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_259;
      weight_mem_read_arbxbar_arbiters_next_3_7_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_259;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_14
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_13
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_12
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_11
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_10
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_9
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_8
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_7
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_0
          <= 1'b0;
      weight_mem_read_arbxbar_arbiters_next_4_15_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_14_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_13_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_12_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_11_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_10_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_9_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_6_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_8_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_7_sva <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_4_ssc
        ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_14
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_14;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_13
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_13;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_12
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_12;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_11
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_11;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_10
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_10;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_9
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_9;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_8
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_8;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_7
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_7;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_6
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_6;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_5
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_5;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_4
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_4;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_3
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_3;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_2
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_2;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_1
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_1;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_0
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_0;
      weight_mem_read_arbxbar_arbiters_next_4_15_sva <= Arbiter_16U_Roundrobin_pick_if_1_not_257;
      weight_mem_read_arbxbar_arbiters_next_4_14_sva <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_14
          | Arbiter_16U_Roundrobin_pick_if_1_not_257;
      weight_mem_read_arbxbar_arbiters_next_4_1_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
          | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_257;
      weight_mem_read_arbxbar_arbiters_next_4_13_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_257;
      weight_mem_read_arbxbar_arbiters_next_4_2_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_257;
      weight_mem_read_arbxbar_arbiters_next_4_12_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_257;
      weight_mem_read_arbxbar_arbiters_next_4_3_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_257;
      weight_mem_read_arbxbar_arbiters_next_4_11_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_257;
      weight_mem_read_arbxbar_arbiters_next_4_4_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_257;
      weight_mem_read_arbxbar_arbiters_next_4_10_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_257;
      weight_mem_read_arbxbar_arbiters_next_4_5_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_257;
      weight_mem_read_arbxbar_arbiters_next_4_9_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_257;
      weight_mem_read_arbxbar_arbiters_next_4_6_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_257;
      weight_mem_read_arbxbar_arbiters_next_4_8_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_257;
      weight_mem_read_arbxbar_arbiters_next_4_7_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_257;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_14
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_13
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_12
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_11
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_10
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_9
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_8
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_7
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_0
          <= 1'b0;
      weight_mem_read_arbxbar_arbiters_next_5_15_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_14_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_13_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_12_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_11_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_10_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_9_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_6_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_8_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_7_sva <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_5_ssc
        ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_14
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_14;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_13
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_13;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_12
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_12;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_11
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_11;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_10
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_10;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_9
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_9;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_8
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_8;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_7
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_7;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_6
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_6;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_5
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_5;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_4
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_4;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_3
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_3;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_2
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_2;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_1
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_1;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_0
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_0;
      weight_mem_read_arbxbar_arbiters_next_5_15_sva <= Arbiter_16U_Roundrobin_pick_if_1_not_245;
      weight_mem_read_arbxbar_arbiters_next_5_14_sva <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_14
          | Arbiter_16U_Roundrobin_pick_if_1_not_245;
      weight_mem_read_arbxbar_arbiters_next_5_1_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
          | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_245;
      weight_mem_read_arbxbar_arbiters_next_5_13_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_245;
      weight_mem_read_arbxbar_arbiters_next_5_2_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_245;
      weight_mem_read_arbxbar_arbiters_next_5_12_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_245;
      weight_mem_read_arbxbar_arbiters_next_5_3_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_245;
      weight_mem_read_arbxbar_arbiters_next_5_11_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_245;
      weight_mem_read_arbxbar_arbiters_next_5_4_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_245;
      weight_mem_read_arbxbar_arbiters_next_5_10_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_245;
      weight_mem_read_arbxbar_arbiters_next_5_5_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_245;
      weight_mem_read_arbxbar_arbiters_next_5_9_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_245;
      weight_mem_read_arbxbar_arbiters_next_5_6_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_245;
      weight_mem_read_arbxbar_arbiters_next_5_8_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_245;
      weight_mem_read_arbxbar_arbiters_next_5_7_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_245;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_14
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_13
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_12
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_11
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_10
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_9
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_8
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_7
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_0
          <= 1'b0;
      weight_mem_read_arbxbar_arbiters_next_6_15_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_14_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_13_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_12_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_11_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_10_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_9_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_6_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_8_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_7_sva <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_6_ssc
        ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_14
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_14;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_13
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_13;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_12
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_12;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_11
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_11;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_10
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_10;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_9
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_9;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_8
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_8;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_7
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_7;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_6
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_6;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_5
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_5;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_4
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_4;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_3
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_3;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_2
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_2;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_1
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_1;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_0
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_0;
      weight_mem_read_arbxbar_arbiters_next_6_15_sva <= Arbiter_16U_Roundrobin_pick_if_1_not_269;
      weight_mem_read_arbxbar_arbiters_next_6_14_sva <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_14
          | Arbiter_16U_Roundrobin_pick_if_1_not_269;
      weight_mem_read_arbxbar_arbiters_next_6_1_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
          | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_269;
      weight_mem_read_arbxbar_arbiters_next_6_13_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_269;
      weight_mem_read_arbxbar_arbiters_next_6_2_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_269;
      weight_mem_read_arbxbar_arbiters_next_6_12_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_269;
      weight_mem_read_arbxbar_arbiters_next_6_3_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_269;
      weight_mem_read_arbxbar_arbiters_next_6_11_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_269;
      weight_mem_read_arbxbar_arbiters_next_6_4_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_269;
      weight_mem_read_arbxbar_arbiters_next_6_10_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_269;
      weight_mem_read_arbxbar_arbiters_next_6_5_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_269;
      weight_mem_read_arbxbar_arbiters_next_6_9_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_269;
      weight_mem_read_arbxbar_arbiters_next_6_6_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_269;
      weight_mem_read_arbxbar_arbiters_next_6_8_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_269;
      weight_mem_read_arbxbar_arbiters_next_6_7_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_269;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_14
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_13
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_12
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_11
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_10
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_9
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_8
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_7
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_0
          <= 1'b0;
      weight_mem_read_arbxbar_arbiters_next_7_15_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_14_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_13_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_12_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_11_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_10_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_9_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_6_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_8_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_7_sva <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_7_ssc
        ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_14
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_14;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_13
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_13;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_12
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_12;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_11
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_11;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_10
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_10;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_9
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_9;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_8
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_8;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_7
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_7;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_6
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_6;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_5
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_5;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_4
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_4;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_3
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_3;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_2
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_2;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_1
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_1;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_0
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_0;
      weight_mem_read_arbxbar_arbiters_next_7_15_sva <= Arbiter_16U_Roundrobin_pick_if_1_not_261;
      weight_mem_read_arbxbar_arbiters_next_7_14_sva <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_14
          | Arbiter_16U_Roundrobin_pick_if_1_not_261;
      weight_mem_read_arbxbar_arbiters_next_7_1_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
          | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_261;
      weight_mem_read_arbxbar_arbiters_next_7_13_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_261;
      weight_mem_read_arbxbar_arbiters_next_7_2_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_261;
      weight_mem_read_arbxbar_arbiters_next_7_12_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_261;
      weight_mem_read_arbxbar_arbiters_next_7_3_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_261;
      weight_mem_read_arbxbar_arbiters_next_7_11_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_261;
      weight_mem_read_arbxbar_arbiters_next_7_4_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_261;
      weight_mem_read_arbxbar_arbiters_next_7_10_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_261;
      weight_mem_read_arbxbar_arbiters_next_7_5_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_261;
      weight_mem_read_arbxbar_arbiters_next_7_9_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_261;
      weight_mem_read_arbxbar_arbiters_next_7_6_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_261;
      weight_mem_read_arbxbar_arbiters_next_7_8_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_261;
      weight_mem_read_arbxbar_arbiters_next_7_7_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_261;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_14
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_13
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_12
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_11
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_10
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_9
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_8
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_7
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_0
          <= 1'b0;
      weight_mem_read_arbxbar_arbiters_next_8_15_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_8_14_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_8_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_8_13_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_8_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_8_12_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_8_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_8_11_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_8_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_8_10_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_8_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_8_9_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_8_6_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_8_8_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_8_7_sva <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_8_ssc
        ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_14
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_14;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_13
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_13;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_12
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_12;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_11
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_11;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_10
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_10;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_9
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_9;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_8
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_8;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_7
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_7;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_6
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_6;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_5
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_5;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_4
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_4;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_3
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_3;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_2
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_2;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_1
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_1;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_0
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_0;
      weight_mem_read_arbxbar_arbiters_next_8_15_sva <= Arbiter_16U_Roundrobin_pick_if_1_not_267;
      weight_mem_read_arbxbar_arbiters_next_8_14_sva <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_14
          | Arbiter_16U_Roundrobin_pick_if_1_not_267;
      weight_mem_read_arbxbar_arbiters_next_8_1_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
          | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_267;
      weight_mem_read_arbxbar_arbiters_next_8_13_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_267;
      weight_mem_read_arbxbar_arbiters_next_8_2_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_267;
      weight_mem_read_arbxbar_arbiters_next_8_12_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_267;
      weight_mem_read_arbxbar_arbiters_next_8_3_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_267;
      weight_mem_read_arbxbar_arbiters_next_8_11_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_267;
      weight_mem_read_arbxbar_arbiters_next_8_4_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_267;
      weight_mem_read_arbxbar_arbiters_next_8_10_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_267;
      weight_mem_read_arbxbar_arbiters_next_8_5_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_267;
      weight_mem_read_arbxbar_arbiters_next_8_9_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_267;
      weight_mem_read_arbxbar_arbiters_next_8_6_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_267;
      weight_mem_read_arbxbar_arbiters_next_8_8_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_267;
      weight_mem_read_arbxbar_arbiters_next_8_7_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_267;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_14
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_13
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_12
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_11
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_10
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_9
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_8
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_7
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_0
          <= 1'b0;
      weight_mem_read_arbxbar_arbiters_next_9_15_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_9_14_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_9_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_9_13_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_9_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_9_12_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_9_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_9_11_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_9_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_9_10_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_9_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_9_9_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_9_6_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_9_8_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_9_7_sva <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_9_ssc
        ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_14
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_14;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_13
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_13;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_12
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_12;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_11
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_11;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_10
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_10;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_9
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_9;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_8
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_8;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_7
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_7;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_6
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_6;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_5
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_5;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_4
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_4;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_3
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_3;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_2
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_2;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_1
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_1;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_0
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_0;
      weight_mem_read_arbxbar_arbiters_next_9_15_sva <= Arbiter_16U_Roundrobin_pick_if_1_not_253;
      weight_mem_read_arbxbar_arbiters_next_9_14_sva <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_14
          | Arbiter_16U_Roundrobin_pick_if_1_not_253;
      weight_mem_read_arbxbar_arbiters_next_9_1_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
          | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_253;
      weight_mem_read_arbxbar_arbiters_next_9_13_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_253;
      weight_mem_read_arbxbar_arbiters_next_9_2_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_253;
      weight_mem_read_arbxbar_arbiters_next_9_12_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_253;
      weight_mem_read_arbxbar_arbiters_next_9_3_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_253;
      weight_mem_read_arbxbar_arbiters_next_9_11_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_253;
      weight_mem_read_arbxbar_arbiters_next_9_4_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_253;
      weight_mem_read_arbxbar_arbiters_next_9_10_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_253;
      weight_mem_read_arbxbar_arbiters_next_9_5_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_253;
      weight_mem_read_arbxbar_arbiters_next_9_9_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_253;
      weight_mem_read_arbxbar_arbiters_next_9_6_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_253;
      weight_mem_read_arbxbar_arbiters_next_9_8_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_253;
      weight_mem_read_arbxbar_arbiters_next_9_7_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_253;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_14
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_13
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_12
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_11
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_10
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_9
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_8
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_7
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_0
          <= 1'b0;
      weight_mem_read_arbxbar_arbiters_next_10_15_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_10_14_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_10_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_10_13_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_10_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_10_12_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_10_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_10_11_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_10_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_10_10_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_10_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_10_9_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_10_6_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_10_8_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_10_7_sva <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_10_ssc
        ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_14
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_14;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_13
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_13;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_12
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_12;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_11
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_11;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_10
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_10;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_9
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_9;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_8
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_8;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_7
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_7;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_6
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_6;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_5
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_5;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_4
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_4;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_3
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_3;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_2
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_2;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_1
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_1;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_0
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_0;
      weight_mem_read_arbxbar_arbiters_next_10_15_sva <= Arbiter_16U_Roundrobin_pick_if_1_not_263;
      weight_mem_read_arbxbar_arbiters_next_10_14_sva <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_14
          | Arbiter_16U_Roundrobin_pick_if_1_not_263;
      weight_mem_read_arbxbar_arbiters_next_10_1_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
          | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_263;
      weight_mem_read_arbxbar_arbiters_next_10_13_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_263;
      weight_mem_read_arbxbar_arbiters_next_10_2_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_263;
      weight_mem_read_arbxbar_arbiters_next_10_12_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_263;
      weight_mem_read_arbxbar_arbiters_next_10_3_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_263;
      weight_mem_read_arbxbar_arbiters_next_10_11_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_263;
      weight_mem_read_arbxbar_arbiters_next_10_4_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_263;
      weight_mem_read_arbxbar_arbiters_next_10_10_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_263;
      weight_mem_read_arbxbar_arbiters_next_10_5_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_263;
      weight_mem_read_arbxbar_arbiters_next_10_9_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_263;
      weight_mem_read_arbxbar_arbiters_next_10_6_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_263;
      weight_mem_read_arbxbar_arbiters_next_10_8_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_263;
      weight_mem_read_arbxbar_arbiters_next_10_7_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_263;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_14
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_13
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_12
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_11
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_10
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_9
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_8
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_7
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_0
          <= 1'b0;
      weight_mem_read_arbxbar_arbiters_next_11_15_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_11_14_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_11_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_11_13_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_11_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_11_12_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_11_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_11_11_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_11_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_11_10_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_11_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_11_9_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_11_6_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_11_8_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_11_7_sva <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_11_ssc
        ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_14
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_14;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_13
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_13;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_12
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_12;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_11
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_11;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_10
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_10;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_9
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_9;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_8
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_8;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_7
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_7;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_6
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_6;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_5
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_5;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_4
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_4;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_3
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_3;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_2
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_2;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_1
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_1;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_0
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_0;
      weight_mem_read_arbxbar_arbiters_next_11_15_sva <= Arbiter_16U_Roundrobin_pick_if_1_not_271;
      weight_mem_read_arbxbar_arbiters_next_11_14_sva <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_14
          | Arbiter_16U_Roundrobin_pick_if_1_not_271;
      weight_mem_read_arbxbar_arbiters_next_11_1_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
          | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_271;
      weight_mem_read_arbxbar_arbiters_next_11_13_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_271;
      weight_mem_read_arbxbar_arbiters_next_11_2_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_271;
      weight_mem_read_arbxbar_arbiters_next_11_12_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_271;
      weight_mem_read_arbxbar_arbiters_next_11_3_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_271;
      weight_mem_read_arbxbar_arbiters_next_11_11_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_271;
      weight_mem_read_arbxbar_arbiters_next_11_4_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_271;
      weight_mem_read_arbxbar_arbiters_next_11_10_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_271;
      weight_mem_read_arbxbar_arbiters_next_11_5_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_271;
      weight_mem_read_arbxbar_arbiters_next_11_9_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_271;
      weight_mem_read_arbxbar_arbiters_next_11_6_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_271;
      weight_mem_read_arbxbar_arbiters_next_11_8_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_271;
      weight_mem_read_arbxbar_arbiters_next_11_7_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_271;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_14
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_13
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_12
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_11
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_10
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_9
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_8
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_7
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_0
          <= 1'b0;
      weight_mem_read_arbxbar_arbiters_next_12_15_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_12_14_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_12_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_12_13_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_12_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_12_12_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_12_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_12_11_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_12_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_12_10_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_12_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_12_9_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_12_6_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_12_8_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_12_7_sva <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_12_ssc
        ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_14
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_14;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_13
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_13;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_12
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_12;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_11
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_11;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_10
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_10;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_9
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_9;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_8
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_8;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_7
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_7;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_6
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_6;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_5
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_5;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_4
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_4;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_3
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_3;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_2
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_2;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_1
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_1;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_0
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_0;
      weight_mem_read_arbxbar_arbiters_next_12_15_sva <= Arbiter_16U_Roundrobin_pick_if_1_not_265;
      weight_mem_read_arbxbar_arbiters_next_12_14_sva <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_14
          | Arbiter_16U_Roundrobin_pick_if_1_not_265;
      weight_mem_read_arbxbar_arbiters_next_12_1_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
          | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_265;
      weight_mem_read_arbxbar_arbiters_next_12_13_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_265;
      weight_mem_read_arbxbar_arbiters_next_12_2_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_265;
      weight_mem_read_arbxbar_arbiters_next_12_12_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_265;
      weight_mem_read_arbxbar_arbiters_next_12_3_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_265;
      weight_mem_read_arbxbar_arbiters_next_12_11_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_265;
      weight_mem_read_arbxbar_arbiters_next_12_4_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_265;
      weight_mem_read_arbxbar_arbiters_next_12_10_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_265;
      weight_mem_read_arbxbar_arbiters_next_12_5_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_265;
      weight_mem_read_arbxbar_arbiters_next_12_9_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_265;
      weight_mem_read_arbxbar_arbiters_next_12_6_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_265;
      weight_mem_read_arbxbar_arbiters_next_12_8_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_265;
      weight_mem_read_arbxbar_arbiters_next_12_7_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_265;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_14
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_13
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_12
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_11
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_10
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_9
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_8
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_7
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_0
          <= 1'b0;
      weight_mem_read_arbxbar_arbiters_next_13_15_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_13_14_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_13_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_13_13_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_13_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_13_12_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_13_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_13_11_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_13_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_13_10_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_13_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_13_9_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_13_6_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_13_8_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_13_7_sva <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_13_ssc
        ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_14
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_14;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_13
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_13;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_12
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_12;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_11
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_11;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_10
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_10;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_9
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_9;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_8
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_8;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_7
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_7;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_6
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_6;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_5
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_5;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_4
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_4;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_3
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_3;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_2
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_2;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_1
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_1;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_0
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_0;
      weight_mem_read_arbxbar_arbiters_next_13_15_sva <= Arbiter_16U_Roundrobin_pick_if_1_not_241;
      weight_mem_read_arbxbar_arbiters_next_13_14_sva <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_14
          | Arbiter_16U_Roundrobin_pick_if_1_not_241;
      weight_mem_read_arbxbar_arbiters_next_13_1_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
          | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_241;
      weight_mem_read_arbxbar_arbiters_next_13_13_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_241;
      weight_mem_read_arbxbar_arbiters_next_13_2_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_241;
      weight_mem_read_arbxbar_arbiters_next_13_12_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_241;
      weight_mem_read_arbxbar_arbiters_next_13_3_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_241;
      weight_mem_read_arbxbar_arbiters_next_13_11_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_241;
      weight_mem_read_arbxbar_arbiters_next_13_4_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_241;
      weight_mem_read_arbxbar_arbiters_next_13_10_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_241;
      weight_mem_read_arbxbar_arbiters_next_13_5_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_241;
      weight_mem_read_arbxbar_arbiters_next_13_9_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_241;
      weight_mem_read_arbxbar_arbiters_next_13_6_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_241;
      weight_mem_read_arbxbar_arbiters_next_13_8_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_241;
      weight_mem_read_arbxbar_arbiters_next_13_7_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_241;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_14
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_13
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_12
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_11
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_10
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_9
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_8
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_7
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_0
          <= 1'b0;
      weight_mem_read_arbxbar_arbiters_next_14_15_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_14_14_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_14_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_14_13_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_14_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_14_12_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_14_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_14_11_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_14_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_14_10_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_14_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_14_9_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_14_6_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_14_8_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_14_7_sva <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_14_ssc
        ) begin
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_14
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_14;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_13
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_13;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_12
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_12;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_11
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_11;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_10
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_10;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_9
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_9;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_8
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_8;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_7
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_7;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_6
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_6;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_5
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_5;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_4
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_4;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_3
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_3;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_2
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_2;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_1
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_1;
      nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_0
          <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_0;
      weight_mem_read_arbxbar_arbiters_next_14_15_sva <= Arbiter_16U_Roundrobin_pick_if_1_not_255;
      weight_mem_read_arbxbar_arbiters_next_14_14_sva <= nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_14
          | Arbiter_16U_Roundrobin_pick_if_1_not_255;
      weight_mem_read_arbxbar_arbiters_next_14_1_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
          | nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_255;
      weight_mem_read_arbxbar_arbiters_next_14_13_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_255;
      weight_mem_read_arbxbar_arbiters_next_14_2_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_255;
      weight_mem_read_arbxbar_arbiters_next_14_12_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_255;
      weight_mem_read_arbxbar_arbiters_next_14_3_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_255;
      weight_mem_read_arbxbar_arbiters_next_14_11_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_255;
      weight_mem_read_arbxbar_arbiters_next_14_4_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_255;
      weight_mem_read_arbxbar_arbiters_next_14_10_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_255;
      weight_mem_read_arbxbar_arbiters_next_14_5_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_255;
      weight_mem_read_arbxbar_arbiters_next_14_9_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_255;
      weight_mem_read_arbxbar_arbiters_next_14_6_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_255;
      weight_mem_read_arbxbar_arbiters_next_14_8_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_255;
      weight_mem_read_arbxbar_arbiters_next_14_7_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_255;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd
          <= 1'b0;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_1
          <= 1'b0;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_2
          <= 1'b0;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_3
          <= 1'b0;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_4
          <= 1'b0;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_5
          <= 1'b0;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_6
          <= 1'b0;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_7
          <= 1'b0;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_8
          <= 1'b0;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_9
          <= 1'b0;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_10
          <= 1'b0;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_11
          <= 1'b0;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_12
          <= 1'b0;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_13
          <= 1'b0;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_14
          <= 1'b0;
      weight_mem_read_arbxbar_arbiters_next_15_15_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_15_14_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_15_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_15_13_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_15_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_15_12_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_15_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_15_11_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_15_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_15_10_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_15_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_15_9_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_15_6_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_15_8_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_15_7_sva <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_15_cse
        ) begin
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd
          <= weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_itm;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_1
          <= weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_1_itm;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_2
          <= weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_2_itm;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_3
          <= weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_3_itm;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_4
          <= weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_4_itm;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_5
          <= weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_5_itm;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_6
          <= weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_6_itm;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_7
          <= weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_7_itm;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_8
          <= weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_8_itm;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_9
          <= weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_9_itm;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_10
          <= weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_10_itm;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_11
          <= weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_11_itm;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_12
          <= weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_12_itm;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_13
          <= weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_13_itm;
      reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_14
          <= weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_14_itm;
      weight_mem_read_arbxbar_arbiters_next_15_15_sva <= Arbiter_16U_Roundrobin_pick_if_1_not_243;
      weight_mem_read_arbxbar_arbiters_next_15_14_sva <= weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_itm
          | Arbiter_16U_Roundrobin_pick_if_1_not_243;
      weight_mem_read_arbxbar_arbiters_next_15_1_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
          | weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_13_itm
          | Arbiter_16U_Roundrobin_pick_if_1_not_243;
      weight_mem_read_arbxbar_arbiters_next_15_13_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_243;
      weight_mem_read_arbxbar_arbiters_next_15_2_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_243;
      weight_mem_read_arbxbar_arbiters_next_15_12_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_243;
      weight_mem_read_arbxbar_arbiters_next_15_3_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_243;
      weight_mem_read_arbxbar_arbiters_next_15_11_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_243;
      weight_mem_read_arbxbar_arbiters_next_15_4_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_243;
      weight_mem_read_arbxbar_arbiters_next_15_10_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_243;
      weight_mem_read_arbxbar_arbiters_next_15_5_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_243;
      weight_mem_read_arbxbar_arbiters_next_15_9_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_243;
      weight_mem_read_arbxbar_arbiters_next_15_6_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_243;
      weight_mem_read_arbxbar_arbiters_next_15_8_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_243;
      weight_mem_read_arbxbar_arbiters_next_15_7_sva <= Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
          | Arbiter_16U_Roundrobin_pick_if_1_not_243;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      PECore_CheckStart_start_reg_sva <= 1'b0;
      PECore_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva
          <= 1'b0;
    end
    else if ( PECore_CheckStart_start_reg_and_cse ) begin
      PECore_CheckStart_start_reg_sva <= MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0,
          start_PopNB_mioi_idat_mxwt, PECore_DecodeAxiRead_switch_lp_and_3_rgt);
      PECore_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva
          <= MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0, start_PopNB_mioi_ivld_mxwt,
          PECore_DecodeAxiRead_switch_lp_and_3_rgt);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      PECore_RunBias_if_for_11_operator_4_false_slc_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_0_itm
          <= 1'b0;
      PECore_RunBias_if_for_10_operator_4_false_slc_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_0_itm
          <= 1'b0;
      PECore_RunBias_if_for_7_operator_4_false_slc_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_0_itm
          <= 1'b0;
      adpfloat_tmp_is_zero_land_7_lpi_1_dfm <= 1'b0;
      PECore_RunBias_if_for_6_operator_4_false_slc_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_0_itm
          <= 1'b0;
      adpfloat_tmp_is_zero_land_6_lpi_1_dfm <= 1'b0;
      PECore_RunBias_if_for_16_operator_32_true_slc_operator_32_true_acc_13_svs <=
          1'b0;
      PECore_RunBias_if_for_15_operator_32_true_slc_operator_32_true_acc_13_svs <=
          1'b0;
      PECore_RunBias_if_for_14_operator_32_true_slc_operator_32_true_acc_13_svs <=
          1'b0;
      PECore_RunBias_if_for_13_operator_32_true_slc_operator_32_true_acc_13_svs <=
          1'b0;
    end
    else if ( operator_4_false_and_cse ) begin
      PECore_RunBias_if_for_11_operator_4_false_slc_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_0_itm
          <= adpfloat_tmp_to_fixed_20U_14U_acc_sdt_11_sva_1[0];
      PECore_RunBias_if_for_10_operator_4_false_slc_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_0_itm
          <= adpfloat_tmp_to_fixed_20U_14U_acc_sdt_10_sva_1[0];
      PECore_RunBias_if_for_7_operator_4_false_slc_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_0_itm
          <= adpfloat_tmp_to_fixed_20U_14U_acc_sdt_7_sva_1[0];
      adpfloat_tmp_is_zero_land_7_lpi_1_dfm <= adpfloat_tmp_is_zero_land_7_lpi_1_dfm_mx1w0;
      PECore_RunBias_if_for_6_operator_4_false_slc_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_0_itm
          <= adpfloat_tmp_to_fixed_20U_14U_acc_sdt_6_sva_1[0];
      adpfloat_tmp_is_zero_land_6_lpi_1_dfm <= adpfloat_tmp_is_zero_land_6_lpi_1_dfm_mx1w0;
      PECore_RunBias_if_for_16_operator_32_true_slc_operator_32_true_acc_13_svs <=
          ~((input_mem_banks_write_if_for_if_mux_cse[38:32]!=7'b0000000));
      PECore_RunBias_if_for_15_operator_32_true_slc_operator_32_true_acc_13_svs <=
          ~((input_mem_banks_write_if_for_if_mux_cse[30:24]!=7'b0000000));
      PECore_RunBias_if_for_14_operator_32_true_slc_operator_32_true_acc_13_svs <=
          ~((input_mem_banks_write_if_for_if_mux_cse[22:16]!=7'b0000000));
      PECore_RunBias_if_for_13_operator_32_true_slc_operator_32_true_acc_13_svs <=
          ~((input_mem_banks_write_if_for_if_mux_cse[14:8]!=7'b0000000));
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      adpfloat_tmp_is_zero_land_11_lpi_1_dfm <= 1'b0;
      adpfloat_tmp_is_zero_land_10_lpi_1_dfm <= 1'b0;
    end
    else if ( adpfloat_tmp_is_zero_aelse_and_cse ) begin
      adpfloat_tmp_is_zero_land_11_lpi_1_dfm <= MUX_s_1_2_2(z_out_13_13, adpfloat_tmp_is_zero_land_11_lpi_1_dfm_mx1w0,
          operator_32_true_and_6_rgt);
      adpfloat_tmp_is_zero_land_10_lpi_1_dfm <= MUX_s_1_2_2(z_out_11_13, adpfloat_tmp_is_zero_land_10_lpi_1_dfm_mx1w0,
          operator_32_true_and_6_rgt);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_11_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~(PECore_RunBias_if_for_and_47_cse | PECore_RunBias_if_for_and_48_cse))
        ) begin
      PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_11_sva <= MUX_v_32_2_2(z_out_37,
          z_out_38, PECore_RunBias_if_for_and_50_rgt);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      PECore_RunBias_if_for_12_operator_32_true_slc_operator_32_true_acc_13_svs <=
          1'b0;
      PECore_RunBias_if_for_1_operator_32_true_slc_operator_32_true_acc_13_svs <=
          1'b0;
      PECore_RunBias_if_for_2_operator_32_true_slc_operator_32_true_acc_13_svs <=
          1'b0;
    end
    else if ( operator_32_true_and_12_cse ) begin
      PECore_RunBias_if_for_12_operator_32_true_slc_operator_32_true_acc_13_svs <=
          ~((input_mem_banks_write_if_for_if_mux_cse[94:88]!=7'b0000000));
      PECore_RunBias_if_for_1_operator_32_true_slc_operator_32_true_acc_13_svs <=
          ~((input_mem_banks_write_if_for_if_mux_cse[62:56]!=7'b0000000));
      PECore_RunBias_if_for_2_operator_32_true_slc_operator_32_true_acc_13_svs <=
          ~((input_mem_banks_write_if_for_if_mux_cse[70:64]!=7'b0000000));
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_10_0_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_10_1_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_10_2_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_10_3_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_10_4_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_10_5_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_10_6_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_10_7_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_10_8_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_10_9_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_10_10_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_10_11_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_10_12_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_10_13_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_10_14_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_10_15_sva_dfm <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_216_cse ) begin
      weight_port_read_out_data_10_0_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1;
      weight_port_read_out_data_10_1_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1;
      weight_port_read_out_data_10_2_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1;
      weight_port_read_out_data_10_3_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1;
      weight_port_read_out_data_10_4_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1;
      weight_port_read_out_data_10_5_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1;
      weight_port_read_out_data_10_6_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1;
      weight_port_read_out_data_10_7_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1;
      weight_port_read_out_data_10_8_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1;
      weight_port_read_out_data_10_9_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1;
      weight_port_read_out_data_10_10_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1;
      weight_port_read_out_data_10_11_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1;
      weight_port_read_out_data_10_12_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1;
      weight_port_read_out_data_10_13_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1;
      weight_port_read_out_data_10_14_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1;
      weight_port_read_out_data_10_15_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_9_0_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_9_1_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_9_2_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_9_3_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_9_4_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_9_5_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_9_6_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_9_7_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_9_8_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_9_9_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_9_10_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_9_11_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_9_12_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_9_13_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_9_14_sva_dfm <= 8'b00000000;
      weight_port_read_out_data_9_15_sva_dfm <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_232_cse ) begin
      weight_port_read_out_data_9_0_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44;
      weight_port_read_out_data_9_1_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42;
      weight_port_read_out_data_9_2_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40;
      weight_port_read_out_data_9_3_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
      weight_port_read_out_data_9_4_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
      weight_port_read_out_data_9_5_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
      weight_port_read_out_data_9_6_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
      weight_port_read_out_data_9_7_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
      weight_port_read_out_data_9_8_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
      weight_port_read_out_data_9_9_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
      weight_port_read_out_data_9_10_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
      weight_port_read_out_data_9_11_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
      weight_port_read_out_data_9_12_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
      weight_port_read_out_data_9_13_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
      weight_port_read_out_data_9_14_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16;
      weight_port_read_out_data_9_15_sva_dfm <= crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      adpfloat_tmp_is_zero_land_11_lpi_1_dfm_st <= 1'b0;
      adpfloat_tmp_is_zero_land_10_lpi_1_dfm_st <= 1'b0;
    end
    else if ( adpfloat_tmp_is_zero_aelse_and_4_cse ) begin
      adpfloat_tmp_is_zero_land_11_lpi_1_dfm_st <= MUX_s_1_2_2(z_out_12_13, adpfloat_tmp_is_zero_land_11_lpi_1_dfm_mx1w0,
          operator_32_true_and_2_rgt);
      adpfloat_tmp_is_zero_land_10_lpi_1_dfm_st <= MUX_s_1_2_2(z_out_10_13, adpfloat_tmp_is_zero_land_10_lpi_1_dfm_mx1w0,
          operator_32_true_and_2_rgt);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      accum_vector_data_9_sva <= 32'b00000000000000000000000000000000;
      accum_vector_data_6_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( accum_vector_data_and_15_cse ) begin
      accum_vector_data_9_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_2_cse;
      accum_vector_data_6_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_3_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      adpfloat_tmp_is_zero_land_7_lpi_1_dfm_st <= 1'b0;
      adpfloat_tmp_is_zero_land_6_lpi_1_dfm_st <= 1'b0;
    end
    else if ( adpfloat_tmp_is_zero_aelse_and_6_cse ) begin
      adpfloat_tmp_is_zero_land_7_lpi_1_dfm_st <= adpfloat_tmp_is_zero_land_7_lpi_1_dfm_mx1w0;
      adpfloat_tmp_is_zero_land_6_lpi_1_dfm_st <= adpfloat_tmp_is_zero_land_6_lpi_1_dfm_mx1w0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      accum_vector_data_5_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (PECore_UpdateFSM_switch_lp_equal_tmp_1 | input_mem_banks_load_store_for_else_and_cse)
        & while_stage_0_2 & (fsm_output[2]) ) begin
      accum_vector_data_5_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_4_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      PECore_RunBias_if_accum_vector_out_data_14_lpi_1_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~(or_dcpl_718 | (state_2_0_sva_0 & or_dcpl_370) |
        nor_499_cse)) ) begin
      PECore_RunBias_if_accum_vector_out_data_14_lpi_1_dfm <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_1_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      PECore_RunBias_if_accum_vector_out_data_15_lpi_1_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~ or_dcpl_718) & (fsm_output[2]) ) begin
      PECore_RunBias_if_accum_vector_out_data_15_lpi_1_dfm <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_1_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      PECore_RunMac_if_mux_160_itm <= 8'b00000000;
      PECore_RunMac_if_mux_161_itm <= 8'b00000000;
      PECore_RunMac_if_mux_162_itm <= 8'b00000000;
      PECore_RunMac_if_mux_163_itm <= 8'b00000000;
      PECore_RunMac_if_mux_164_itm <= 8'b00000000;
      PECore_RunMac_if_mux_165_itm <= 8'b00000000;
      PECore_RunMac_if_mux_166_itm <= 8'b00000000;
      PECore_RunMac_if_mux_167_itm <= 8'b00000000;
      PECore_RunMac_if_mux_168_itm <= 8'b00000000;
      PECore_RunMac_if_mux_169_itm <= 8'b00000000;
      PECore_RunMac_if_mux_170_itm <= 8'b00000000;
      PECore_RunMac_if_mux_171_itm <= 8'b00000000;
      PECore_RunMac_if_mux_172_itm <= 8'b00000000;
      PECore_RunMac_if_mux_173_itm <= 8'b00000000;
      PECore_RunMac_if_mux_174_itm <= 8'b00000000;
      PECore_RunMac_if_mux_175_itm <= 8'b00000000;
    end
    else if ( PECore_RunMac_if_and_685_cse ) begin
      PECore_RunMac_if_mux_160_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_for_mux_94_nl,
          weight_port_read_out_data_10_0_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_675_rgt , PECore_RunMac_if_and_676_rgt});
      PECore_RunMac_if_mux_161_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_for_mux_92_nl,
          weight_port_read_out_data_10_1_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_675_rgt , PECore_RunMac_if_and_676_rgt});
      PECore_RunMac_if_mux_162_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_for_mux_90_nl,
          weight_port_read_out_data_10_2_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_675_rgt , PECore_RunMac_if_and_676_rgt});
      PECore_RunMac_if_mux_163_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_for_mux_88_nl,
          weight_port_read_out_data_10_3_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_675_rgt , PECore_RunMac_if_and_676_rgt});
      PECore_RunMac_if_mux_164_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_for_mux_86_nl,
          weight_port_read_out_data_10_4_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_675_rgt , PECore_RunMac_if_and_676_rgt});
      PECore_RunMac_if_mux_165_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_for_mux_84_nl,
          weight_port_read_out_data_10_5_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_675_rgt , PECore_RunMac_if_and_676_rgt});
      PECore_RunMac_if_mux_166_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_for_mux_82_nl,
          weight_port_read_out_data_10_6_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_675_rgt , PECore_RunMac_if_and_676_rgt});
      PECore_RunMac_if_mux_167_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_for_mux_80_nl,
          weight_port_read_out_data_10_7_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_675_rgt , PECore_RunMac_if_and_676_rgt});
      PECore_RunMac_if_mux_168_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_for_mux_81_nl,
          weight_port_read_out_data_10_8_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_675_rgt , PECore_RunMac_if_and_676_rgt});
      PECore_RunMac_if_mux_169_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_for_mux_83_nl,
          weight_port_read_out_data_10_9_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_675_rgt , PECore_RunMac_if_and_676_rgt});
      PECore_RunMac_if_mux_170_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_for_mux_85_nl,
          weight_port_read_out_data_10_10_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_675_rgt , PECore_RunMac_if_and_676_rgt});
      PECore_RunMac_if_mux_171_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_for_mux_87_nl,
          weight_port_read_out_data_10_11_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_675_rgt , PECore_RunMac_if_and_676_rgt});
      PECore_RunMac_if_mux_172_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_for_mux_89_nl,
          weight_port_read_out_data_10_12_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_675_rgt , PECore_RunMac_if_and_676_rgt});
      PECore_RunMac_if_mux_173_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_for_mux_91_nl,
          weight_port_read_out_data_10_13_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_675_rgt , PECore_RunMac_if_and_676_rgt});
      PECore_RunMac_if_mux_174_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_for_mux_93_nl,
          weight_port_read_out_data_10_14_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_675_rgt , PECore_RunMac_if_and_676_rgt});
      PECore_RunMac_if_mux_175_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_for_mux_95_nl,
          weight_port_read_out_data_10_15_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_675_rgt , PECore_RunMac_if_and_676_rgt});
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      PECore_RunMac_if_mux_144_itm <= 8'b00000000;
      PECore_RunMac_if_mux_145_itm <= 8'b00000000;
      PECore_RunMac_if_mux_146_itm <= 8'b00000000;
      PECore_RunMac_if_mux_147_itm <= 8'b00000000;
      PECore_RunMac_if_mux_148_itm <= 8'b00000000;
      PECore_RunMac_if_mux_149_itm <= 8'b00000000;
      PECore_RunMac_if_mux_150_itm <= 8'b00000000;
      PECore_RunMac_if_mux_151_itm <= 8'b00000000;
      PECore_RunMac_if_mux_152_itm <= 8'b00000000;
      PECore_RunMac_if_mux_153_itm <= 8'b00000000;
      PECore_RunMac_if_mux_154_itm <= 8'b00000000;
      PECore_RunMac_if_mux_155_itm <= 8'b00000000;
      PECore_RunMac_if_mux_156_itm <= 8'b00000000;
      PECore_RunMac_if_mux_157_itm <= 8'b00000000;
      PECore_RunMac_if_mux_158_itm <= 8'b00000000;
      PECore_RunMac_if_mux_159_itm <= 8'b00000000;
    end
    else if ( PECore_RunMac_if_and_701_cse ) begin
      PECore_RunMac_if_mux_144_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_1_for_mux_78_nl,
          weight_port_read_out_data_9_0_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_627_rgt , PECore_RunMac_if_and_628_rgt});
      PECore_RunMac_if_mux_145_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_1_for_mux_76_nl,
          weight_port_read_out_data_9_1_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_627_rgt , PECore_RunMac_if_and_628_rgt});
      PECore_RunMac_if_mux_146_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_1_for_mux_74_nl,
          weight_port_read_out_data_9_2_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_627_rgt , PECore_RunMac_if_and_628_rgt});
      PECore_RunMac_if_mux_147_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_1_for_mux_72_nl,
          weight_port_read_out_data_9_3_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_627_rgt , PECore_RunMac_if_and_628_rgt});
      PECore_RunMac_if_mux_148_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_1_for_mux_70_nl,
          weight_port_read_out_data_9_4_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_627_rgt , PECore_RunMac_if_and_628_rgt});
      PECore_RunMac_if_mux_149_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_1_for_mux_68_nl,
          weight_port_read_out_data_9_5_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_627_rgt , PECore_RunMac_if_and_628_rgt});
      PECore_RunMac_if_mux_150_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_1_for_mux_66_nl,
          weight_port_read_out_data_9_6_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_627_rgt , PECore_RunMac_if_and_628_rgt});
      PECore_RunMac_if_mux_151_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_1_for_mux_64_nl,
          weight_port_read_out_data_9_7_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_627_rgt , PECore_RunMac_if_and_628_rgt});
      PECore_RunMac_if_mux_152_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_1_for_mux_65_nl,
          weight_port_read_out_data_9_8_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_627_rgt , PECore_RunMac_if_and_628_rgt});
      PECore_RunMac_if_mux_153_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_1_for_mux_67_nl,
          weight_port_read_out_data_9_9_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_627_rgt , PECore_RunMac_if_and_628_rgt});
      PECore_RunMac_if_mux_154_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_1_for_mux_69_nl,
          weight_port_read_out_data_9_10_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_627_rgt , PECore_RunMac_if_and_628_rgt});
      PECore_RunMac_if_mux_155_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_1_for_mux_71_nl,
          weight_port_read_out_data_9_11_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_627_rgt , PECore_RunMac_if_and_628_rgt});
      PECore_RunMac_if_mux_156_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_1_for_mux_73_nl,
          weight_port_read_out_data_9_12_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_627_rgt , PECore_RunMac_if_and_628_rgt});
      PECore_RunMac_if_mux_157_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_1_for_mux_75_nl,
          weight_port_read_out_data_9_13_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_627_rgt , PECore_RunMac_if_and_628_rgt});
      PECore_RunMac_if_mux_158_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_1_for_mux_77_nl,
          weight_port_read_out_data_9_14_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_627_rgt , PECore_RunMac_if_and_628_rgt});
      PECore_RunMac_if_mux_159_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_1_for_mux_79_nl,
          weight_port_read_out_data_9_15_sva_dfm, crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
          {PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_627_rgt , PECore_RunMac_if_and_628_rgt});
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      PECore_RunMac_if_mux_96_itm <= 8'b00000000;
      PECore_RunMac_if_mux_97_itm <= 8'b00000000;
      PECore_RunMac_if_mux_98_itm <= 8'b00000000;
      PECore_RunMac_if_mux_99_itm <= 8'b00000000;
      PECore_RunMac_if_mux_107_itm <= 8'b00000000;
      PECore_RunMac_if_mux_108_itm <= 8'b00000000;
      PECore_RunMac_if_mux_109_itm <= 8'b00000000;
      PECore_RunMac_if_mux_110_itm <= 8'b00000000;
      PECore_RunMac_if_mux_111_itm <= 8'b00000000;
      PECore_RunMac_if_mux_80_itm <= 8'b00000000;
      PECore_RunMac_if_mux_81_itm <= 8'b00000000;
      PECore_RunMac_if_mux_82_itm <= 8'b00000000;
      PECore_RunMac_if_mux_83_itm <= 8'b00000000;
      PECore_RunMac_if_mux_84_itm <= 8'b00000000;
      PECore_RunMac_if_mux_85_itm <= 8'b00000000;
      PECore_RunMac_if_mux_86_itm <= 8'b00000000;
      PECore_RunMac_if_mux_87_itm <= 8'b00000000;
      PECore_RunMac_if_mux_88_itm <= 8'b00000000;
      PECore_RunMac_if_mux_89_itm <= 8'b00000000;
      PECore_RunMac_if_mux_90_itm <= 8'b00000000;
      PECore_RunMac_if_mux_91_itm <= 8'b00000000;
      PECore_RunMac_if_mux_92_itm <= 8'b00000000;
      PECore_RunMac_if_mux_93_itm <= 8'b00000000;
      PECore_RunMac_if_mux_94_itm <= 8'b00000000;
      PECore_RunMac_if_mux_95_itm <= 8'b00000000;
    end
    else if ( PECore_RunMac_if_and_717_cse ) begin
      PECore_RunMac_if_mux_96_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_for_mux_62_nl,
          weight_port_read_out_data_6_0_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_97_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_for_mux_60_nl,
          weight_port_read_out_data_6_1_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_98_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_for_mux_58_nl,
          weight_port_read_out_data_6_2_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_99_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_for_mux_56_nl,
          weight_port_read_out_data_6_3_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_107_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_for_mux_55_nl,
          weight_port_read_out_data_6_11_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_108_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_for_mux_57_nl,
          weight_port_read_out_data_6_12_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_109_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_for_mux_59_nl,
          weight_port_read_out_data_6_13_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_110_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_for_mux_61_nl,
          weight_port_read_out_data_6_14_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_111_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_for_mux_63_nl,
          weight_port_read_out_data_6_15_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_80_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_1_for_mux_46_nl,
          weight_port_read_out_data_5_0_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_81_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_1_for_mux_44_nl,
          weight_port_read_out_data_5_1_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_82_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_1_for_mux_42_nl,
          weight_port_read_out_data_5_2_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_83_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_1_for_mux_40_nl,
          weight_port_read_out_data_5_3_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_84_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_1_for_mux_38_nl,
          weight_port_read_out_data_5_4_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_85_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_1_for_mux_36_nl,
          weight_port_read_out_data_5_5_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_86_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_1_for_mux_34_nl,
          weight_port_read_out_data_5_6_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_87_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_1_for_mux_32_nl,
          weight_port_read_out_data_5_7_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_88_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_1_for_mux_33_nl,
          weight_port_read_out_data_5_8_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_89_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_1_for_mux_35_nl,
          weight_port_read_out_data_5_9_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_90_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_1_for_mux_37_nl,
          weight_port_read_out_data_5_10_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_91_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_1_for_mux_39_nl,
          weight_port_read_out_data_5_11_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_92_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_1_for_mux_41_nl,
          weight_port_read_out_data_5_12_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_93_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_1_for_mux_43_nl,
          weight_port_read_out_data_5_13_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_94_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_1_for_mux_45_nl,
          weight_port_read_out_data_5_14_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
      PECore_RunMac_if_mux_95_itm <= MUX_v_8_2_2(PEManager_16U_ClusterLookup_1_for_mux_47_nl,
          weight_port_read_out_data_5_15_sva_dfm_mx1, PECore_RunMac_if_and_580_rgt);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_PECore_RunMac_if_mux_100_ftd <= 3'b000;
      reg_PECore_RunMac_if_mux_101_ftd <= 3'b000;
      reg_PECore_RunMac_if_mux_103_ftd <= 3'b000;
      reg_PECore_RunMac_if_mux_104_ftd <= 3'b000;
    end
    else if ( PECore_RunMac_if_and_721_ssc ) begin
      reg_PECore_RunMac_if_mux_100_ftd <= MUX_v_3_2_2(PEManager_16U_ClusterLookup_for_mux_54_nl,
          (weight_port_read_out_data_6_4_sva_dfm_mx1[7:5]), PECore_RunMac_if_and_570_rgt);
      reg_PECore_RunMac_if_mux_101_ftd <= MUX_v_3_2_2(PEManager_16U_ClusterLookup_for_mux_52_nl,
          (weight_port_read_out_data_6_5_sva_dfm_mx1[7:5]), PECore_RunMac_if_and_570_rgt);
      reg_PECore_RunMac_if_mux_103_ftd <= MUX_v_3_2_2(PEManager_16U_ClusterLookup_for_mux_48_nl,
          (weight_port_read_out_data_6_7_sva_dfm_mx1[7:5]), PECore_RunMac_if_and_570_rgt);
      reg_PECore_RunMac_if_mux_104_ftd <= MUX_v_3_2_2(PEManager_16U_ClusterLookup_for_mux_49_nl,
          (weight_port_read_out_data_6_8_sva_dfm_mx1[7:5]), PECore_RunMac_if_and_570_rgt);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_PECore_RunMac_if_mux_100_ftd_1 <= 5'b00000;
      reg_PECore_RunMac_if_mux_101_ftd_1 <= 5'b00000;
      reg_PECore_RunMac_if_mux_103_ftd_1 <= 5'b00000;
      reg_PECore_RunMac_if_mux_104_ftd_1 <= 5'b00000;
    end
    else if ( PECore_RunMac_if_and_867_cse ) begin
      reg_PECore_RunMac_if_mux_100_ftd_1 <= MUX1HOT_v_5_3_2(PECore_RunBias_if_for_10_operator_34_true_acc_nl,
          PEManager_16U_ClusterLookup_for_mux_139_nl, (weight_port_read_out_data_6_4_sva_dfm_mx1[4:0]),
          {PECore_RunMac_if_and_834_rgt , PECore_RunMac_if_and_569_rgt , PECore_RunMac_if_and_570_rgt});
      reg_PECore_RunMac_if_mux_101_ftd_1 <= MUX1HOT_v_5_3_2(PECore_RunBias_if_for_11_operator_34_true_acc_nl,
          PEManager_16U_ClusterLookup_for_mux_140_nl, (weight_port_read_out_data_6_5_sva_dfm_mx1[4:0]),
          {PECore_RunMac_if_and_834_rgt , PECore_RunMac_if_and_569_rgt , PECore_RunMac_if_and_570_rgt});
      reg_PECore_RunMac_if_mux_103_ftd_1 <= MUX1HOT_v_5_3_2(PECore_RunBias_if_for_6_operator_34_true_acc_nl,
          PEManager_16U_ClusterLookup_for_mux_142_nl, (weight_port_read_out_data_6_7_sva_dfm_mx1[4:0]),
          {PECore_RunMac_if_and_834_rgt , PECore_RunMac_if_and_569_rgt , PECore_RunMac_if_and_570_rgt});
      reg_PECore_RunMac_if_mux_104_ftd_1 <= MUX1HOT_v_5_3_2(PECore_RunBias_if_for_7_operator_34_true_acc_nl,
          PEManager_16U_ClusterLookup_for_mux_143_nl, (weight_port_read_out_data_6_8_sva_dfm_mx1[4:0]),
          {PECore_RunMac_if_and_834_rgt , PECore_RunMac_if_and_569_rgt , PECore_RunMac_if_and_570_rgt});
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_PECore_RunMac_if_mux_102_ftd <= 3'b000;
    end
    else if ( PECore_RunMac_if_and_723_ssc ) begin
      reg_PECore_RunMac_if_mux_102_ftd <= MUX_v_3_2_2(PEManager_16U_ClusterLookup_for_mux_50_nl,
          (weight_port_read_out_data_6_6_sva_dfm_mx1[7:5]), PECore_RunMac_if_and_570_rgt);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_PECore_RunMac_if_mux_102_ftd_1 <= 5'b00000;
    end
    else if ( PECore_RunMac_if_and_723_ssc & (~((fsm_output[3]) & PECore_RunMac_if_or_143_m1c))
        ) begin
      reg_PECore_RunMac_if_mux_102_ftd_1 <= MUX1HOT_v_5_3_2(PEManager_16U_ClusterLookup_for_mux_141_nl,
          (weight_port_read_out_data_6_6_sva_dfm_mx1[4:0]), PECore_RunBias_if_for_5_operator_34_true_acc_nl,
          {PECore_RunMac_if_and_569_rgt , PECore_RunMac_if_and_570_rgt , PECore_RunMac_if_and_829_nl});
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      PECore_RunMac_if_mux_105_itm <= 8'b00000000;
      PECore_RunMac_if_mux_106_itm <= 8'b00000000;
    end
    else if ( PECore_RunMac_if_and_726_cse ) begin
      PECore_RunMac_if_mux_105_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_for_mux_51_nl,
          weight_port_read_out_data_6_9_sva_dfm_mx1, ({3'b000 , PECore_RunBias_if_for_8_operator_34_true_acc_nl}),
          {PECore_RunMac_if_and_569_rgt , PECore_RunMac_if_and_570_rgt , PECore_RunMac_if_and_571_rgt});
      PECore_RunMac_if_mux_106_itm <= MUX1HOT_v_8_3_2(PEManager_16U_ClusterLookup_for_mux_53_nl,
          weight_port_read_out_data_6_10_sva_dfm_mx1, ({3'b000 , PECore_RunBias_if_for_9_operator_34_true_acc_nl}),
          {PECore_RunMac_if_and_569_rgt , PECore_RunMac_if_and_570_rgt , PECore_RunMac_if_and_571_rgt});
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & (fsm_output[2]) ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_1 <= and_5871_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      input_mem_banks_load_store_for_else_and_cse <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (fsm_output[1])) ) begin
      input_mem_banks_load_store_for_else_and_cse <= MUX_s_1_2_2(input_mem_banks_load_store_for_else_and_cse_1,
          while_and_30_itm_1, fsm_output[4]);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_and_2_itm <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_2_itm <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_and_5_itm <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_and_itm <= 1'b0;
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm <= 1'b0;
      w_axi_rsp_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_and_2_itm <= MUX_s_1_2_2(PECore_DecodeAxiRead_case_4_switch_lp_and_2_nl,
          pe_config_is_bias_sva, fsm_output[4]);
      PECore_DecodeAxiRead_switch_lp_nor_2_itm <= PECore_DecodeAxiRead_switch_lp_nor_2_itm_mx0w0;
      PECore_DecodeAxiRead_case_4_switch_lp_and_5_itm <= PECore_DecodeAxiRead_case_4_switch_lp_mux1h_13_nl
          & (~ PECore_DecodeAxiWrite_case_4_switch_lp_nor_tmp_1);
      PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm <= PECore_DecodeAxiRead_case_4_switch_lp_mux1h_11_nl
          & (~ PECore_DecodeAxiWrite_case_4_switch_lp_nor_tmp_1);
      PECore_DecodeAxiRead_case_4_switch_lp_and_itm <= PECore_DecodeAxiRead_case_4_switch_lp_mux1h_16_nl
          & (~ PECore_DecodeAxiWrite_case_4_switch_lp_nor_tmp_1);
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm <= ~(crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_tmp
          | (~ weight_read_ack_0_lpi_1_dfm_15_mx0));
      w_axi_rsp_lpi_1_dfm_1 <= ~((rva_in_PopNB_mio_mrgout_dat_sva_1[168]) | (~ rva_in_PopNB_mioi_ivld_mxwt)
          | is_start_sva);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~(PECore_RunBias_if_for_and_47_cse | PECore_RunBias_if_for_and_42_cse
        | PECore_DecodeAxiRead_switch_lp_and_3_rgt)) ) begin
      PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_1_sva <= MUX1HOT_v_32_3_2(z_out_38,
          z_out_40, z_out_39, {PECore_RunBias_if_for_and_49_nl , PECore_RunBias_if_for_and_45_rgt
          , PECore_DecodeAxiRead_switch_lp_and_2_cse});
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_4_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~((~(is_start_sva | (~((fsm_output[2:1]!=2'b00)))))
        | ((~ is_start_sva) & or_dcpl_251))) ) begin
      PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_4_sva <= MUX_v_32_2_2(z_out_39,
          z_out_40, PECore_RunBias_if_for_and_40_nl);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_5_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~(PECore_RunBias_if_for_and_cse | PECore_RunBias_if_for_and_48_cse
        | and_2966_cse)) ) begin
      PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_5_sva <= MUX1HOT_v_32_3_2(z_out_40,
          z_out_37, z_out_39, {PECore_RunBias_if_for_and_34_rgt , PECore_RunBias_if_for_and_50_rgt
          , PECore_RunBias_if_for_and_36_nl});
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_reg_data_asn_1_itm <= 20'b00000000000000000000;
    end
    else if ( act_port_reg_data_and_enex5 ) begin
      act_port_reg_data_asn_1_itm <= act_port_reg_data_14_sva;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_reg_data_asn_2_itm <= 20'b00000000000000000000;
    end
    else if ( act_port_reg_data_and_28_enex5 ) begin
      act_port_reg_data_asn_2_itm <= act_port_reg_data_13_sva;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_reg_data_asn_3_itm <= 20'b00000000000000000000;
    end
    else if ( act_port_reg_data_and_29_enex5 ) begin
      act_port_reg_data_asn_3_itm <= act_port_reg_data_12_sva;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_reg_data_asn_itm <= 20'b00000000000000000000;
    end
    else if ( act_port_reg_data_and_30_enex5 ) begin
      act_port_reg_data_asn_itm <= act_port_reg_data_15_sva;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_nor_tmp <= 1'b0;
    end
    else if ( PECoreRun_wen & (is_start_sva | (~ (fsm_output[2]))) ) begin
      PECore_DecodeAxiRead_switch_lp_nor_tmp <= MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_nor_tmp_mx0w0,
          adpfloat_tmp_is_zero_if_adpfloat_tmp_is_zero_if_nor_nl, fsm_output[2]);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_out_reg_data_103_96_sva_dfm_4 <= 8'b00000000;
      rva_out_reg_data_111_104_sva_dfm_4 <= 8'b00000000;
      rva_out_reg_data_119_112_sva_dfm_4 <= 8'b00000000;
      rva_out_reg_data_127_120_sva_dfm_4 <= 8'b00000000;
      rva_out_reg_data_87_80_sva_dfm_4 <= 8'b00000000;
      rva_out_reg_data_95_88_sva_dfm_4 <= 8'b00000000;
      rva_out_reg_data_71_64_sva_dfm_4 <= 8'b00000000;
      rva_out_reg_data_79_72_sva_dfm_4 <= 8'b00000000;
      rva_out_reg_data_55_48_sva_dfm_4 <= 8'b00000000;
      rva_out_reg_data_63_56_sva_dfm_4 <= 8'b00000000;
      rva_out_reg_data_47_40_sva_dfm_4 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_91_cse ) begin
      rva_out_reg_data_103_96_sva_dfm_4 <= MUX1HOT_v_8_5_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_29_nl,
          (input_mem_banks_bank_array_impl_data0_rsci_q_d[103:96]), crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18,
          PEManager_16U_ClusterLookup_1_for_mux_62_nl, weight_port_read_out_data_7_0_sva_dfm_mx1,
          {(~ (fsm_output[2])) , rva_out_reg_data_and_87_rgt , rva_out_reg_data_and_88_rgt
          , PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_580_rgt});
      rva_out_reg_data_111_104_sva_dfm_4 <= MUX1HOT_v_8_5_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_28_nl,
          (input_mem_banks_bank_array_impl_data0_rsci_q_d[111:104]), crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20,
          PEManager_16U_ClusterLookup_1_for_mux_60_nl, weight_port_read_out_data_7_1_sva_dfm_mx1,
          {(~ (fsm_output[2])) , rva_out_reg_data_and_87_rgt , rva_out_reg_data_and_88_rgt
          , PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_580_rgt});
      rva_out_reg_data_119_112_sva_dfm_4 <= MUX1HOT_v_8_5_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_27_nl,
          (input_mem_banks_bank_array_impl_data0_rsci_q_d[119:112]), crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22,
          PEManager_16U_ClusterLookup_1_for_mux_58_nl, weight_port_read_out_data_7_2_sva_dfm_mx1,
          {(~ (fsm_output[2])) , rva_out_reg_data_and_87_rgt , rva_out_reg_data_and_88_rgt
          , PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_580_rgt});
      rva_out_reg_data_127_120_sva_dfm_4 <= MUX1HOT_v_8_5_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_26_nl,
          (input_mem_banks_bank_array_impl_data0_rsci_q_d[127:120]), crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_2,
          PEManager_16U_ClusterLookup_1_for_mux_56_nl, weight_port_read_out_data_7_3_sva_dfm_mx1,
          {(~ (fsm_output[2])) , rva_out_reg_data_and_87_rgt , rva_out_reg_data_and_88_rgt
          , PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_580_rgt});
      rva_out_reg_data_87_80_sva_dfm_4 <= MUX1HOT_v_8_5_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_25_nl,
          (input_mem_banks_bank_array_impl_data0_rsci_q_d[87:80]), crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24,
          PEManager_16U_ClusterLookup_1_for_mux_49_nl, weight_port_read_out_data_7_8_sva_dfm_mx1,
          {(~ (fsm_output[2])) , rva_out_reg_data_and_87_rgt , rva_out_reg_data_and_88_rgt
          , PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_580_rgt});
      rva_out_reg_data_95_88_sva_dfm_4 <= MUX1HOT_v_8_5_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl,
          (input_mem_banks_bank_array_impl_data0_rsci_q_d[95:88]), crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26,
          PEManager_16U_ClusterLookup_1_for_mux_51_nl, weight_port_read_out_data_7_9_sva_dfm_mx1,
          {(~ (fsm_output[2])) , rva_out_reg_data_and_87_rgt , rva_out_reg_data_and_88_rgt
          , PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_580_rgt});
      rva_out_reg_data_71_64_sva_dfm_4 <= MUX1HOT_v_8_5_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl,
          (input_mem_banks_bank_array_impl_data0_rsci_q_d[71:64]), crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28,
          PEManager_16U_ClusterLookup_1_for_mux_48_nl, weight_port_read_out_data_7_7_sva_dfm_mx1,
          {(~ (fsm_output[2])) , rva_out_reg_data_and_87_rgt , rva_out_reg_data_and_88_rgt
          , PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_580_rgt});
      rva_out_reg_data_79_72_sva_dfm_4 <= MUX1HOT_v_8_5_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl,
          (input_mem_banks_bank_array_impl_data0_rsci_q_d[79:72]), crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30,
          PEManager_16U_ClusterLookup_for_mux_4_nl, weight_port_read_out_data_0_12_sva_dfm_mx1,
          {(~ (fsm_output[2])) , rva_out_reg_data_and_87_rgt , rva_out_reg_data_and_88_rgt
          , PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_580_rgt});
      rva_out_reg_data_55_48_sva_dfm_4 <= MUX1HOT_v_8_5_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl,
          (input_mem_banks_bank_array_impl_data0_rsci_q_d[55:48]), crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32,
          PEManager_16U_ClusterLookup_1_for_mux_52_nl, weight_port_read_out_data_7_5_sva_dfm_mx1,
          {(~ (fsm_output[2])) , rva_out_reg_data_and_87_rgt , rva_out_reg_data_and_88_rgt
          , PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_580_rgt});
      rva_out_reg_data_63_56_sva_dfm_4 <= MUX1HOT_v_8_5_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_20_nl,
          (input_mem_banks_bank_array_impl_data0_rsci_q_d[63:56]), crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34,
          PEManager_16U_ClusterLookup_1_for_mux_50_nl, weight_port_read_out_data_7_6_sva_dfm_mx1,
          {(~ (fsm_output[2])) , rva_out_reg_data_and_87_rgt , rva_out_reg_data_and_88_rgt
          , PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_580_rgt});
      rva_out_reg_data_47_40_sva_dfm_4 <= MUX1HOT_v_8_5_2(PECore_DecodeAxiRead_case_4_switch_lp_and_3_nl,
          (input_mem_banks_bank_array_impl_data0_rsci_q_d[47:40]), crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36,
          PEManager_16U_ClusterLookup_1_for_mux_54_nl, weight_port_read_out_data_7_4_sva_dfm_mx1,
          {(~ (fsm_output[2])) , rva_out_reg_data_and_87_rgt , rva_out_reg_data_and_88_rgt
          , PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_580_rgt});
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_1_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]))
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_1_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= weight_mem_read_arbxbar_xbar_for_3_1_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_2_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]))
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_2_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= weight_mem_read_arbxbar_xbar_for_3_2_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_3_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]))
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_3_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= weight_mem_read_arbxbar_xbar_for_3_3_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_4_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]))
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_4_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= weight_mem_read_arbxbar_xbar_for_3_4_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_5_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]))
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_5_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= weight_mem_read_arbxbar_xbar_for_3_5_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_6_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]))
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_6_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= weight_mem_read_arbxbar_xbar_for_3_6_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_7_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]))
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_7_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= weight_mem_read_arbxbar_xbar_for_3_7_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_8_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]))
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_8_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= weight_mem_read_arbxbar_xbar_for_3_8_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_9_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8]))
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_9_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= weight_mem_read_arbxbar_xbar_for_3_9_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_10_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[9]))
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_10_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= weight_mem_read_arbxbar_xbar_for_3_10_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_11_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[10]))
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_11_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= weight_mem_read_arbxbar_xbar_for_3_11_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_12_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11]))
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_12_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= weight_mem_read_arbxbar_xbar_for_3_12_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_13_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12]))
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_13_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= weight_mem_read_arbxbar_xbar_for_3_13_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_14_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13]))
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_14_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= weight_mem_read_arbxbar_xbar_for_3_14_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_15_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14]))
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_15_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= weight_mem_read_arbxbar_xbar_for_3_15_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_for_3_16_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]))
        ) begin
      weight_mem_read_arbxbar_xbar_for_3_16_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva
          <= weight_mem_read_arbxbar_xbar_for_3_16_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_pe_config_UpdateInputCounter_if_nor_svs
          <= 1'b0;
      PECore_UpdateFSM_case_4_is_output_end_pe_config_UpdateManagerCounter_nand_itm
          <= 1'b0;
      PECore_UpdateFSM_switch_lp_unequal_tmp <= 1'b0;
      PECore_RunMac_nor_tmp <= 1'b0;
    end
    else if ( pe_config_UpdateInputCounter_if_and_cse ) begin
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_pe_config_UpdateInputCounter_if_nor_svs
          <= pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_pe_config_UpdateInputCounter_if_nor_svs_1;
      PECore_UpdateFSM_case_4_is_output_end_pe_config_UpdateManagerCounter_nand_itm
          <= ~(pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1
          & pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_nor_svs_1);
      PECore_UpdateFSM_switch_lp_unequal_tmp <= PECore_UpdateFSM_switch_lp_unequal_tmp_1;
      PECore_RunMac_nor_tmp <= MUX_s_1_2_2(PECore_RunMac_nor_nl, PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl,
          state_2_0_sva_0);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_PECore_RunMac_if_mux_1_ftd_1 <= 5'b00000;
      reg_PECore_RunMac_if_mux_10_ftd_1 <= 5'b00000;
      PECore_RunMac_if_mux_64_itm <= 8'b00000000;
      PECore_RunMac_if_mux_65_itm <= 8'b00000000;
      PECore_RunMac_if_mux_66_itm <= 8'b00000000;
      PECore_RunMac_if_mux_67_itm <= 8'b00000000;
      PECore_RunMac_if_mux_68_itm <= 8'b00000000;
      PECore_RunMac_if_mux_69_itm <= 8'b00000000;
      PECore_RunMac_if_mux_70_itm <= 8'b00000000;
      PECore_RunMac_if_mux_71_itm <= 8'b00000000;
      PECore_RunMac_if_mux_72_itm <= 8'b00000000;
      PECore_RunMac_if_mux_73_itm <= 8'b00000000;
      PECore_RunMac_if_mux_74_itm <= 8'b00000000;
      PECore_RunMac_if_mux_75_itm <= 8'b00000000;
      PECore_RunMac_if_mux_76_itm <= 8'b00000000;
      PECore_RunMac_if_mux_77_itm <= 8'b00000000;
      PECore_RunMac_if_mux_78_itm <= 8'b00000000;
      PECore_RunMac_if_mux_79_itm <= 8'b00000000;
      PECore_RunMac_if_mux_48_itm <= 8'b00000000;
      PECore_RunMac_if_mux_49_itm <= 8'b00000000;
      PECore_RunMac_if_mux_50_itm <= 8'b00000000;
      PECore_RunMac_if_mux_51_itm <= 8'b00000000;
      PECore_RunMac_if_mux_52_itm <= 8'b00000000;
      PECore_RunMac_if_mux_53_itm <= 8'b00000000;
      PECore_RunMac_if_mux_54_itm <= 8'b00000000;
      PECore_RunMac_if_mux_55_itm <= 8'b00000000;
      PECore_RunMac_if_mux_56_itm <= 8'b00000000;
      PECore_RunMac_if_mux_57_itm <= 8'b00000000;
      PECore_RunMac_if_mux_58_itm <= 8'b00000000;
      PECore_RunMac_if_mux_59_itm <= 8'b00000000;
      PECore_RunMac_if_mux_60_itm <= 8'b00000000;
      PECore_RunMac_if_mux_61_itm <= 8'b00000000;
      PECore_RunMac_if_mux_62_itm <= 8'b00000000;
      PECore_RunMac_if_mux_63_itm <= 8'b00000000;
      PECore_RunMac_if_mux_32_itm <= 8'b00000000;
      PECore_RunMac_if_mux_33_itm <= 8'b00000000;
      PECore_RunMac_if_mux_34_itm <= 8'b00000000;
      PECore_RunMac_if_mux_35_itm <= 8'b00000000;
      PECore_RunMac_if_mux_36_itm <= 8'b00000000;
      PECore_RunMac_if_mux_37_itm <= 8'b00000000;
      PECore_RunMac_if_mux_38_itm <= 8'b00000000;
      PECore_RunMac_if_mux_39_itm <= 8'b00000000;
      PECore_RunMac_if_mux_40_itm <= 8'b00000000;
      PECore_RunMac_if_mux_41_itm <= 8'b00000000;
      PECore_RunMac_if_mux_42_itm <= 8'b00000000;
      PECore_RunMac_if_mux_43_itm <= 8'b00000000;
      PECore_RunMac_if_mux_44_itm <= 8'b00000000;
      PECore_RunMac_if_mux_45_itm <= 8'b00000000;
      PECore_RunMac_if_mux_46_itm <= 8'b00000000;
      PECore_RunMac_if_mux_47_itm <= 8'b00000000;
      reg_PECore_RunMac_if_mux_124_ftd_1 <= 4'b0000;
      reg_PECore_RunMac_if_mux_125_ftd_1 <= 4'b0000;
      reg_PECore_RunMac_if_mux_126_ftd_1 <= 4'b0000;
      reg_PECore_RunMac_if_mux_127_ftd_1 <= 4'b0000;
    end
    else if ( PECore_RunMac_if_and_872_cse ) begin
      reg_PECore_RunMac_if_mux_1_ftd_1 <= MUX1HOT_v_5_5_2(({2'b00 , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_3_1_lpi_1_dfm_1}),
          PEManager_16U_ClusterLookup_for_mux_145_nl, (weight_port_read_out_data_0_1_sva_dfm_mx1[4:0]),
          (crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_12_mx1w2[4:0]),
          PECore_RunBias_if_for_3_operator_34_true_acc_nl, {(fsm_output[1]) , PECore_RunMac_if_and_569_rgt
          , PECore_RunMac_if_and_570_rgt , PECore_RunBias_if_for_and_42_cse , PECore_RunMac_if_and_820_rgt});
      reg_PECore_RunMac_if_mux_10_ftd_1 <= MUX1HOT_v_5_5_2(({3'b000 , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_13_1_0_lpi_1_dfm_1}),
          PEManager_16U_ClusterLookup_for_mux_144_nl, (weight_port_read_out_data_0_10_sva_dfm_mx1[4:0]),
          (crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_11_mx1w2[4:0]),
          PECore_RunBias_if_for_4_operator_34_true_acc_nl, {(fsm_output[1]) , PECore_RunMac_if_and_569_rgt
          , PECore_RunMac_if_and_570_rgt , PECore_RunBias_if_for_and_42_cse , PECore_RunMac_if_and_820_rgt});
      PECore_RunMac_if_mux_64_itm <= MUX_v_8_2_2(weight_port_read_out_data_4_0_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_46_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_65_itm <= MUX_v_8_2_2(weight_port_read_out_data_4_1_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_44_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_66_itm <= MUX_v_8_2_2(weight_port_read_out_data_4_2_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_42_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_67_itm <= MUX_v_8_2_2(weight_port_read_out_data_4_3_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_40_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_68_itm <= MUX_v_8_2_2(weight_port_read_out_data_4_4_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_38_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_69_itm <= MUX_v_8_2_2(weight_port_read_out_data_4_5_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_36_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_70_itm <= MUX_v_8_2_2(weight_port_read_out_data_4_6_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_34_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_71_itm <= MUX_v_8_2_2(weight_port_read_out_data_4_7_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_32_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_72_itm <= MUX_v_8_2_2(weight_port_read_out_data_4_8_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_33_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_73_itm <= MUX_v_8_2_2(weight_port_read_out_data_4_9_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_35_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_74_itm <= MUX_v_8_2_2(weight_port_read_out_data_4_10_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_37_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_75_itm <= MUX_v_8_2_2(weight_port_read_out_data_4_11_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_39_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_76_itm <= MUX_v_8_2_2(weight_port_read_out_data_4_12_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_41_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_77_itm <= MUX_v_8_2_2(weight_port_read_out_data_4_13_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_43_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_78_itm <= MUX_v_8_2_2(weight_port_read_out_data_4_14_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_45_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_79_itm <= MUX_v_8_2_2(weight_port_read_out_data_4_15_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_47_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_48_itm <= MUX_v_8_2_2(weight_port_read_out_data_3_0_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_30_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_49_itm <= MUX_v_8_2_2(weight_port_read_out_data_3_1_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_28_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_50_itm <= MUX_v_8_2_2(weight_port_read_out_data_3_2_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_26_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_51_itm <= MUX_v_8_2_2(weight_port_read_out_data_3_3_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_24_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_52_itm <= MUX_v_8_2_2(weight_port_read_out_data_3_4_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_22_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_53_itm <= MUX_v_8_2_2(weight_port_read_out_data_3_5_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_20_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_54_itm <= MUX_v_8_2_2(weight_port_read_out_data_3_6_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_18_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_55_itm <= MUX_v_8_2_2(weight_port_read_out_data_3_7_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_16_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_56_itm <= MUX_v_8_2_2(weight_port_read_out_data_3_8_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_17_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_57_itm <= MUX_v_8_2_2(weight_port_read_out_data_3_9_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_19_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_58_itm <= MUX_v_8_2_2(weight_port_read_out_data_3_10_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_21_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_59_itm <= MUX_v_8_2_2(weight_port_read_out_data_3_11_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_23_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_60_itm <= MUX_v_8_2_2(weight_port_read_out_data_3_12_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_25_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_61_itm <= MUX_v_8_2_2(weight_port_read_out_data_3_13_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_27_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_62_itm <= MUX_v_8_2_2(weight_port_read_out_data_3_14_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_29_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_63_itm <= MUX_v_8_2_2(weight_port_read_out_data_3_15_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_31_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_32_itm <= MUX_v_8_2_2(weight_port_read_out_data_2_0_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_30_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_33_itm <= MUX_v_8_2_2(weight_port_read_out_data_2_1_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_28_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_34_itm <= MUX_v_8_2_2(weight_port_read_out_data_2_2_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_26_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_35_itm <= MUX_v_8_2_2(weight_port_read_out_data_2_3_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_24_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_36_itm <= MUX_v_8_2_2(weight_port_read_out_data_2_4_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_22_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_37_itm <= MUX_v_8_2_2(weight_port_read_out_data_2_5_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_20_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_38_itm <= MUX_v_8_2_2(weight_port_read_out_data_2_6_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_18_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_39_itm <= MUX_v_8_2_2(weight_port_read_out_data_2_7_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_16_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_40_itm <= MUX_v_8_2_2(weight_port_read_out_data_2_8_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_17_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_41_itm <= MUX_v_8_2_2(weight_port_read_out_data_2_9_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_19_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_42_itm <= MUX_v_8_2_2(weight_port_read_out_data_2_10_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_21_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_43_itm <= MUX_v_8_2_2(weight_port_read_out_data_2_11_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_23_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_44_itm <= MUX_v_8_2_2(weight_port_read_out_data_2_12_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_25_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_45_itm <= MUX_v_8_2_2(weight_port_read_out_data_2_13_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_27_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_46_itm <= MUX_v_8_2_2(weight_port_read_out_data_2_14_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_29_nl, PECore_RunMac_if_and_346_rgt);
      PECore_RunMac_if_mux_47_itm <= MUX_v_8_2_2(weight_port_read_out_data_2_15_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_31_nl, PECore_RunMac_if_and_346_rgt);
      reg_PECore_RunMac_if_mux_124_ftd_1 <= MUX1HOT_v_4_4_2(crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_12_lpi_1_dfm_1,
          adpfloat_tmp_to_fixed_20U_14U_acc_sdt_2_sva_mx0w1, PEManager_16U_ClusterLookup_1_for_mux_131_nl,
          (weight_port_read_out_data_7_12_sva_dfm_mx1[3:0]), {(fsm_output[1]) , PECore_RunMac_if_and_571_rgt
          , PECore_RunMac_if_and_472_rgt , PECore_RunMac_if_and_470_cse});
      reg_PECore_RunMac_if_mux_125_ftd_1 <= MUX1HOT_v_4_4_2(crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_14_lpi_1_dfm_1,
          adpfloat_tmp_to_fixed_20U_14U_acc_sdt_3_sva_mx0w1, PEManager_16U_ClusterLookup_1_for_mux_130_nl,
          (weight_port_read_out_data_7_13_sva_dfm_mx1[3:0]), {(fsm_output[1]) , PECore_RunMac_if_and_571_rgt
          , PECore_RunMac_if_and_472_rgt , PECore_RunMac_if_and_470_cse});
      reg_PECore_RunMac_if_mux_126_ftd_1 <= MUX1HOT_v_4_4_2(({crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_15_lpi_1_dfm_1_3_1
          , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_15_lpi_1_dfm_1_0}),
          adpfloat_tmp_to_fixed_20U_14U_acc_sdt_4_sva_mx0w1, PEManager_16U_ClusterLookup_1_for_mux_129_nl,
          (weight_port_read_out_data_7_14_sva_dfm_mx1[3:0]), {(fsm_output[1]) , PECore_RunMac_if_and_571_rgt
          , PECore_RunMac_if_and_472_rgt , PECore_RunMac_if_and_470_cse});
      reg_PECore_RunMac_if_mux_127_ftd_1 <= MUX1HOT_v_4_4_2(crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_2_lpi_1_dfm_1,
          adpfloat_tmp_to_fixed_20U_14U_acc_sdt_5_sva_mx0w1, PEManager_16U_ClusterLookup_1_for_mux_128_nl,
          (weight_port_read_out_data_7_15_sva_dfm_mx1[3:0]), {(fsm_output[1]) , PECore_RunMac_if_and_571_rgt
          , PECore_RunMac_if_and_472_rgt , PECore_RunMac_if_and_470_cse});
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      PECore_RunMac_if_mux_176_itm <= 8'b00000000;
      PECore_RunMac_if_mux_177_itm <= 8'b00000000;
      PECore_RunMac_if_mux_178_itm <= 8'b00000000;
      PECore_RunMac_if_mux_179_itm <= 8'b00000000;
      PECore_RunMac_if_mux_180_itm <= 8'b00000000;
      PECore_RunMac_if_mux_181_itm <= 8'b00000000;
      PECore_RunMac_if_mux_182_itm <= 8'b00000000;
      PECore_RunMac_if_mux_183_itm <= 8'b00000000;
      PECore_RunMac_if_mux_184_itm <= 8'b00000000;
      PECore_RunMac_if_mux_185_itm <= 8'b00000000;
      PECore_RunMac_if_mux_186_itm <= 8'b00000000;
      PECore_RunMac_if_mux_187_itm <= 8'b00000000;
      PECore_RunMac_if_mux_188_itm <= 8'b00000000;
      PECore_RunMac_if_mux_189_itm <= 8'b00000000;
      PECore_RunMac_if_mux_190_itm <= 8'b00000000;
      PECore_RunMac_if_mux_191_itm <= 8'b00000000;
      PECore_RunMac_if_mux_16_itm <= 8'b00000000;
      PECore_RunMac_if_mux_17_itm <= 8'b00000000;
      PECore_RunMac_if_mux_18_itm <= 8'b00000000;
      PECore_RunMac_if_mux_19_itm <= 8'b00000000;
      PECore_RunMac_if_mux_20_itm <= 8'b00000000;
      PECore_RunMac_if_mux_21_itm <= 8'b00000000;
      PECore_RunMac_if_mux_22_itm <= 8'b00000000;
      PECore_RunMac_if_mux_23_itm <= 8'b00000000;
      PECore_RunMac_if_mux_24_itm <= 8'b00000000;
      PECore_RunMac_if_mux_25_itm <= 8'b00000000;
      PECore_RunMac_if_mux_26_itm <= 8'b00000000;
      PECore_RunMac_if_mux_27_itm <= 8'b00000000;
      PECore_RunMac_if_mux_28_itm <= 8'b00000000;
      PECore_RunMac_if_mux_29_itm <= 8'b00000000;
      PECore_RunMac_if_mux_30_itm <= 8'b00000000;
      PECore_RunMac_if_mux_31_itm <= 8'b00000000;
      PECore_RunMac_if_mux_itm <= 8'b00000000;
      PECore_RunMac_if_mux_2_itm <= 8'b00000000;
      PECore_RunMac_if_mux_3_itm <= 8'b00000000;
      PECore_RunMac_if_mux_4_itm <= 8'b00000000;
      PECore_RunMac_if_mux_5_itm <= 8'b00000000;
      PECore_RunMac_if_mux_6_itm <= 8'b00000000;
      PECore_RunMac_if_mux_7_itm <= 8'b00000000;
      PECore_RunMac_if_mux_8_itm <= 8'b00000000;
      PECore_RunMac_if_mux_9_itm <= 8'b00000000;
      PECore_RunMac_if_mux_15_itm <= 8'b00000000;
    end
    else if ( PECore_RunMac_if_and_cse ) begin
      PECore_RunMac_if_mux_176_itm <= MUX_v_8_2_2(weight_mem_run_1_for_5_mux_30_nl,
          PEManager_16U_ClusterLookup_1_for_mux_94_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_177_itm <= MUX_v_8_2_2(weight_mem_run_1_for_5_mux_31_nl,
          PEManager_16U_ClusterLookup_1_for_mux_92_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_178_itm <= MUX_v_8_2_2(weight_mem_run_1_for_5_mux_32_nl,
          PEManager_16U_ClusterLookup_1_for_mux_90_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_179_itm <= MUX_v_8_2_2(weight_mem_run_1_for_5_mux_33_nl,
          PEManager_16U_ClusterLookup_1_for_mux_88_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_180_itm <= MUX_v_8_2_2(weight_mem_run_1_for_5_mux_34_nl,
          PEManager_16U_ClusterLookup_1_for_mux_86_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_181_itm <= MUX_v_8_2_2(weight_mem_run_1_for_5_mux_35_nl,
          PEManager_16U_ClusterLookup_1_for_mux_84_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_182_itm <= MUX_v_8_2_2(weight_mem_run_1_for_5_mux_36_nl,
          PEManager_16U_ClusterLookup_1_for_mux_82_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_183_itm <= MUX_v_8_2_2(weight_mem_run_1_for_5_mux_37_nl,
          PEManager_16U_ClusterLookup_1_for_mux_80_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_184_itm <= MUX_v_8_2_2(weight_mem_run_1_for_5_mux_38_nl,
          PEManager_16U_ClusterLookup_1_for_mux_81_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_185_itm <= MUX_v_8_2_2(weight_mem_run_1_for_5_mux_39_nl,
          PEManager_16U_ClusterLookup_1_for_mux_83_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_186_itm <= MUX_v_8_2_2(weight_mem_run_1_for_5_mux_40_nl,
          PEManager_16U_ClusterLookup_1_for_mux_85_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_187_itm <= MUX_v_8_2_2(weight_mem_run_1_for_5_mux_41_nl,
          PEManager_16U_ClusterLookup_1_for_mux_87_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_188_itm <= MUX_v_8_2_2(weight_mem_run_1_for_5_mux_42_nl,
          PEManager_16U_ClusterLookup_1_for_mux_89_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_189_itm <= MUX_v_8_2_2(weight_mem_run_1_for_5_mux_43_nl,
          PEManager_16U_ClusterLookup_1_for_mux_91_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_190_itm <= MUX_v_8_2_2(weight_mem_run_1_for_5_mux_44_nl,
          PEManager_16U_ClusterLookup_1_for_mux_93_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_191_itm <= MUX_v_8_2_2(data_in_tmp_operator_for_mux_34_nl,
          PEManager_16U_ClusterLookup_1_for_mux_95_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_16_itm <= MUX_v_8_2_2(weight_port_read_out_data_1_0_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_17_itm <= MUX_v_8_2_2(weight_port_read_out_data_1_1_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_1_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_18_itm <= MUX_v_8_2_2(weight_port_read_out_data_1_2_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_2_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_19_itm <= MUX_v_8_2_2(weight_port_read_out_data_1_3_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_3_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_20_itm <= MUX_v_8_2_2(weight_port_read_out_data_1_4_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_4_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_21_itm <= MUX_v_8_2_2(weight_port_read_out_data_1_5_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_5_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_22_itm <= MUX_v_8_2_2(weight_port_read_out_data_1_6_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_6_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_23_itm <= MUX_v_8_2_2(weight_port_read_out_data_1_7_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_7_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_24_itm <= MUX_v_8_2_2(weight_port_read_out_data_1_8_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_8_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_25_itm <= MUX_v_8_2_2(weight_port_read_out_data_1_9_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_9_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_26_itm <= MUX_v_8_2_2(weight_port_read_out_data_1_10_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_10_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_27_itm <= MUX_v_8_2_2(weight_port_read_out_data_1_11_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_11_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_28_itm <= MUX_v_8_2_2(weight_port_read_out_data_1_12_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_12_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_29_itm <= MUX_v_8_2_2(weight_port_read_out_data_1_13_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_13_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_30_itm <= MUX_v_8_2_2(weight_port_read_out_data_1_14_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_14_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_31_itm <= MUX_v_8_2_2(weight_port_read_out_data_1_15_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_1_for_mux_15_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_itm <= MUX_v_8_2_2(weight_port_read_out_data_0_0_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_2_itm <= MUX_v_8_2_2(weight_port_read_out_data_0_2_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_14_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_3_itm <= MUX_v_8_2_2(weight_port_read_out_data_0_3_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_13_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_4_itm <= MUX_v_8_2_2(weight_port_read_out_data_0_4_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_12_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_5_itm <= MUX_v_8_2_2(weight_port_read_out_data_0_5_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_11_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_6_itm <= MUX_v_8_2_2(weight_port_read_out_data_0_6_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_10_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_7_itm <= MUX_v_8_2_2(weight_port_read_out_data_0_7_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_9_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_8_itm <= MUX_v_8_2_2(weight_port_read_out_data_0_8_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_8_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_9_itm <= MUX_v_8_2_2(weight_port_read_out_data_0_9_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_7_nl, pe_config_is_cluster_sva);
      PECore_RunMac_if_mux_15_itm <= MUX_v_8_2_2(weight_port_read_out_data_0_15_sva_dfm_mx1,
          PEManager_16U_ClusterLookup_for_mux_1_nl, pe_config_is_cluster_sva);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_PECore_RunBias_if_accum_vector_out_data_6_lpi_1_dfm_ftd_12 <= 20'b00000000000000000000;
      reg_PECore_RunBias_if_accum_vector_out_data_7_lpi_1_dfm_ftd_12 <= 20'b00000000000000000000;
      reg_PECore_RunBias_if_accum_vector_out_data_10_lpi_1_dfm_ftd_12 <= 20'b00000000000000000000;
      reg_PECore_RunBias_if_accum_vector_out_data_11_lpi_1_dfm_ftd_12 <= 20'b00000000000000000000;
    end
    else if ( PECore_RunBias_if_accum_vector_out_data_and_17_cse ) begin
      reg_PECore_RunBias_if_accum_vector_out_data_6_lpi_1_dfm_ftd_12 <= MUX_v_20_2_2((z_out_31[19:0]),
          (PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_4_sva[19:0]),
          PECore_RunBias_if_accum_vector_out_data_and_15_rgt);
      reg_PECore_RunBias_if_accum_vector_out_data_7_lpi_1_dfm_ftd_12 <= MUX_v_20_2_2((z_out_32[19:0]),
          (PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_5_sva[19:0]),
          PECore_RunBias_if_accum_vector_out_data_and_15_rgt);
      reg_PECore_RunBias_if_accum_vector_out_data_10_lpi_1_dfm_ftd_12 <= MUX_v_20_2_2((z_out_29[19:0]),
          (PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_1_sva[19:0]),
          PECore_RunBias_if_accum_vector_out_data_and_15_rgt);
      reg_PECore_RunBias_if_accum_vector_out_data_11_lpi_1_dfm_ftd_12 <= MUX_v_20_2_2((z_out_30[19:0]),
          (PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_11_sva[19:0]),
          PECore_RunBias_if_accum_vector_out_data_and_15_rgt);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_PECore_RunMac_if_mux_122_ftd_1 <= 4'b0000;
    end
    else if ( PECoreRun_wen & (~(and_4616_cse & PECore_RunMac_if_or_140_m1c)) ) begin
      reg_PECore_RunMac_if_mux_122_ftd_1 <= MUX1HOT_v_4_4_2((rva_in_PopNB_mioi_idat_mxwt[151:148]),
          z_out_50, PEManager_16U_ClusterLookup_1_for_mux_133_nl, (weight_port_read_out_data_7_10_sva_dfm_mx1[3:0]),
          {PECore_RunBias_if_for_and_cse , PECore_RunBias_if_for_and_34_rgt , PECore_RunMac_if_and_569_rgt
          , PECore_RunMac_if_and_570_rgt});
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_PECore_RunMac_if_mux_123_ftd_1 <= 4'b0000;
    end
    else if ( PECore_RunMac_if_and_854_tmp ) begin
      reg_PECore_RunMac_if_mux_123_ftd_1 <= MUX1HOT_v_4_7_2(({crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1_3
          , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1_2 ,
          crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1_1 , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1_0}),
          PECore_DecodeAxiRead_case_4_switch_lp_and_1_nl, adpfloat_tmp_to_fixed_20U_14U_acc_sdt_1_sva_mx0w2,
          (input_mem_banks_bank_array_impl_data0_rsci_q_d[35:32]), (crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38[3:0]),
          PEManager_16U_ClusterLookup_1_for_mux_132_nl, (weight_port_read_out_data_7_11_sva_dfm_mx1[3:0]),
          {and_5134_nl , and_5136_nl , PECore_RunMac_if_and_817_rgt , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_and_1_nl
          , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_and_2_nl , PECore_RunMac_if_and_569_rgt
          , PECore_RunMac_if_and_570_rgt});
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_PECore_RunMac_if_mux_137_ftd_1 <= 2'b00;
      reg_PECore_RunMac_if_mux_139_ftd_1 <= 2'b00;
      reg_PECore_RunMac_if_mux_140_ftd_1 <= 2'b00;
      reg_PECore_RunMac_if_mux_143_ftd_1 <= 7'b0000000;
    end
    else if ( PECore_RunMac_if_and_859_cse ) begin
      reg_PECore_RunMac_if_mux_137_ftd_1 <= MUX1HOT_v_2_4_2(PECore_DecodeAxiRead_case_4_switch_lp_and_9_nl,
          PEManager_16U_ClusterLookup_for_mux_135_nl, (weight_port_read_out_data_8_9_sva_dfm[1:0]),
          (crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1[1:0]),
          {(~ (fsm_output[2])) , PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_398_cse
          , PECore_RunMac_if_and_399_cse});
      reg_PECore_RunMac_if_mux_139_ftd_1 <= MUX1HOT_v_2_4_2(PECore_DecodeAxiRead_case_4_switch_lp_and_7_nl,
          PEManager_16U_ClusterLookup_for_mux_133_nl, (weight_port_read_out_data_8_11_sva_dfm[1:0]),
          (crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1[1:0]),
          {(~ (fsm_output[2])) , PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_398_cse
          , PECore_RunMac_if_and_399_cse});
      reg_PECore_RunMac_if_mux_140_ftd_1 <= MUX1HOT_v_2_4_2(PECore_DecodeAxiRead_case_4_switch_lp_and_6_nl,
          PEManager_16U_ClusterLookup_for_mux_131_nl, (weight_port_read_out_data_8_12_sva_dfm[1:0]),
          (crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1[1:0]),
          {(~ (fsm_output[2])) , PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_398_cse
          , PECore_RunMac_if_and_399_cse});
      reg_PECore_RunMac_if_mux_143_ftd_1 <= MUX1HOT_v_7_4_2(PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_13_nl,
          PEManager_16U_ClusterLookup_for_mux_128_nl, (weight_port_read_out_data_8_15_sva_dfm[6:0]),
          (crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1[6:0]),
          {(~ (fsm_output[2])) , PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_398_cse
          , PECore_RunMac_if_and_399_cse});
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_PECore_RunMac_if_mux_138_ftd_1 <= 5'b00000;
      reg_PECore_RunMac_if_mux_14_ftd_1 <= 5'b00000;
    end
    else if ( PECore_RunMac_if_and_860_cse ) begin
      reg_PECore_RunMac_if_mux_138_ftd_1 <= MUX1HOT_v_5_5_2(PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_12_nl,
          PECore_RunBias_if_for_12_operator_34_true_acc_nl, PEManager_16U_ClusterLookup_for_mux_134_nl,
          (weight_port_read_out_data_8_10_sva_dfm[4:0]), (crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1[4:0]),
          {(fsm_output[1]) , PECore_RunMac_if_and_817_rgt , PECore_RunMac_if_and_569_rgt
          , PECore_RunMac_if_and_390_cse , PECore_RunMac_if_and_391_cse});
      reg_PECore_RunMac_if_mux_14_ftd_1 <= MUX1HOT_v_5_4_2(PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_10_nl,
          z_out_4, PEManager_16U_ClusterLookup_for_mux_132_nl, (weight_port_read_out_data_0_14_sva_dfm_mx1[4:0]),
          {(fsm_output[1]) , PECore_RunMac_if_and_817_rgt , PECore_RunMac_if_and_569_rgt
          , PECore_RunMac_if_and_570_rgt});
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_PECore_RunMac_if_mux_141_ftd_1 <= 5'b00000;
    end
    else if ( PECoreRun_wen & (~((fsm_output[3]) | PECore_RunBias_if_for_and_42_cse))
        ) begin
      reg_PECore_RunMac_if_mux_141_ftd_1 <= MUX1HOT_v_5_5_2(PEManager_16U_ClusterLookup_for_mux_130_nl,
          (weight_port_read_out_data_8_13_sva_dfm[4:0]), (crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1[4:0]),
          PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_11_nl,
          PECore_RunBias_if_for_2_operator_34_true_acc_nl, {PECore_RunMac_if_and_359_cse
          , PECore_RunMac_if_and_360_cse , PECore_RunMac_if_and_361_cse , (fsm_output[1])
          , PECore_RunMac_if_and_803_nl});
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_PECore_RunMac_if_mux_142_ftd_1 <= 4'b0000;
    end
    else if ( PECore_RunMac_if_and_865_tmp ) begin
      reg_PECore_RunMac_if_mux_142_ftd_1 <= MUX1HOT_v_4_7_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl,
          pe_config_manager_counter_sva, (input_mem_banks_bank_array_impl_data0_rsci_q_d[39:36]),
          (crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38[7:4]),
          PEManager_16U_ClusterLookup_for_mux_129_nl, (weight_port_read_out_data_8_14_sva_dfm[3:0]),
          (crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1[3:0]),
          {PECore_RunBias_if_for_and_cse , PECore_RunBias_if_for_and_34_rgt , rva_out_reg_data_and_1_nl
          , PECore_RunMac_if_and_801_nl , PECore_RunMac_if_and_674_rgt , PECore_RunMac_if_and_398_cse
          , PECore_RunMac_if_and_399_cse});
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_Datapath_for_conc_4_ftd <= 8'b00000000;
      reg_Datapath_for_conc_4_ftd_1 <= 8'b00000000;
      reg_Datapath_for_conc_4_ftd_2 <= 8'b00000000;
      reg_Datapath_for_conc_4_ftd_3 <= 8'b00000000;
      reg_Datapath_for_conc_4_ftd_4 <= 8'b00000000;
      reg_Datapath_for_conc_4_ftd_5 <= 8'b00000000;
      reg_Datapath_for_conc_4_ftd_6 <= 8'b00000000;
      reg_Datapath_for_conc_4_ftd_7 <= 8'b00000000;
      reg_Datapath_for_conc_4_ftd_8 <= 8'b00000000;
      reg_Datapath_for_conc_4_ftd_9 <= 8'b00000000;
      reg_Datapath_for_conc_4_ftd_10 <= 8'b00000000;
      reg_Datapath_for_conc_4_ftd_11 <= 8'b00000000;
      reg_Datapath_for_conc_4_ftd_12 <= 8'b00000000;
      reg_Datapath_for_conc_4_ftd_13 <= 8'b00000000;
      reg_Datapath_for_conc_4_ftd_14 <= 8'b00000000;
      reg_Datapath_for_conc_4_ftd_15 <= 8'b00000000;
    end
    else if ( Datapath_for_and_enex5 ) begin
      reg_Datapath_for_conc_4_ftd <= PECore_RunMac_if_mux_31_itm;
      reg_Datapath_for_conc_4_ftd_1 <= PECore_RunMac_if_mux_30_itm;
      reg_Datapath_for_conc_4_ftd_2 <= PECore_RunMac_if_mux_29_itm;
      reg_Datapath_for_conc_4_ftd_3 <= PECore_RunMac_if_mux_28_itm;
      reg_Datapath_for_conc_4_ftd_4 <= PECore_RunMac_if_mux_27_itm;
      reg_Datapath_for_conc_4_ftd_5 <= PECore_RunMac_if_mux_26_itm;
      reg_Datapath_for_conc_4_ftd_6 <= PECore_RunMac_if_mux_25_itm;
      reg_Datapath_for_conc_4_ftd_7 <= PECore_RunMac_if_mux_24_itm;
      reg_Datapath_for_conc_4_ftd_8 <= PECore_RunMac_if_mux_23_itm;
      reg_Datapath_for_conc_4_ftd_9 <= PECore_RunMac_if_mux_22_itm;
      reg_Datapath_for_conc_4_ftd_10 <= PECore_RunMac_if_mux_21_itm;
      reg_Datapath_for_conc_4_ftd_11 <= PECore_RunMac_if_mux_20_itm;
      reg_Datapath_for_conc_4_ftd_12 <= PECore_RunMac_if_mux_19_itm;
      reg_Datapath_for_conc_4_ftd_13 <= PECore_RunMac_if_mux_18_itm;
      reg_Datapath_for_conc_4_ftd_14 <= PECore_RunMac_if_mux_17_itm;
      reg_Datapath_for_conc_4_ftd_15 <= PECore_RunMac_if_mux_16_itm;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_PECore_RunMac_if_mux_123_1_enexo <= 1'b1;
    end
    else if ( PECore_RunMac_if_and_854_tmp | PECore_PushAxiRsp_if_and_47_enex5 )
        begin
      reg_PECore_RunMac_if_mux_123_1_enexo <= PECore_RunMac_if_and_854_tmp;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_PECore_RunMac_if_mux_142_1_enexo <= 1'b1;
    end
    else if ( PECore_RunMac_if_and_865_tmp | PECore_PushAxiRsp_if_and_48_enex5 )
        begin
      reg_PECore_RunMac_if_mux_142_1_enexo <= PECore_RunMac_if_and_865_tmp;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_47_40_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_91_cse | PECore_PushAxiRsp_if_and_49_enex5 ) begin
      reg_rva_out_reg_data_47_40_sva_dfm_4_enexo <= rva_out_reg_data_and_91_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_91_cse | PECore_PushAxiRsp_if_and_50_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_enexo <= rva_out_reg_data_and_91_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_63_56_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_91_cse | PECore_PushAxiRsp_if_and_51_enex5 ) begin
      reg_rva_out_reg_data_63_56_sva_dfm_4_enexo <= rva_out_reg_data_and_91_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_71_64_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_91_cse | PECore_PushAxiRsp_if_and_52_enex5 ) begin
      reg_rva_out_reg_data_71_64_sva_dfm_4_enexo <= rva_out_reg_data_and_91_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_72_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_91_cse | PECore_PushAxiRsp_if_and_53_enex5 ) begin
      reg_rva_out_reg_data_79_72_sva_dfm_4_enexo <= rva_out_reg_data_and_91_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_91_cse | PECore_PushAxiRsp_if_and_54_enex5 ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_enexo <= rva_out_reg_data_and_91_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_95_88_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_91_cse | PECore_PushAxiRsp_if_and_55_enex5 ) begin
      reg_rva_out_reg_data_95_88_sva_dfm_4_enexo <= rva_out_reg_data_and_91_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_91_cse | PECore_PushAxiRsp_if_and_56_enex5 ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_enexo <= rva_out_reg_data_and_91_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_111_104_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_91_cse | PECore_PushAxiRsp_if_and_57_enex5 ) begin
      reg_rva_out_reg_data_111_104_sva_dfm_4_enexo <= rva_out_reg_data_and_91_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_119_112_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_91_cse | PECore_PushAxiRsp_if_and_58_enex5 ) begin
      reg_rva_out_reg_data_119_112_sva_dfm_4_enexo <= rva_out_reg_data_and_91_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_127_120_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_91_cse | PECore_PushAxiRsp_if_and_59_enex5 ) begin
      reg_rva_out_reg_data_127_120_sva_dfm_4_enexo <= rva_out_reg_data_and_91_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_0_enexo <= 1'b1;
    end
    else if ( accum_vector_data_and_9_cse | PECore_PushOutput_if_and_16_enex5 ) begin
      reg_act_port_reg_data_0_enexo <= accum_vector_data_and_9_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_1_enexo <= 1'b1;
    end
    else if ( is_start_and_cse | PECore_PushOutput_if_and_17_enex5 ) begin
      reg_act_port_reg_data_1_enexo <= is_start_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_2_enexo <= 1'b1;
    end
    else if ( is_start_and_cse | PECore_PushOutput_if_and_18_enex5 ) begin
      reg_act_port_reg_data_2_enexo <= is_start_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_3_enexo <= 1'b1;
    end
    else if ( is_start_and_cse | PECore_PushOutput_if_and_19_enex5 ) begin
      reg_act_port_reg_data_3_enexo <= is_start_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_4_enexo <= 1'b1;
    end
    else if ( is_start_and_cse | PECore_PushOutput_if_and_20_enex5 ) begin
      reg_act_port_reg_data_4_enexo <= is_start_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_5_enexo <= 1'b1;
    end
    else if ( act_port_reg_data_and_8_cse | PECore_PushOutput_if_and_21_enex5 ) begin
      reg_act_port_reg_data_5_enexo <= act_port_reg_data_and_8_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_6_enexo <= 1'b1;
    end
    else if ( act_port_reg_data_and_8_cse | PECore_PushOutput_if_and_22_enex5 ) begin
      reg_act_port_reg_data_6_enexo <= act_port_reg_data_and_8_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_9_enexo <= 1'b1;
    end
    else if ( act_port_reg_data_and_8_cse | PECore_PushOutput_if_and_25_enex5 ) begin
      reg_act_port_reg_data_9_enexo <= act_port_reg_data_and_8_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_10_enexo <= 1'b1;
    end
    else if ( act_port_reg_data_and_8_cse | PECore_PushOutput_if_and_26_enex5 ) begin
      reg_act_port_reg_data_10_enexo <= act_port_reg_data_and_8_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_asn_3_enexo <= 1'b1;
    end
    else if ( act_port_reg_data_and_29_enex5 | PECore_PushOutput_if_and_28_enex5
        ) begin
      reg_act_port_reg_data_asn_3_enexo <= act_port_reg_data_and_29_enex5;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_asn_2_enexo <= 1'b1;
    end
    else if ( act_port_reg_data_and_28_enex5 | PECore_PushOutput_if_and_29_enex5
        ) begin
      reg_act_port_reg_data_asn_2_enexo <= act_port_reg_data_and_28_enex5;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_asn_1_enexo <= 1'b1;
    end
    else if ( act_port_reg_data_and_enex5 | PECore_PushOutput_if_and_30_enex5 ) begin
      reg_act_port_reg_data_asn_1_enexo <= act_port_reg_data_and_enex5;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_asn_enexo <= 1'b1;
    end
    else if ( act_port_reg_data_and_30_enex5 | PECore_PushOutput_if_and_31_enex5
        ) begin
      reg_act_port_reg_data_asn_enexo <= act_port_reg_data_and_30_enex5;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_14_enexo <= 1'b1;
    end
    else if ( and_5872_cse | act_port_reg_data_and_enex5 ) begin
      reg_act_port_reg_data_14_enexo <= and_5872_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_13_enexo <= 1'b1;
    end
    else if ( and_5872_cse | act_port_reg_data_and_28_enex5 ) begin
      reg_act_port_reg_data_13_enexo <= and_5872_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_12_enexo <= 1'b1;
    end
    else if ( and_5872_cse | act_port_reg_data_and_29_enex5 ) begin
      reg_act_port_reg_data_12_enexo <= and_5872_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_15_enexo <= 1'b1;
    end
    else if ( and_5872_cse | act_port_reg_data_and_30_enex5 ) begin
      reg_act_port_reg_data_15_enexo <= and_5872_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_PECore_RunMac_if_mux_31_enexo <= 1'b1;
    end
    else if ( PECore_RunMac_if_and_cse | Datapath_for_and_enex5 ) begin
      reg_PECore_RunMac_if_mux_31_enexo <= PECore_RunMac_if_and_cse;
    end
  end
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_or_1_nl
      = input_read_req_valid_lpi_1_dfm_6 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
  assign PECore_DecodeAxi_if_mux_67_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_or_1_nl,
      input_read_req_valid_lpi_1_dfm_6, rva_in_PopNB_mioi_idat_mxwt[168]);
  assign PECore_DecodeAxi_mux_133_nl = MUX_s_1_2_2(input_read_req_valid_lpi_1_dfm_6,
      PECore_DecodeAxi_if_mux_67_nl, rva_in_PopNB_mioi_ivld_mxwt);
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_or_nl
      = input_write_req_valid_lpi_1_dfm_6 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
  assign PECore_DecodeAxi_if_mux_125_nl = MUX_s_1_2_2(input_write_req_valid_lpi_1_dfm_6,
      PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_or_nl,
      rva_in_PopNB_mioi_idat_mxwt[168]);
  assign PECore_DecodeAxi_mux_138_nl = MUX_s_1_2_2(input_write_req_valid_lpi_1_dfm_6,
      PECore_DecodeAxi_if_mux_125_nl, rva_in_PopNB_mioi_ivld_mxwt);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_258_nl = MUX_s_1_16_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[9]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[10]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]), crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_lpi_1_dfm_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_257_nl = MUX_s_1_16_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[9]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[10]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]), {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_15_lpi_1_dfm_1_3_1
      , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_15_lpi_1_dfm_1_0});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_256_nl = MUX_s_1_16_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[9]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[10]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]), crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_14_lpi_1_dfm_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_255_nl = MUX_s_1_16_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[9]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[10]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]), {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_13_3_2_lpi_1_dfm_1
      , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_13_1_0_lpi_1_dfm_1});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_254_nl = MUX_s_1_16_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[9]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[10]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]), crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_12_lpi_1_dfm_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_251_nl = MUX_s_1_16_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[9]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[10]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]), {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm_1
      , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_2_0_lpi_1_dfm_1});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_250_nl = MUX_s_1_16_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[9]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[10]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]), crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_8_lpi_1_dfm_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_249_nl = MUX_s_1_16_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[9]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[10]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]), {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_3_1_lpi_1_dfm_1
      , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm_1});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_248_nl = MUX_s_1_16_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[9]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[10]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]), crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_6_lpi_1_dfm_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_247_nl = MUX_s_1_16_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[9]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[10]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]), {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_5_3_2_lpi_1_dfm_1
      , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_5_1_0_lpi_1_dfm_1});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_246_nl = MUX_s_1_16_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[9]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[10]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]), crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_4_lpi_1_dfm_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_245_nl = MUX_s_1_16_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[9]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[10]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]), {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_3_1_lpi_1_dfm_1
      , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm_1});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_244_nl = MUX_s_1_16_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[9]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[10]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]), crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_2_lpi_1_dfm_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_253_nl = MUX_s_1_16_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[9]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[10]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]), {crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_3_1_lpi_1_dfm_1
      , crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm_1});
  assign PEManager_16U_ClusterLookup_for_mux_15_nl = MUX_v_3_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:5]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_0_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_6_nl = MUX_v_3_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:5]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_5_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_3_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_6_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_74_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_1_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_72_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_1_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_70_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_2_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_68_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_2_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_66_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_3_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_64_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_3_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_65_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_4_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_53_nl = MUX_v_4_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:4]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_13_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_5_nl = MUX_v_4_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:4]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_5_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_138_nl = MUX_v_4_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[3:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_5_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_55_nl = MUX_v_4_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:4]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_13_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_57_nl = MUX_v_4_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:4]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_14_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_59_nl = MUX_v_4_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:4]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_14_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_61_nl = MUX_v_4_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:4]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_15_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_63_nl = MUX_v_4_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:4]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_15_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_78_nl = MUX_v_4_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:4]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_0_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_137_nl = MUX_v_4_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[3:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_0_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_76_nl = MUX_v_4_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:4]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_0_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_136_nl = MUX_v_4_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[3:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_0_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_67_nl = MUX_v_6_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:2]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_4_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_69_nl = MUX_v_3_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:5]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_5_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_71_nl = MUX_v_6_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:2]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_5_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_2_nl = MUX_v_3_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:5]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_7_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_73_nl = MUX_v_6_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:2]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:2]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:2]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_6_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_75_nl = MUX_v_3_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:5]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_6_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_77_nl = MUX_v_4_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:4]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:4]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:4]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_7_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_79_nl = MUX_s_1_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_7_sva_dfm_mx1[7:4])});
  assign PECore_DecodeAxiRead_switch_lp_mux_11_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[0]),
      PECore_DecodeAxiRead_case_4_switch_lp_and_5_itm, PECore_DecodeAxiRead_switch_lp_equal_tmp_5);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_19_nl
      = PECore_DecodeAxiRead_switch_lp_mux_11_nl & PECore_DecodeAxiRead_switch_lp_nor_10_cse_1;
  assign PECore_DecodeAxi_if_mux_74_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_19_nl,
      PECore_DecodeAxiRead_case_4_switch_lp_and_2_itm, rva_in_PopNB_mio_mrgout_dat_sva[168]);
  assign PECore_DecodeAxi_mux_139_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_case_4_switch_lp_and_2_itm,
      PECore_DecodeAxi_if_mux_74_nl, PECore_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva);
  assign PECore_PushAxiRsp_if_else_mux_14_nl = MUX_s_1_2_2(PECore_DecodeAxi_mux_139_nl,
      (input_mem_banks_read_read_data_lpi_1[0]), input_mem_banks_load_store_for_else_and_cse);
  assign PECore_DecodeAxiRead_switch_lp_mux_8_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[8]),
      PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm, PECore_DecodeAxiRead_switch_lp_equal_tmp_5);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_17_nl
      = PECore_DecodeAxiRead_switch_lp_mux_8_nl & PECore_DecodeAxiRead_switch_lp_nor_10_cse_1;
  assign PECore_DecodeAxi_if_mux_126_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_17_nl,
      PECore_DecodeAxiRead_case_4_switch_lp_and_itm, rva_in_PopNB_mio_mrgout_dat_sva[168]);
  assign PECore_DecodeAxi_mux_141_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_case_4_switch_lp_and_itm,
      PECore_DecodeAxi_if_mux_126_nl, PECore_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva);
  assign PECore_PushAxiRsp_if_else_mux_15_nl = MUX_s_1_2_2(PECore_DecodeAxi_mux_141_nl,
      (input_mem_banks_read_read_data_lpi_1[8]), input_mem_banks_load_store_for_else_and_cse);
  assign PECore_DecodeAxiRead_switch_lp_mux_5_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[16]),
      PECore_DecodeAxiRead_case_4_switch_lp_and_2_itm, PECore_DecodeAxiRead_switch_lp_equal_tmp_5);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_13_nl
      = PECore_DecodeAxiRead_switch_lp_mux_5_nl & PECore_DecodeAxiRead_switch_lp_nor_10_cse_1;
  assign PECore_DecodeAxi_if_mux_127_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_13_nl,
      PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm, rva_in_PopNB_mio_mrgout_dat_sva[168]);
  assign PECore_DecodeAxi_mux_143_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm,
      PECore_DecodeAxi_if_mux_127_nl, PECore_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva);
  assign PECore_PushAxiRsp_if_else_mux_16_nl = MUX_s_1_2_2(PECore_DecodeAxi_mux_143_nl,
      (input_mem_banks_read_read_data_lpi_1[16]), input_mem_banks_load_store_for_else_and_cse);
  assign PECore_DecodeAxiRead_switch_lp_mux_12_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[24]),
      PECore_DecodeAxiRead_case_4_switch_lp_and_itm, PECore_DecodeAxiRead_switch_lp_equal_tmp_5);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl =
      PECore_DecodeAxiRead_switch_lp_mux_12_nl & PECore_DecodeAxiRead_switch_lp_nor_10_cse_1;
  assign PECore_DecodeAxi_if_mux_128_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl,
      PECore_DecodeAxiRead_case_4_switch_lp_and_5_itm, rva_in_PopNB_mio_mrgout_dat_sva[168]);
  assign PECore_DecodeAxi_mux_145_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_case_4_switch_lp_and_5_itm,
      PECore_DecodeAxi_if_mux_128_nl, PECore_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva);
  assign PECore_PushAxiRsp_if_else_mux_17_nl = MUX_s_1_2_2(PECore_DecodeAxi_mux_145_nl,
      (input_mem_banks_read_read_data_lpi_1[24]), input_mem_banks_load_store_for_else_and_cse);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_18_nl
      = MUX_v_7_2_2(7'b0000000, (SC_SRAM_CONFIG[7:1]), PECore_DecodeAxiRead_switch_lp_nor_10_cse_1);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl
      = MUX_v_2_2_2(2'b00, (SC_SRAM_CONFIG[10:9]), PECore_DecodeAxiRead_switch_lp_nor_10_cse_1);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_15_nl
      = MUX_v_5_2_2(5'b00000, (SC_SRAM_CONFIG[15:11]), PECore_DecodeAxiRead_switch_lp_nor_10_cse_1);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_12_nl
      = MUX_v_2_2_2(2'b00, (SC_SRAM_CONFIG[18:17]), PECore_DecodeAxiRead_switch_lp_nor_10_cse_1);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_10_nl
      = MUX_v_5_2_2(5'b00000, (SC_SRAM_CONFIG[23:19]), PECore_DecodeAxiRead_switch_lp_nor_10_cse_1);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_9_nl =
      MUX_v_2_2_2(2'b00, (SC_SRAM_CONFIG[26:25]), PECore_DecodeAxiRead_switch_lp_nor_10_cse_1);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl
      = MUX_v_5_2_2(5'b00000, (SC_SRAM_CONFIG[31:27]), PECore_DecodeAxiRead_switch_lp_nor_10_cse_1);
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_7_nl = or_1521_cse
      & PECore_UpdateFSM_case_4_is_output_end_pe_config_UpdateManagerCounter_nand_itm;
  assign PECore_UpdateFSM_switch_lp_mux_6_nl = MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_7_nl,
      or_1521_cse, PECore_UpdateFSM_switch_lp_unequal_tmp);
  assign and_3383_nl = (~ state_2_0_sva_2) & (fsm_output[4]);
  assign PECore_UpdateFSM_switch_lp_mux1h_42_nl = MUX1HOT_s_1_3_2(or_1521_cse, PECore_RunMac_nor_tmp,
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_pe_config_UpdateInputCounter_if_nor_svs,
      {PECore_RunFSM_switch_lp_equal_tmp , PECore_UpdateFSM_switch_lp_equal_tmp_1
      , PECore_RunFSM_switch_lp_equal_tmp_1});
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_252_nl = MUX_s_1_16_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[8]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[9]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[10]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[11]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[12]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[13]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[14]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]), crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_10_lpi_1_dfm_1);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_for_if_1_crossbar_spec_PE_Weight_WordType_16U_16U_for_if_1_crossbar_spec_PE_Weight_WordType_16U_16U_for_if_1_nor_5_nl
      = ~(crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_252_nl | (~ weight_read_ack_9_lpi_1_dfm_15_mx0));
  assign pe_config_UpdateManagerCounter_if_not_7_nl = ~ pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_nor_svs_1;
  assign pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_and_1_nl =
      MUX_v_4_2_2(4'b0000, (z_out_4[3:0]), pe_config_UpdateManagerCounter_if_not_7_nl);
  assign and_3501_nl = and_5844_cse & (fsm_output[1]);
  assign while_and_202_nl = and_dcpl_700 & while_and_81_m1c;
  assign while_and_203_nl = and_dcpl_702 & while_and_81_m1c;
  assign while_and_204_nl = or_dcpl_370 & while_and_81_m1c;
  assign PECore_RunBias_if_for_and_25_nl = z_out_21_32 & (~ PECore_RunBias_if_for_13_operator_32_true_slc_operator_32_true_acc_13_svs_mx1)
      & while_and_48_tmp_1;
  assign while_and_82_nl = PECore_RunBias_if_for_13_operator_32_true_slc_operator_32_true_acc_13_svs_mx1
      & while_and_48_tmp_1;
  assign while_while_mux1h_12_nl = MUX1HOT_v_20_5_2((z_out_29[19:0]), (PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_1_sva[19:0]),
      (PECore_RunBias_if_accum_vector_out_data_13_lpi_1_dfm[19:0]), 20'b10000000000000000001,
      20'b01111111111111111111, {while_and_202_nl , while_and_203_nl , while_and_204_nl
      , PECore_RunBias_if_for_and_25_nl , while_and_82_nl});
  assign PECore_UpdateFSM_switch_lp_not_36_nl = ~ and_5871_cse;
  assign while_and_199_nl = and_dcpl_700 & while_and_83_m1c;
  assign while_and_200_nl = and_dcpl_702 & while_and_83_m1c;
  assign while_and_201_nl = or_dcpl_370 & while_and_83_m1c;
  assign PECore_RunBias_if_for_and_27_nl = z_out_24_32 & (~ PECore_RunBias_if_for_14_operator_32_true_slc_operator_32_true_acc_13_svs_mx1)
      & while_and_48_tmp_1;
  assign while_and_84_nl = PECore_RunBias_if_for_14_operator_32_true_slc_operator_32_true_acc_13_svs_mx1
      & while_and_48_tmp_1;
  assign while_while_mux1h_13_nl = MUX1HOT_v_20_5_2((z_out_30[19:0]), (PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_11_sva[19:0]),
      (PECore_RunBias_if_accum_vector_out_data_14_lpi_1_dfm[19:0]), 20'b10000000000000000001,
      20'b01111111111111111111, {while_and_199_nl , while_and_200_nl , while_and_201_nl
      , PECore_RunBias_if_for_and_27_nl , while_and_84_nl});
  assign PECore_UpdateFSM_switch_lp_not_64_nl = ~ and_5871_cse;
  assign while_and_196_nl = and_dcpl_700 & while_and_85_m1c;
  assign while_and_197_nl = and_dcpl_702 & while_and_85_m1c;
  assign while_and_198_nl = or_dcpl_370 & while_and_85_m1c;
  assign PECore_RunBias_if_for_and_29_nl = z_out_23_32 & (~ PECore_RunBias_if_for_15_operator_32_true_slc_operator_32_true_acc_13_svs_mx1)
      & while_and_48_tmp_1;
  assign while_and_86_nl = PECore_RunBias_if_for_15_operator_32_true_slc_operator_32_true_acc_13_svs_mx1
      & while_and_48_tmp_1;
  assign while_while_mux1h_14_nl = MUX1HOT_v_20_5_2((z_out_31[19:0]), (PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_4_sva[19:0]),
      (PECore_RunBias_if_accum_vector_out_data_15_lpi_1_dfm[19:0]), 20'b10000000000000000001,
      20'b01111111111111111111, {while_and_196_nl , while_and_197_nl , while_and_198_nl
      , PECore_RunBias_if_for_and_29_nl , while_and_86_nl});
  assign PECore_UpdateFSM_switch_lp_not_63_nl = ~ and_5871_cse;
  assign while_and_193_nl = and_dcpl_700 & while_and_87_m1c;
  assign while_and_194_nl = and_dcpl_702 & while_and_87_m1c;
  assign while_and_195_nl = or_dcpl_370 & while_and_87_m1c;
  assign PECore_RunBias_if_for_and_31_nl = z_out_22_32 & (~ PECore_RunBias_if_for_16_operator_32_true_slc_operator_32_true_acc_13_svs_mx1)
      & while_and_48_tmp_1;
  assign while_and_88_nl = PECore_RunBias_if_for_16_operator_32_true_slc_operator_32_true_acc_13_svs_mx1
      & while_and_48_tmp_1;
  assign while_while_mux1h_15_nl = MUX1HOT_v_20_5_2((z_out_32[19:0]), (PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_5_sva[19:0]),
      (PECore_RunBias_if_accum_vector_out_data_lpi_1_dfm[19:0]), 20'b10000000000000000001,
      20'b01111111111111111111, {while_and_193_nl , while_and_194_nl , while_and_195_nl
      , PECore_RunBias_if_for_and_31_nl , while_and_88_nl});
  assign PECore_UpdateFSM_switch_lp_not_62_nl = ~ and_5871_cse;
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl
      = pe_config_is_zero_first_sva_dfm_4_mx0 & (~ pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1);
  assign pe_config_UpdateManagerCounter_mux_1_nl = MUX_s_1_2_2(pe_config_is_zero_first_sva_dfm_4_mx0,
      pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl,
      pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_nor_svs_1);
  assign PECore_UpdateFSM_switch_lp_mux_7_nl = MUX_s_1_2_2(pe_config_UpdateManagerCounter_mux_1_nl,
      pe_config_is_zero_first_sva_dfm_4_mx0, PECore_UpdateFSM_switch_lp_unequal_tmp_1);
  assign and_3991_nl = (~ state_2_0_sva_2) & (fsm_output[1]);
  assign pe_config_UpdateInputCounter_if_not_2_nl = ~ pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_pe_config_UpdateInputCounter_if_nor_svs_1;
  assign pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl = MUX_v_8_2_2(8'b00000000,
      z_out_5, pe_config_UpdateInputCounter_if_not_2_nl);
  assign PECore_UpdateFSM_switch_lp_and_nl = (~ or_dcpl_724) & and_4031_m1c;
  assign pe_config_UpdateManagerCounter_if_not_9_nl = ~ pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1;
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl
      = MUX_v_8_2_2(8'b00000000, z_out_5, pe_config_UpdateManagerCounter_if_not_9_nl);
  assign and_4037_nl = and_5844_cse & pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_nor_svs_1
      & (fsm_output[1]);
  assign PEManager_16U_ClusterLookup_for_mux_94_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_0_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_92_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_0_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_90_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_1_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_88_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_1_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_86_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_2_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_84_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_2_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_82_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_3_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_80_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_3_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_81_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_4_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_83_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_4_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_85_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_5_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_87_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_5_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_89_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_6_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_91_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_6_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_93_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_7_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_95_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_7_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_78_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_8_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_76_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_8_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_74_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_9_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_72_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_9_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_70_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_10_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_68_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_10_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_66_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_11_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_64_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_11_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_65_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_12_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_67_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_12_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_69_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_13_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_71_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_13_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_73_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_14_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_75_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_14_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_77_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_15_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_79_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_15_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_62_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_0_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_60_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_0_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_58_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_1_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_56_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_1_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_55_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_5_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_57_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_6_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_59_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_6_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_61_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_7_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_63_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_7_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_46_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_8_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_44_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_8_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_42_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_9_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_40_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_9_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_38_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_10_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_36_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_10_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_34_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_11_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_32_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_11_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_33_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_12_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_35_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_12_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_37_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_13_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_39_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_13_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_41_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_14_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_43_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_14_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_45_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_15_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_47_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_15_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_54_nl = MUX_v_3_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:5]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_2_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_52_nl = MUX_v_3_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:5]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_2_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_48_nl = MUX_v_3_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:5]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_3_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_49_nl = MUX_v_3_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:5]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_4_sva_dfm_mx1[3:0])});
  assign nl_PECore_RunBias_if_for_10_operator_33_true_acc_nl = (operator_4_false_acc_psp_10_sva_1[3:1])
      + 3'b111;
  assign PECore_RunBias_if_for_10_operator_33_true_acc_nl = nl_PECore_RunBias_if_for_10_operator_33_true_acc_nl[2:0];
  assign nl_PECore_RunBias_if_for_10_operator_34_true_acc_nl = conv_s2s_4_5({PECore_RunBias_if_for_10_operator_33_true_acc_nl
      , (operator_4_false_acc_psp_10_sva_1[0])}) + 5'b00111;
  assign PECore_RunBias_if_for_10_operator_34_true_acc_nl = nl_PECore_RunBias_if_for_10_operator_34_true_acc_nl[4:0];
  assign PEManager_16U_ClusterLookup_for_mux_139_nl = MUX_v_5_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[4:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_2_sva_dfm_mx1[3:0])});
  assign nl_PECore_RunBias_if_for_11_operator_33_true_acc_nl = (operator_4_false_acc_psp_11_sva_1[3:1])
      + 3'b111;
  assign PECore_RunBias_if_for_11_operator_33_true_acc_nl = nl_PECore_RunBias_if_for_11_operator_33_true_acc_nl[2:0];
  assign nl_PECore_RunBias_if_for_11_operator_34_true_acc_nl = conv_s2s_4_5({PECore_RunBias_if_for_11_operator_33_true_acc_nl
      , (operator_4_false_acc_psp_11_sva_1[0])}) + 5'b00111;
  assign PECore_RunBias_if_for_11_operator_34_true_acc_nl = nl_PECore_RunBias_if_for_11_operator_34_true_acc_nl[4:0];
  assign PEManager_16U_ClusterLookup_for_mux_140_nl = MUX_v_5_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[4:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_2_sva_dfm_mx1[7:4])});
  assign nl_PECore_RunBias_if_for_6_operator_33_true_acc_nl = (operator_4_false_acc_psp_6_sva_1[3:1])
      + 3'b111;
  assign PECore_RunBias_if_for_6_operator_33_true_acc_nl = nl_PECore_RunBias_if_for_6_operator_33_true_acc_nl[2:0];
  assign nl_PECore_RunBias_if_for_6_operator_34_true_acc_nl = conv_s2s_4_5({PECore_RunBias_if_for_6_operator_33_true_acc_nl
      , (operator_4_false_acc_psp_6_sva_1[0])}) + 5'b00111;
  assign PECore_RunBias_if_for_6_operator_34_true_acc_nl = nl_PECore_RunBias_if_for_6_operator_34_true_acc_nl[4:0];
  assign PEManager_16U_ClusterLookup_for_mux_142_nl = MUX_v_5_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[4:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_3_sva_dfm_mx1[7:4])});
  assign nl_PECore_RunBias_if_for_7_operator_33_true_acc_nl = (operator_4_false_acc_psp_7_sva_1[3:1])
      + 3'b111;
  assign PECore_RunBias_if_for_7_operator_33_true_acc_nl = nl_PECore_RunBias_if_for_7_operator_33_true_acc_nl[2:0];
  assign nl_PECore_RunBias_if_for_7_operator_34_true_acc_nl = conv_s2s_4_5({PECore_RunBias_if_for_7_operator_33_true_acc_nl
      , (operator_4_false_acc_psp_7_sva_1[0])}) + 5'b00111;
  assign PECore_RunBias_if_for_7_operator_34_true_acc_nl = nl_PECore_RunBias_if_for_7_operator_34_true_acc_nl[4:0];
  assign PEManager_16U_ClusterLookup_for_mux_143_nl = MUX_v_5_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[4:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_4_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_50_nl = MUX_v_3_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[7:5]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[7:5]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[7:5]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_3_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_141_nl = MUX_v_5_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[4:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_3_sva_dfm_mx1[3:0])});
  assign nl_PECore_RunBias_if_for_5_operator_33_true_acc_nl = (operator_4_false_acc_psp_5_sva_1[3:1])
      + 3'b111;
  assign PECore_RunBias_if_for_5_operator_33_true_acc_nl = nl_PECore_RunBias_if_for_5_operator_33_true_acc_nl[2:0];
  assign nl_PECore_RunBias_if_for_5_operator_34_true_acc_nl = conv_s2s_4_5({PECore_RunBias_if_for_5_operator_33_true_acc_nl
      , (operator_4_false_acc_psp_5_sva_1[0])}) + 5'b00111;
  assign PECore_RunBias_if_for_5_operator_34_true_acc_nl = nl_PECore_RunBias_if_for_5_operator_34_true_acc_nl[4:0];
  assign PECore_RunMac_if_and_829_nl = (~ (fsm_output[3])) & PECore_RunMac_if_or_143_m1c;
  assign PEManager_16U_ClusterLookup_for_mux_51_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_4_sva_dfm_mx1[7:4])});
  assign nl_PECore_RunBias_if_for_8_operator_33_true_acc_nl = (operator_4_false_acc_psp_8_sva_1[3:1])
      + 3'b111;
  assign PECore_RunBias_if_for_8_operator_33_true_acc_nl = nl_PECore_RunBias_if_for_8_operator_33_true_acc_nl[2:0];
  assign nl_PECore_RunBias_if_for_8_operator_34_true_acc_nl = conv_s2u_4_5({PECore_RunBias_if_for_8_operator_33_true_acc_nl
      , (operator_4_false_acc_psp_8_sva_1[0])}) + 5'b00111;
  assign PECore_RunBias_if_for_8_operator_34_true_acc_nl = nl_PECore_RunBias_if_for_8_operator_34_true_acc_nl[4:0];
  assign PEManager_16U_ClusterLookup_for_mux_53_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_5_sva_dfm_mx1[3:0])});
  assign nl_PECore_RunBias_if_for_9_operator_33_true_acc_nl = (operator_4_false_acc_psp_9_sva_1[3:1])
      + 3'b111;
  assign PECore_RunBias_if_for_9_operator_33_true_acc_nl = nl_PECore_RunBias_if_for_9_operator_33_true_acc_nl[2:0];
  assign nl_PECore_RunBias_if_for_9_operator_34_true_acc_nl = conv_s2u_4_5({PECore_RunBias_if_for_9_operator_33_true_acc_nl
      , (operator_4_false_acc_psp_9_sva_1[0])}) + 5'b00111;
  assign PECore_RunBias_if_for_9_operator_34_true_acc_nl = nl_PECore_RunBias_if_for_9_operator_34_true_acc_nl[4:0];
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux1h_6_nl = MUX1HOT_s_1_5_2(pe_config_is_cluster_sva,
      (pe_manager_adplfloat_bias_bias_0_sva[0]), crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm,
      (pe_manager_adplfloat_bias_bias_1_sva[0]), pe_manager_cluster_lut_data_1_2_sva_0,
      {PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_5 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5});
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_2_nl = PECore_DecodeAxiRead_case_4_switch_lp_mux1h_6_nl
      & (~ PECore_DecodeAxiWrite_case_4_switch_lp_nor_tmp_1);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux1h_13_nl = MUX1HOT_s_1_5_2(pe_config_is_valid_sva,
      pe_manager_zero_active_0_sva, crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm,
      pe_manager_zero_active_1_sva, pe_manager_cluster_lut_data_1_0_sva_0, {PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_5
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5});
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux1h_11_nl = MUX1HOT_s_1_5_2(pe_config_is_zero_first_sva,
      (pe_manager_adplfloat_bias_weight_0_sva[0]), crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm,
      (pe_manager_adplfloat_bias_weight_1_sva[0]), pe_manager_cluster_lut_data_1_1_sva_0,
      {PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_5 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5});
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux1h_16_nl = MUX1HOT_s_1_5_2(pe_config_is_bias_sva,
      (pe_manager_adplfloat_bias_input_0_sva[0]), crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm,
      (pe_manager_adplfloat_bias_input_1_sva[0]), pe_manager_cluster_lut_data_1_3_sva_0,
      {PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_5 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5});
  assign PECore_RunBias_if_for_and_49_nl = is_start_sva & or_3399_cse;
  assign PECore_RunBias_if_for_and_40_nl = is_start_sva & or_dcpl_251;
  assign PECore_RunBias_if_for_and_36_nl = is_start_sva & (fsm_output[3]);
  assign adpfloat_tmp_is_zero_if_adpfloat_tmp_is_zero_if_nor_nl = ~((input_mem_banks_write_if_for_if_mux_cse[6:0]!=7'b0000000));
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_7_nl = MUX_v_8_2_2(pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_12_sva_dfm_4, PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_29_nl
      = PECore_DecodeAxiRead_case_4_switch_lp_mux_7_nl & ({{7{PECore_DecodeAxiRead_case_4_switch_lp_nor_13_cse_1}},
      PECore_DecodeAxiRead_case_4_switch_lp_nor_13_cse_1}) & ({{7{PECore_DecodeAxiRead_switch_lp_nor_14_cse_1}},
      PECore_DecodeAxiRead_switch_lp_nor_14_cse_1});
  assign PEManager_16U_ClusterLookup_1_for_mux_62_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_8_sva_dfm_mx1[3:0])});
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_8_nl = MUX_v_8_2_2(pe_manager_cluster_lut_data_0_13_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_28_nl
      = PECore_DecodeAxiRead_case_4_switch_lp_mux_8_nl & ({{7{PECore_DecodeAxiRead_case_4_switch_lp_nor_13_cse_1}},
      PECore_DecodeAxiRead_case_4_switch_lp_nor_13_cse_1}) & ({{7{PECore_DecodeAxiRead_switch_lp_nor_14_cse_1}},
      PECore_DecodeAxiRead_switch_lp_nor_14_cse_1});
  assign PEManager_16U_ClusterLookup_1_for_mux_60_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_8_sva_dfm_mx1[7:4])});
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_9_nl = MUX_v_8_2_2(pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_14_sva_dfm_4, PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_27_nl
      = PECore_DecodeAxiRead_case_4_switch_lp_mux_9_nl & ({{7{PECore_DecodeAxiRead_case_4_switch_lp_nor_13_cse_1}},
      PECore_DecodeAxiRead_case_4_switch_lp_nor_13_cse_1}) & ({{7{PECore_DecodeAxiRead_switch_lp_nor_14_cse_1}},
      PECore_DecodeAxiRead_switch_lp_nor_14_cse_1});
  assign PEManager_16U_ClusterLookup_1_for_mux_58_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_9_sva_dfm_mx1[3:0])});
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_10_nl = MUX_v_8_2_2(pe_manager_cluster_lut_data_0_15_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_26_nl
      = PECore_DecodeAxiRead_case_4_switch_lp_mux_10_nl & ({{7{PECore_DecodeAxiRead_case_4_switch_lp_nor_13_cse_1}},
      PECore_DecodeAxiRead_case_4_switch_lp_nor_13_cse_1}) & ({{7{PECore_DecodeAxiRead_switch_lp_nor_14_cse_1}},
      PECore_DecodeAxiRead_switch_lp_nor_14_cse_1});
  assign PEManager_16U_ClusterLookup_1_for_mux_56_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_9_sva_dfm_mx1[7:4])});
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux1h_19_nl = MUX1HOT_v_8_4_2((pe_manager_base_input_0_sva[7:0]),
      pe_manager_cluster_lut_data_0_10_sva_dfm_4, (pe_manager_base_input_1_sva[7:0]),
      pe_manager_cluster_lut_data_1_10_sva_dfm_4, {PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5});
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_25_nl
      = PECore_DecodeAxiRead_case_4_switch_lp_mux1h_19_nl & ({{7{PECore_DecodeAxiRead_case_4_switch_lp_nor_12_cse_1}},
      PECore_DecodeAxiRead_case_4_switch_lp_nor_12_cse_1}) & ({{7{PECore_DecodeAxiRead_switch_lp_nor_14_cse_1}},
      PECore_DecodeAxiRead_switch_lp_nor_14_cse_1});
  assign PEManager_16U_ClusterLookup_1_for_mux_49_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_12_sva_dfm_mx1[3:0])});
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux1h_18_nl = MUX1HOT_v_8_4_2((pe_manager_base_input_0_sva[15:8]),
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, (pe_manager_base_input_1_sva[15:8]),
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, {PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5});
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl
      = PECore_DecodeAxiRead_case_4_switch_lp_mux1h_18_nl & ({{7{PECore_DecodeAxiRead_case_4_switch_lp_nor_12_cse_1}},
      PECore_DecodeAxiRead_case_4_switch_lp_nor_12_cse_1}) & ({{7{PECore_DecodeAxiRead_switch_lp_nor_14_cse_1}},
      PECore_DecodeAxiRead_switch_lp_nor_14_cse_1});
  assign PEManager_16U_ClusterLookup_1_for_mux_51_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_12_sva_dfm_mx1[7:4])});
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux1h_20_nl = MUX1HOT_v_8_4_2((pe_manager_base_bias_0_sva[7:0]),
      pe_manager_cluster_lut_data_0_8_sva_dfm_4, (pe_manager_base_bias_1_sva[7:0]),
      pe_manager_cluster_lut_data_1_8_sva_dfm_4, {PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5});
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl
      = PECore_DecodeAxiRead_case_4_switch_lp_mux1h_20_nl & ({{7{PECore_DecodeAxiRead_case_4_switch_lp_nor_12_cse_1}},
      PECore_DecodeAxiRead_case_4_switch_lp_nor_12_cse_1}) & ({{7{PECore_DecodeAxiRead_switch_lp_nor_14_cse_1}},
      PECore_DecodeAxiRead_switch_lp_nor_14_cse_1});
  assign PEManager_16U_ClusterLookup_1_for_mux_48_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_11_sva_dfm_mx1[7:4])});
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux1h_21_nl = MUX1HOT_v_8_4_2((pe_manager_base_bias_0_sva[15:8]),
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, (pe_manager_base_bias_1_sva[15:8]),
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, {PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5});
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl
      = PECore_DecodeAxiRead_case_4_switch_lp_mux1h_21_nl & ({{7{PECore_DecodeAxiRead_case_4_switch_lp_nor_12_cse_1}},
      PECore_DecodeAxiRead_case_4_switch_lp_nor_12_cse_1}) & ({{7{PECore_DecodeAxiRead_switch_lp_nor_14_cse_1}},
      PECore_DecodeAxiRead_switch_lp_nor_14_cse_1});
  assign PEManager_16U_ClusterLookup_for_mux_4_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_6_sva_dfm_mx1[3:0])});
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux1h_22_nl = MUX1HOT_v_8_4_2((pe_manager_base_weight_0_sva[7:0]),
      pe_manager_cluster_lut_data_0_6_sva_dfm_4, (pe_manager_base_weight_1_sva[7:0]),
      pe_manager_cluster_lut_data_1_6_sva_dfm_4, {PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5});
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl
      = PECore_DecodeAxiRead_case_4_switch_lp_mux1h_22_nl & ({{7{PECore_DecodeAxiRead_case_4_switch_lp_nor_12_cse_1}},
      PECore_DecodeAxiRead_case_4_switch_lp_nor_12_cse_1}) & ({{7{PECore_DecodeAxiRead_switch_lp_nor_14_cse_1}},
      PECore_DecodeAxiRead_switch_lp_nor_14_cse_1});
  assign PEManager_16U_ClusterLookup_1_for_mux_52_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_10_sva_dfm_mx1[7:4])});
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux1h_23_nl = MUX1HOT_v_8_4_2((pe_manager_base_weight_0_sva[15:8]),
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, (pe_manager_base_weight_1_sva[15:8]),
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, {PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5});
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_20_nl
      = PECore_DecodeAxiRead_case_4_switch_lp_mux1h_23_nl & ({{7{PECore_DecodeAxiRead_case_4_switch_lp_nor_12_cse_1}},
      PECore_DecodeAxiRead_case_4_switch_lp_nor_12_cse_1}) & ({{7{PECore_DecodeAxiRead_switch_lp_nor_14_cse_1}},
      PECore_DecodeAxiRead_switch_lp_nor_14_cse_1});
  assign PEManager_16U_ClusterLookup_1_for_mux_50_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_11_sva_dfm_mx1[3:0])});
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux1h_9_nl = MUX1HOT_v_8_3_2(pe_config_num_output_sva,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_1_5_sva_dfm_4,
      {PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_5 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5});
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_11_nl = ~(PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6
      | PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8 | PECore_DecodeAxiWrite_case_4_switch_lp_nor_tmp_1);
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_3_nl = PECore_DecodeAxiRead_case_4_switch_lp_mux1h_9_nl
      & (signext_8_1(PECore_DecodeAxiRead_case_4_switch_lp_nor_11_nl)) & ({{7{PECore_DecodeAxiRead_switch_lp_nor_14_cse_1}},
      PECore_DecodeAxiRead_switch_lp_nor_14_cse_1});
  assign PEManager_16U_ClusterLookup_1_for_mux_54_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_10_sva_dfm_mx1[3:0])});
  assign PECore_RunMac_nor_nl = ~(PECore_RunFSM_switch_lp_equal_tmp_5 | PECore_RunFSM_switch_lp_equal_tmp_4
      | PECore_RunMac_PECore_RunMac_and_2_cse);
  assign PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_32_nl
      = MUX_s_1_2_2(pe_manager_zero_active_0_sva, (rva_in_PopNB_mioi_idat_mxwt[0]),
      PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6);
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_34_nl
      = MUX_s_1_2_2(pe_manager_zero_active_0_sva, PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_32_nl,
      PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_31);
  assign PECore_DecodeAxi_if_mux_57_nl = MUX_s_1_2_2(pe_manager_zero_active_0_sva,
      PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_34_nl,
      rva_in_PopNB_mioi_idat_mxwt[168]);
  assign PECore_DecodeAxi_mux_127_nl = MUX_s_1_2_2(pe_manager_zero_active_0_sva,
      PECore_DecodeAxi_if_mux_57_nl, rva_in_PopNB_mioi_ivld_mxwt);
  assign pe_manager_zero_active_mux_nl = MUX_s_1_2_2(PECore_DecodeAxi_mux_127_nl,
      pe_manager_zero_active_0_sva, is_start_sva);
  assign PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_33_nl
      = MUX_s_1_2_2(pe_manager_zero_active_1_sva, (rva_in_PopNB_mioi_idat_mxwt[0]),
      PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8);
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_35_nl
      = MUX_s_1_2_2(pe_manager_zero_active_1_sva, PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_33_nl,
      PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_31);
  assign PECore_DecodeAxi_if_mux_55_nl = MUX_s_1_2_2(pe_manager_zero_active_1_sva,
      PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_35_nl,
      rva_in_PopNB_mioi_idat_mxwt[168]);
  assign PECore_DecodeAxi_mux_125_nl = MUX_s_1_2_2(pe_manager_zero_active_1_sva,
      PECore_DecodeAxi_if_mux_55_nl, rva_in_PopNB_mioi_ivld_mxwt);
  assign pe_manager_zero_active_mux_1_nl = MUX_s_1_2_2(PECore_DecodeAxi_mux_125_nl,
      pe_manager_zero_active_1_sva, is_start_sva);
  assign PECore_UpdateFSM_case_1_if_mux_nl = MUX_s_1_2_2(pe_manager_zero_active_mux_nl,
      pe_manager_zero_active_mux_1_nl, pe_config_manager_counter_sva_dfm_4_mx0_0);
  assign PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl = pe_config_is_zero_first_sva_dfm_4_mx0
      & PECore_UpdateFSM_case_1_if_mux_nl;
  assign PEManager_16U_ClusterLookup_for_mux_145_nl = MUX_v_5_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[4:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_0_sva_dfm_mx1[7:4])});
  assign nl_PECore_RunBias_if_for_3_operator_33_true_acc_nl = (operator_4_false_acc_psp_3_sva_1[3:1])
      + 3'b111;
  assign PECore_RunBias_if_for_3_operator_33_true_acc_nl = nl_PECore_RunBias_if_for_3_operator_33_true_acc_nl[2:0];
  assign nl_PECore_RunBias_if_for_3_operator_34_true_acc_nl = conv_s2s_4_5({PECore_RunBias_if_for_3_operator_33_true_acc_nl
      , (operator_4_false_acc_psp_3_sva_1[0])}) + 5'b00111;
  assign PECore_RunBias_if_for_3_operator_34_true_acc_nl = nl_PECore_RunBias_if_for_3_operator_34_true_acc_nl[4:0];
  assign PEManager_16U_ClusterLookup_for_mux_144_nl = MUX_v_5_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[4:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_5_sva_dfm_mx1[3:0])});
  assign nl_PECore_RunBias_if_for_4_operator_33_true_acc_nl = (operator_4_false_acc_psp_4_sva_1[3:1])
      + 3'b111;
  assign PECore_RunBias_if_for_4_operator_33_true_acc_nl = nl_PECore_RunBias_if_for_4_operator_33_true_acc_nl[2:0];
  assign nl_PECore_RunBias_if_for_4_operator_34_true_acc_nl = conv_s2s_4_5({PECore_RunBias_if_for_4_operator_33_true_acc_nl
      , (operator_4_false_acc_psp_4_sva_1[0])}) + 5'b00111;
  assign PECore_RunBias_if_for_4_operator_34_true_acc_nl = nl_PECore_RunBias_if_for_4_operator_34_true_acc_nl[4:0];
  assign PEManager_16U_ClusterLookup_for_mux_46_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_0_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_44_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_0_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_42_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_1_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_40_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_1_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_38_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_2_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_36_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_2_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_34_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_3_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_32_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_3_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_33_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_4_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_35_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_4_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_37_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_5_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_39_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_5_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_41_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_6_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_43_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_6_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_45_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_7_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_47_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_2_7_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_30_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_8_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_28_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_8_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_26_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_9_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_24_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_9_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_22_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_10_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_20_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_10_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_18_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_11_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_16_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_11_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_17_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_12_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_19_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_12_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_21_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_13_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_23_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_13_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_25_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_14_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_27_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_14_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_29_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_15_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_31_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_15_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_30_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_0_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_28_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_0_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_26_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_1_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_24_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_1_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_22_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_2_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_20_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_2_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_18_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_3_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_16_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_3_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_17_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_4_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_19_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_4_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_21_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_5_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_23_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_5_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_25_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_6_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_27_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_6_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_29_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_7_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_31_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_1_7_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_131_nl = MUX_v_4_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[3:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_14_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_130_nl = MUX_v_4_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[3:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_14_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_129_nl = MUX_v_4_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[3:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_15_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_128_nl = MUX_v_4_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[3:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_15_sva_dfm_mx1[7:4])});
  assign weight_mem_run_1_for_5_mux_30_nl = MUX_v_8_2_2(weight_port_read_out_data_11_0_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm);
  assign PEManager_16U_ClusterLookup_1_for_mux_94_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_8_sva_dfm_mx1[3:0])});
  assign weight_mem_run_1_for_5_mux_31_nl = MUX_v_8_2_2(weight_port_read_out_data_11_1_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm);
  assign PEManager_16U_ClusterLookup_1_for_mux_92_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_8_sva_dfm_mx1[7:4])});
  assign weight_mem_run_1_for_5_mux_32_nl = MUX_v_8_2_2(weight_port_read_out_data_11_2_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm);
  assign PEManager_16U_ClusterLookup_1_for_mux_90_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_9_sva_dfm_mx1[3:0])});
  assign weight_mem_run_1_for_5_mux_33_nl = MUX_v_8_2_2(weight_port_read_out_data_11_3_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm);
  assign PEManager_16U_ClusterLookup_1_for_mux_88_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_9_sva_dfm_mx1[7:4])});
  assign weight_mem_run_1_for_5_mux_34_nl = MUX_v_8_2_2(weight_port_read_out_data_11_4_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm);
  assign PEManager_16U_ClusterLookup_1_for_mux_86_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_10_sva_dfm_mx1[3:0])});
  assign weight_mem_run_1_for_5_mux_35_nl = MUX_v_8_2_2(weight_port_read_out_data_11_5_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm);
  assign PEManager_16U_ClusterLookup_1_for_mux_84_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_10_sva_dfm_mx1[7:4])});
  assign weight_mem_run_1_for_5_mux_36_nl = MUX_v_8_2_2(weight_port_read_out_data_11_6_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm);
  assign PEManager_16U_ClusterLookup_1_for_mux_82_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_11_sva_dfm_mx1[3:0])});
  assign weight_mem_run_1_for_5_mux_37_nl = MUX_v_8_2_2(weight_port_read_out_data_11_7_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm);
  assign PEManager_16U_ClusterLookup_1_for_mux_80_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_11_sva_dfm_mx1[7:4])});
  assign weight_mem_run_1_for_5_mux_38_nl = MUX_v_8_2_2(weight_port_read_out_data_11_8_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm);
  assign PEManager_16U_ClusterLookup_1_for_mux_81_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_12_sva_dfm_mx1[3:0])});
  assign weight_mem_run_1_for_5_mux_39_nl = MUX_v_8_2_2(weight_port_read_out_data_11_9_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm);
  assign PEManager_16U_ClusterLookup_1_for_mux_83_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_12_sva_dfm_mx1[7:4])});
  assign weight_mem_run_1_for_5_mux_40_nl = MUX_v_8_2_2(weight_port_read_out_data_11_10_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm);
  assign PEManager_16U_ClusterLookup_1_for_mux_85_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_13_sva_dfm_mx1[3:0])});
  assign weight_mem_run_1_for_5_mux_41_nl = MUX_v_8_2_2(weight_port_read_out_data_11_11_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm);
  assign PEManager_16U_ClusterLookup_1_for_mux_87_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_13_sva_dfm_mx1[7:4])});
  assign weight_mem_run_1_for_5_mux_42_nl = MUX_v_8_2_2(weight_port_read_out_data_11_12_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm);
  assign PEManager_16U_ClusterLookup_1_for_mux_89_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_14_sva_dfm_mx1[3:0])});
  assign weight_mem_run_1_for_5_mux_43_nl = MUX_v_8_2_2(weight_port_read_out_data_11_13_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm);
  assign PEManager_16U_ClusterLookup_1_for_mux_91_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_14_sva_dfm_mx1[7:4])});
  assign weight_mem_run_1_for_5_mux_44_nl = MUX_v_8_2_2(weight_port_read_out_data_11_14_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm);
  assign PEManager_16U_ClusterLookup_1_for_mux_93_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_15_sva_dfm_mx1[3:0])});
  assign data_in_tmp_operator_for_mux_34_nl = MUX_v_8_2_2(weight_port_read_out_data_11_15_sva_dfm,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1,
      crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm);
  assign PEManager_16U_ClusterLookup_1_for_mux_95_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_5_15_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_8_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_1_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_8_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_2_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_9_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_3_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_9_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_4_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_10_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_5_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_10_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_6_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_11_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_7_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_11_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_8_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_12_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_9_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_12_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_10_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_13_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_11_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_13_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_12_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_14_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_13_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_14_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_14_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_15_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_1_for_mux_15_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_15_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_0_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_14_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_1_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_13_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_1_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_12_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_2_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_11_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_2_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_10_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_3_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_9_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_3_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_8_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_4_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_7_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_4_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_for_mux_1_nl = MUX_v_8_32_2(pe_manager_cluster_lut_data_0_0_sva_dfm_4,
      pe_manager_cluster_lut_data_0_1_sva_dfm_4, pe_manager_cluster_lut_data_0_2_sva_dfm_4,
      pe_manager_cluster_lut_data_0_3_sva_dfm_4, pe_manager_cluster_lut_data_0_4_sva_dfm_4,
      pe_manager_cluster_lut_data_0_5_sva_dfm_4, pe_manager_cluster_lut_data_0_6_sva_dfm_4,
      pe_manager_cluster_lut_data_0_7_sva_dfm_4, pe_manager_cluster_lut_data_0_8_sva_dfm_4,
      pe_manager_cluster_lut_data_0_9_sva_dfm_4, pe_manager_cluster_lut_data_0_10_sva_dfm_4,
      pe_manager_cluster_lut_data_0_11_sva_dfm_4, pe_manager_cluster_lut_data_0_12_sva_dfm_4,
      pe_manager_cluster_lut_data_0_13_sva_dfm_4, pe_manager_cluster_lut_data_0_14_sva_dfm_4,
      pe_manager_cluster_lut_data_0_15_sva_dfm_4, pe_manager_cluster_lut_data_1_0_sva_dfm_4,
      pe_manager_cluster_lut_data_1_1_sva_dfm_4, pe_manager_cluster_lut_data_1_2_sva_dfm_4,
      pe_manager_cluster_lut_data_1_3_sva_dfm_4, pe_manager_cluster_lut_data_1_4_sva_dfm_4,
      pe_manager_cluster_lut_data_1_5_sva_dfm_4, pe_manager_cluster_lut_data_1_6_sva_dfm_4,
      pe_manager_cluster_lut_data_1_7_sva_dfm_4, pe_manager_cluster_lut_data_1_8_sva_dfm_4,
      pe_manager_cluster_lut_data_1_9_sva_dfm_4, pe_manager_cluster_lut_data_1_10_sva_dfm_4,
      pe_manager_cluster_lut_data_1_11_sva_dfm_4, pe_manager_cluster_lut_data_1_12_sva_dfm_4,
      pe_manager_cluster_lut_data_1_13_sva_dfm_4, pe_manager_cluster_lut_data_1_14_sva_dfm_4,
      pe_manager_cluster_lut_data_1_15_sva_dfm_4, {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_7_sva_dfm_mx1[7:4])});
  assign PEManager_16U_ClusterLookup_1_for_mux_133_nl = MUX_v_4_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[3:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_13_sva_dfm_mx1[3:0])});
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux1h_5_nl = MUX1HOT_v_4_5_2(pe_config_num_manager_sva,
      (pe_manager_num_input_0_sva[3:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[3:0]),
      (pe_manager_num_input_1_sva[3:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[3:0]),
      {PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_5 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5});
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_1_nl = PECore_DecodeAxiRead_case_4_switch_lp_mux1h_5_nl
      & (signext_4_1(~ PECore_DecodeAxiWrite_case_4_switch_lp_nor_tmp_1)) & ({{3{PECore_DecodeAxiRead_switch_lp_nor_14_cse_1}},
      PECore_DecodeAxiRead_switch_lp_nor_14_cse_1});
  assign PEManager_16U_ClusterLookup_1_for_mux_132_nl = MUX_v_4_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[3:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_3_13_sva_dfm_mx1[7:4])});
  assign and_5134_nl = (or_dcpl_34 | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_14
      | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_6 | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_10
      | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_2 | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_4
      | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_0 | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_9
      | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_1 | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_8
      | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_7 | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_3
      | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_11 | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_5
      | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_12 | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_13)
      & (~ crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_tmp) & weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_224_tmp
      & (fsm_output[1]);
  assign and_5136_nl = (((weight_mem_write_arbxbar_xbar_for_lshift_tmp[15]) & weight_mem_read_arbxbar_xbar_for_3_16_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp
      & (~ Arbiter_16U_Roundrobin_pick_mux_2460_tmp_14) & (~(Arbiter_16U_Roundrobin_pick_mux_2460_tmp_6
      | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_10)) & (~(Arbiter_16U_Roundrobin_pick_mux_2460_tmp_2
      | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_4)) & (~(Arbiter_16U_Roundrobin_pick_mux_2460_tmp_0
      | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_9)) & (~(Arbiter_16U_Roundrobin_pick_mux_2460_tmp_1
      | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_8)) & (~(Arbiter_16U_Roundrobin_pick_mux_2460_tmp_7
      | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_3)) & (~(Arbiter_16U_Roundrobin_pick_mux_2460_tmp_11
      | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_5)) & (~(Arbiter_16U_Roundrobin_pick_mux_2460_tmp_12
      | Arbiter_16U_Roundrobin_pick_mux_2460_tmp_13))) | crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_tmp
      | (~ weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_224_tmp)) & (fsm_output[1]);
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_and_1_nl = PECore_PushAxiRsp_if_asn_68
      & PECore_RunBias_if_for_and_42_cse;
  assign crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_and_2_nl = crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm
      & PECore_RunBias_if_for_and_42_cse;
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux1h_10_nl = MUX1HOT_v_2_4_2((pe_manager_adplfloat_bias_weight_0_sva[2:1]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[2:1]), (pe_manager_adplfloat_bias_weight_1_sva[2:1]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[2:1]), {PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5});
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_9_nl = MUX_v_2_2_2(2'b00, PECore_DecodeAxiRead_case_4_switch_lp_mux1h_10_nl,
      PECore_DecodeAxiRead_case_4_switch_lp_nor_12_cse_1);
  assign PEManager_16U_ClusterLookup_for_mux_135_nl = MUX_v_2_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[1:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_4_sva_dfm_mx1[7:4])});
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux1h_4_nl = MUX1HOT_v_2_4_2((pe_manager_adplfloat_bias_bias_0_sva[2:1]),
      (pe_manager_cluster_lut_data_0_2_sva_dfm_4[2:1]), (pe_manager_adplfloat_bias_bias_1_sva[2:1]),
      (pe_manager_cluster_lut_data_1_2_sva_dfm_4[2:1]), {PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5});
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_7_nl = MUX_v_2_2_2(2'b00, PECore_DecodeAxiRead_case_4_switch_lp_mux1h_4_nl,
      PECore_DecodeAxiRead_case_4_switch_lp_nor_12_cse_1);
  assign PEManager_16U_ClusterLookup_for_mux_133_nl = MUX_v_2_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[1:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_5_sva_dfm_mx1[7:4])});
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux1h_1_nl = MUX1HOT_v_2_4_2((pe_manager_adplfloat_bias_input_0_sva[2:1]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[2:1]), (pe_manager_adplfloat_bias_input_1_sva[2:1]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[2:1]), {PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5});
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_6_nl = MUX_v_2_2_2(2'b00, PECore_DecodeAxiRead_case_4_switch_lp_mux1h_1_nl,
      PECore_DecodeAxiRead_case_4_switch_lp_nor_12_cse_1);
  assign PEManager_16U_ClusterLookup_for_mux_131_nl = MUX_v_2_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[1:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[1:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[1:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_6_sva_dfm_mx1[3:0])});
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl = MUX_v_7_2_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[7:1]),
      (pe_manager_cluster_lut_data_1_0_sva_dfm_4[7:1]), PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5);
  assign PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_13_nl
      = MUX_v_7_2_2(7'b0000000, PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl, PECore_DecodeAxiRead_case_4_switch_lp_nor_13_cse_1);
  assign PEManager_16U_ClusterLookup_for_mux_128_nl = MUX_v_7_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[6:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[6:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[6:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[6:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[6:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[6:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[6:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[6:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[6:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[6:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[6:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[6:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[6:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[6:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[6:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[6:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[6:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[6:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[6:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[6:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[6:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[6:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[6:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[6:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[6:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[6:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[6:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[6:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[6:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[6:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[6:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[6:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_7_sva_dfm_mx1[7:4])});
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_2_nl = MUX_v_5_2_2((pe_manager_cluster_lut_data_0_1_sva_dfm_4[7:3]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[7:3]), PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5);
  assign PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_12_nl
      = MUX_v_5_2_2(5'b00000, PECore_DecodeAxiRead_case_4_switch_lp_mux_2_nl, PECore_DecodeAxiRead_case_4_switch_lp_nor_13_cse_1);
  assign nl_PECore_RunBias_if_for_12_operator_33_true_acc_nl = (operator_4_false_acc_psp_12_sva_1[3:1])
      + 3'b111;
  assign PECore_RunBias_if_for_12_operator_33_true_acc_nl = nl_PECore_RunBias_if_for_12_operator_33_true_acc_nl[2:0];
  assign nl_PECore_RunBias_if_for_12_operator_34_true_acc_nl = conv_s2s_4_5({PECore_RunBias_if_for_12_operator_33_true_acc_nl
      , (operator_4_false_acc_psp_12_sva_1[0])}) + 5'b00111;
  assign PECore_RunBias_if_for_12_operator_34_true_acc_nl = nl_PECore_RunBias_if_for_12_operator_34_true_acc_nl[4:0];
  assign PEManager_16U_ClusterLookup_for_mux_134_nl = MUX_v_5_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[4:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_5_sva_dfm_mx1[3:0])});
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_nl = MUX_v_5_2_2((pe_manager_cluster_lut_data_0_2_sva_dfm_4[7:3]),
      (pe_manager_cluster_lut_data_1_2_sva_dfm_4[7:3]), PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5);
  assign PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_10_nl
      = MUX_v_5_2_2(5'b00000, PECore_DecodeAxiRead_case_4_switch_lp_mux_nl, PECore_DecodeAxiRead_case_4_switch_lp_nor_13_cse_1);
  assign PEManager_16U_ClusterLookup_for_mux_132_nl = MUX_v_5_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[4:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_0_7_sva_dfm_mx1[3:0])});
  assign PEManager_16U_ClusterLookup_for_mux_130_nl = MUX_v_5_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[4:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[4:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[4:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_6_sva_dfm_mx1[7:4])});
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_1_nl = MUX_v_5_2_2((pe_manager_cluster_lut_data_0_3_sva_dfm_4[7:3]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[7:3]), PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5);
  assign PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_11_nl
      = MUX_v_5_2_2(5'b00000, PECore_DecodeAxiRead_case_4_switch_lp_mux_1_nl, PECore_DecodeAxiRead_case_4_switch_lp_nor_13_cse_1);
  assign nl_PECore_RunBias_if_for_2_operator_33_true_acc_nl = (operator_4_false_acc_psp_2_sva_1[3:1])
      + 3'b111;
  assign PECore_RunBias_if_for_2_operator_33_true_acc_nl = nl_PECore_RunBias_if_for_2_operator_33_true_acc_nl[2:0];
  assign nl_PECore_RunBias_if_for_2_operator_34_true_acc_nl = conv_s2s_4_5({PECore_RunBias_if_for_2_operator_33_true_acc_nl
      , (operator_4_false_acc_psp_2_sva_1[0])}) + 5'b00111;
  assign PECore_RunBias_if_for_2_operator_34_true_acc_nl = nl_PECore_RunBias_if_for_2_operator_34_true_acc_nl[4:0];
  assign PECore_RunMac_if_and_803_nl = PECore_RunBias_if_for_and_45_rgt & (or_dcpl_247
      | or_3399_cse);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux1h_24_nl = MUX1HOT_v_4_4_2((pe_manager_num_input_0_sva[7:4]),
      (pe_manager_cluster_lut_data_0_4_sva_dfm_4[7:4]), (pe_manager_num_input_1_sva[7:4]),
      (pe_manager_cluster_lut_data_1_4_sva_dfm_4[7:4]), {PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7 , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8
      , PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5});
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl
      = PECore_DecodeAxiRead_case_4_switch_lp_mux1h_24_nl & ({{3{PECore_DecodeAxiRead_case_4_switch_lp_nor_12_cse_1}},
      PECore_DecodeAxiRead_case_4_switch_lp_nor_12_cse_1}) & ({{3{PECore_DecodeAxiRead_switch_lp_nor_14_cse_1}},
      PECore_DecodeAxiRead_switch_lp_nor_14_cse_1});
  assign PEManager_16U_ClusterLookup_for_mux_129_nl = MUX_v_4_32_2((pe_manager_cluster_lut_data_0_0_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_1_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_2_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_3_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_4_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_5_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_6_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_7_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_8_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_9_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_10_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_11_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_12_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_13_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_0_14_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_0_15_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_0_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_1_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_2_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_3_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_4_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_5_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_6_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_7_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_8_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_9_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_10_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_11_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_12_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_13_sva_dfm_4[3:0]), (pe_manager_cluster_lut_data_1_14_sva_dfm_4[3:0]),
      (pe_manager_cluster_lut_data_1_15_sva_dfm_4[3:0]), {(reg_PECore_RunMac_if_mux_142_ftd_1[0])
      , (weight_port_read_out_data_4_7_sva_dfm_mx1[3:0])});
  assign rva_out_reg_data_and_1_nl = PECore_PushAxiRsp_if_asn_68 & (fsm_output[2])
      & PECore_RunMac_if_nand_56_rgt;
  assign PECore_RunMac_if_and_801_nl = rva_out_reg_data_and_2_cse & PECore_RunMac_if_nand_56_rgt;
  assign nl_PECore_RunBias_if_for_1_operator_33_true_acc_1_nl = (operator_4_false_acc_psp_1_sva_1[3:1])
      + 3'b111;
  assign PECore_RunBias_if_for_1_operator_33_true_acc_1_nl = nl_PECore_RunBias_if_for_1_operator_33_true_acc_1_nl[2:0];
  assign operator_4_false_mux_2_nl = MUX_v_4_2_2(pe_config_manager_counter_sva_dfm_4_mx1,
      ({PECore_RunBias_if_for_1_operator_33_true_acc_1_nl , (operator_4_false_acc_psp_1_sva_1[0])}),
      fsm_output[2]);
  assign nl_z_out_4 = conv_s2u_4_5(operator_4_false_mux_2_nl) + conv_u2u_3_5(signext_3_2({(fsm_output[2])
      , 1'b1}));
  assign z_out_4 = nl_z_out_4[4:0];
  assign and_5952_nl = state_2_0_sva_2 & (fsm_output[1]);
  assign operator_8_false_mux_2_nl = MUX_v_8_2_2(pe_config_input_counter_sva_dfm_4_mx0,
      pe_config_output_counter_sva_dfm_4_mx0, and_5952_nl);
  assign nl_z_out_5 = operator_8_false_mux_2_nl + 8'b00000001;
  assign z_out_5 = nl_z_out_5[7:0];
  assign operator_16_false_1_mux_16_cse = MUX_v_16_2_2(({PEManager_16U_GetWeightAddr_1_else_acc_2_psp_sva_1
      , (PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx1[3:0])}),
      ({PEManager_16U_GetWeightAddr_if_acc_2_psp_sva_1 , (PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx0_3_0[2:0])}),
      and_5541_cse);
  assign operator_32_true_mux1h_40_nl = MUX1HOT_v_13_3_2((~ (PECore_RunBias_if_accum_vector_out_data_11_lpi_1_dfm_mx2[31:19])),
      (~ (PECore_RunBias_if_accum_vector_out_data_mux_11_cse[31:19])), (~ (PECore_RunBias_if_accum_vector_out_data_mux_5_cse[31:19])),
      {(fsm_output[1]) , (fsm_output[2]) , or_dcpl_251});
  assign nl_operator_32_true_acc_nl = conv_s2u_13_14(operator_32_true_mux1h_40_nl)
      + 14'b00000000000001;
  assign operator_32_true_acc_nl = nl_operator_32_true_acc_nl[13:0];
  assign z_out_10_13 = readslicef_14_1_13(operator_32_true_acc_nl);
  assign operator_32_true_mux1h_41_nl = MUX1HOT_v_13_3_2((~ (PECore_RunBias_if_accum_vector_out_data_10_lpi_1_dfm_mx2[31:19])),
      (~ (PECore_RunBias_if_accum_vector_out_data_mux_9_cse[31:19])), (~ (PECore_RunBias_if_accum_vector_out_data_mux_7_cse[31:19])),
      {(fsm_output[1]) , (fsm_output[2]) , or_dcpl_251});
  assign nl_operator_32_true_acc_1_nl = conv_s2u_13_14(operator_32_true_mux1h_41_nl)
      + 14'b00000000000001;
  assign operator_32_true_acc_1_nl = nl_operator_32_true_acc_1_nl[13:0];
  assign z_out_11_13 = readslicef_14_1_13(operator_32_true_acc_1_nl);
  assign operator_32_true_mux1h_42_nl = MUX1HOT_v_13_4_2((~ (PECore_RunBias_if_accum_vector_out_data_7_lpi_1_dfm_mx2[31:19])),
      (~ (PECore_RunBias_if_accum_vector_out_data_mux_7_cse[31:19])), (~ (PECore_RunBias_if_accum_vector_out_data_mux_11_cse[31:19])),
      (~ (PECore_RunBias_if_accum_vector_out_data_mux_9_cse[31:19])), {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])});
  assign nl_operator_32_true_acc_2_nl = conv_s2u_13_14(operator_32_true_mux1h_42_nl)
      + 14'b00000000000001;
  assign operator_32_true_acc_2_nl = nl_operator_32_true_acc_2_nl[13:0];
  assign z_out_12_13 = readslicef_14_1_13(operator_32_true_acc_2_nl);
  assign operator_32_true_mux1h_43_nl = MUX1HOT_v_13_4_2((~ (PECore_RunBias_if_accum_vector_out_data_6_lpi_1_dfm_mx2[31:19])),
      (~ (PECore_RunBias_if_accum_vector_out_data_mux_5_cse[31:19])), (~ (PECore_RunBias_if_accum_vector_out_data_mux_9_cse[31:19])),
      (~ (PECore_RunBias_if_accum_vector_out_data_mux_11_cse[31:19])), {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])});
  assign nl_operator_32_true_acc_3_nl = conv_s2u_13_14(operator_32_true_mux1h_43_nl)
      + 14'b00000000000001;
  assign operator_32_true_acc_3_nl = nl_operator_32_true_acc_3_nl[13:0];
  assign z_out_13_13 = readslicef_14_1_13(operator_32_true_acc_3_nl);
  assign adpfloat_tmp_to_fixed_20U_14U_if_1_adpfloat_tmp_to_fixed_20U_14U_if_1_mux_2_nl
      = MUX_v_20_2_2((~ z_out_46), (~ z_out_49), fsm_output[1]);
  assign nl_z_out_17 = adpfloat_tmp_to_fixed_20U_14U_if_1_adpfloat_tmp_to_fixed_20U_14U_if_1_mux_2_nl
      + 20'b00000000000000000001;
  assign z_out_17 = nl_z_out_17[19:0];
  assign adpfloat_tmp_to_fixed_20U_14U_if_1_mux1h_8_nl = MUX1HOT_v_20_3_2((~ z_out_49),
      (~ z_out_47), (~ z_out_48), {(fsm_output[2]) , or_dcpl_251 , (fsm_output[1])});
  assign nl_z_out_18 = adpfloat_tmp_to_fixed_20U_14U_if_1_mux1h_8_nl + 20'b00000000000000000001;
  assign z_out_18 = nl_z_out_18[19:0];
  assign adpfloat_tmp_to_fixed_20U_14U_if_1_adpfloat_tmp_to_fixed_20U_14U_if_1_mux_3_nl
      = MUX_v_20_2_2((~ z_out_48), (~ z_out_47), fsm_output[1]);
  assign nl_z_out_19 = adpfloat_tmp_to_fixed_20U_14U_if_1_adpfloat_tmp_to_fixed_20U_14U_if_1_mux_3_nl
      + 20'b00000000000000000001;
  assign z_out_19 = nl_z_out_19[19:0];
  assign adpfloat_tmp_to_fixed_20U_14U_if_1_mux1h_9_nl = MUX1HOT_v_20_3_2((~ z_out_47),
      (~ z_out_49), (~ z_out_46), {(fsm_output[2]) , or_dcpl_251 , (fsm_output[1])});
  assign nl_z_out_20 = adpfloat_tmp_to_fixed_20U_14U_if_1_mux1h_9_nl + 20'b00000000000000000001;
  assign z_out_20 = nl_z_out_20[19:0];
  assign operator_32_true_mux1h_8_nl = MUX1HOT_v_32_3_2(PECore_RunBias_if_accum_vector_out_data_6_lpi_1_dfm_mx2,
      PECore_RunBias_if_accum_vector_out_data_mux_5_cse, PECore_RunBias_if_accum_vector_out_data_mux_9_cse,
      {(fsm_output[1]) , and_4616_cse , (fsm_output[4])});
  assign nl_operator_32_true_acc_nl_1 = conv_s2u_32_33(operator_32_true_mux1h_8_nl)
      + 33'b000000000000001111111111111111111;
  assign operator_32_true_acc_nl_1 = nl_operator_32_true_acc_nl_1[32:0];
  assign z_out_21_32 = readslicef_33_1_32(operator_32_true_acc_nl_1);
  assign operator_32_true_mux1h_9_nl = MUX1HOT_v_32_3_2(PECore_RunBias_if_accum_vector_out_data_7_lpi_1_dfm_mx2,
      PECore_RunBias_if_accum_vector_out_data_mux_11_cse, PECore_RunBias_if_accum_vector_out_data_mux_7_cse,
      {(fsm_output[1]) , and_4616_cse , (fsm_output[4])});
  assign nl_operator_32_true_acc_1_nl_1 = conv_s2u_32_33(operator_32_true_mux1h_9_nl)
      + 33'b000000000000001111111111111111111;
  assign operator_32_true_acc_1_nl_1 = nl_operator_32_true_acc_1_nl_1[32:0];
  assign z_out_22_32 = readslicef_33_1_32(operator_32_true_acc_1_nl_1);
  assign operator_32_true_mux1h_10_nl = MUX1HOT_v_32_3_2(PECore_RunBias_if_accum_vector_out_data_10_lpi_1_dfm_mx2,
      PECore_RunBias_if_accum_vector_out_data_mux_9_cse, PECore_RunBias_if_accum_vector_out_data_mux_5_cse,
      {(fsm_output[1]) , and_4616_cse , (fsm_output[4])});
  assign nl_operator_32_true_acc_2_nl_1 = conv_s2u_32_33(operator_32_true_mux1h_10_nl)
      + 33'b000000000000001111111111111111111;
  assign operator_32_true_acc_2_nl_1 = nl_operator_32_true_acc_2_nl_1[32:0];
  assign z_out_23_32 = readslicef_33_1_32(operator_32_true_acc_2_nl_1);
  assign operator_32_true_mux1h_11_nl = MUX1HOT_v_32_3_2(PECore_RunBias_if_accum_vector_out_data_11_lpi_1_dfm_mx2,
      PECore_RunBias_if_accum_vector_out_data_mux_7_cse, PECore_RunBias_if_accum_vector_out_data_mux_11_cse,
      {(fsm_output[1]) , and_4616_cse , (fsm_output[4])});
  assign nl_operator_32_true_acc_3_nl_1 = conv_s2u_32_33(operator_32_true_mux1h_11_nl)
      + 33'b000000000000001111111111111111111;
  assign operator_32_true_acc_3_nl_1 = nl_operator_32_true_acc_3_nl_1[32:0];
  assign z_out_24_32 = readslicef_33_1_32(operator_32_true_acc_3_nl_1);
  assign PECore_RunMac_if_for_mux1h_4_nl = MUX1HOT_v_32_4_2(accum_vector_data_4_sva,
      accum_vector_data_13_sva, accum_vector_data_5_sva, PECore_RunBias_if_accum_vector_out_data_lpi_1_dfm,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[2]) , (fsm_output[4])});
  assign nl_z_out_25 = PECore_RunMac_if_for_mux1h_4_nl + Datapath_for_1_ProductSum_cmp_1_out_rsc_z;
  assign z_out_25 = nl_z_out_25[31:0];
  assign PECore_RunMac_if_for_mux1h_5_nl = MUX1HOT_v_32_4_2(accum_vector_data_3_sva,
      accum_vector_data_14_sva, accum_vector_data_8_sva, accum_vector_data_6_sva,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[2])});
  assign nl_z_out_26 = PECore_RunMac_if_for_mux1h_5_nl + Datapath_for_1_ProductSum_cmp_2_out_rsc_z;
  assign z_out_26 = nl_z_out_26[31:0];
  assign PECore_RunMac_if_for_mux1h_6_nl = MUX1HOT_v_32_4_2(accum_vector_data_2_sva,
      accum_vector_data_12_sva, accum_vector_data_7_sva, accum_vector_data_9_sva,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[2])});
  assign nl_z_out_27 = PECore_RunMac_if_for_mux1h_6_nl + Datapath_for_1_ProductSum_cmp_3_out_rsc_z;
  assign z_out_27 = nl_z_out_27[31:0];
  assign PECore_RunMac_if_for_mux1h_7_nl = MUX1HOT_v_32_4_2(accum_vector_data_15_sva,
      PECore_RunBias_if_accum_vector_out_data_13_lpi_1_dfm, PECore_RunBias_if_accum_vector_out_data_14_lpi_1_dfm,
      PECore_RunBias_if_accum_vector_out_data_15_lpi_1_dfm, {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[1]) , (fsm_output[2])});
  assign nl_z_out_28 = PECore_RunMac_if_for_mux1h_7_nl + Datapath_for_1_ProductSum_cmp_out_rsc_z;
  assign z_out_28 = nl_z_out_28[31:0];
  assign adpfloat_tmp_to_fixed_20U_14U_mux1h_28_tmp = MUX1HOT_s_1_3_2((input_mem_banks_write_if_for_if_mux_cse[103]),
      (input_mem_banks_read_read_data_lpi_1[7]), (input_mem_banks_read_read_data_lpi_1[15]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])});
  assign or_3880_tmp = ((~ PECore_DecodeAxiRead_switch_lp_nor_tmp) & (fsm_output[3]))
      | (((input_mem_banks_write_if_for_if_mux_cse[102:96]!=7'b0000000)) & (fsm_output[2]))
      | ((~ PECore_RunBias_if_for_13_operator_32_true_slc_operator_32_true_acc_13_svs)
      & (fsm_output[4]));
  assign PECore_RunBias_if_for_if_and_8_nl = (~(adpfloat_tmp_is_zero_land_10_lpi_1_dfm_st
      | (input_mem_banks_read_read_data_lpi_1[79]))) & (fsm_output[1]);
  assign adpfloat_tmp_to_fixed_20U_14U_and_8_nl = adpfloat_tmp_is_zero_land_10_lpi_1_dfm_st
      & (~ (input_mem_banks_read_read_data_lpi_1[79])) & (fsm_output[1]);
  assign PECore_RunBias_if_for_if_mux1h_4_nl = MUX1HOT_v_20_3_2(z_out_48, act_port_reg_data_asn_1_itm,
      z_out_18, {PECore_RunBias_if_for_if_and_8_nl , adpfloat_tmp_to_fixed_20U_14U_and_8_nl
      , (input_mem_banks_read_read_data_lpi_1[79])});
  assign PECore_RunBias_if_for_if_or_9_nl = (fsm_output[4:2]!=3'b000);
  assign PECore_RunBias_if_for_if_or_8_nl = MUX_v_20_2_2(PECore_RunBias_if_for_if_mux1h_4_nl,
      20'b11111111111111111111, PECore_RunBias_if_for_if_or_9_nl);
  assign adpfloat_tmp_to_fixed_20U_14U_and_nl = (~ (fsm_output[4])) & (~ adpfloat_tmp_to_fixed_20U_14U_mux1h_28_tmp)
      & or_3880_tmp;
  assign adpfloat_tmp_to_fixed_20U_14U_and_12_nl = (fsm_output[4]) & (~ adpfloat_tmp_to_fixed_20U_14U_mux1h_28_tmp)
      & or_3880_tmp;
  assign adpfloat_tmp_to_fixed_20U_14U_and_13_nl = (~ (fsm_output[4])) & adpfloat_tmp_to_fixed_20U_14U_mux1h_28_tmp
      & or_3880_tmp;
  assign adpfloat_tmp_to_fixed_20U_14U_and_14_nl = (fsm_output[4]) & adpfloat_tmp_to_fixed_20U_14U_mux1h_28_tmp
      & or_3880_tmp;
  assign mux1h_16_nl = MUX1HOT_v_20_5_2(PECore_RunBias_if_for_if_or_8_nl, z_out_46,
      z_out_47, z_out_17, z_out_18, {(~ or_3880_tmp) , adpfloat_tmp_to_fixed_20U_14U_and_nl
      , adpfloat_tmp_to_fixed_20U_14U_and_12_nl , adpfloat_tmp_to_fixed_20U_14U_and_13_nl
      , adpfloat_tmp_to_fixed_20U_14U_and_14_nl});
  assign nor_599_nl = ~((PECore_DecodeAxiRead_switch_lp_nor_tmp & (fsm_output[3]))
      | (adpfloat_tmp_is_zero_land_10_lpi_1_dfm & (fsm_output[1])) | ((input_mem_banks_write_if_for_if_mux_cse[102:96]==7'b0000000)
      & (fsm_output[2])) | (PECore_RunBias_if_for_13_operator_32_true_slc_operator_32_true_acc_13_svs
      & (fsm_output[4])));
  assign and_5953_nl = MUX_v_20_2_2(20'b00000000000000000000, mux1h_16_nl, nor_599_nl);
  assign nl_z_out_29 = PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_1_sva
      + conv_s2u_20_32(and_5953_nl);
  assign z_out_29 = nl_z_out_29[31:0];
  assign PECore_RunBias_if_for_if_and_9_nl = (~(adpfloat_tmp_is_zero_land_11_lpi_1_dfm_st
      | (input_mem_banks_read_read_data_lpi_1[87]))) & (fsm_output[1]);
  assign adpfloat_tmp_to_fixed_20U_14U_and_9_nl = adpfloat_tmp_is_zero_land_11_lpi_1_dfm_st
      & (~ (input_mem_banks_read_read_data_lpi_1[87])) & (fsm_output[1]);
  assign PECore_RunBias_if_for_if_and_10_nl = (input_mem_banks_read_read_data_lpi_1[87])
      & (fsm_output[1]);
  assign PECore_RunBias_if_for_if_mux1h_5_nl = MUX1HOT_v_20_4_2(z_out_43, z_out_49,
      act_port_reg_data_asn_2_itm, z_out_17, {(fsm_output[2]) , PECore_RunBias_if_for_if_and_9_nl
      , adpfloat_tmp_to_fixed_20U_14U_and_9_nl , PECore_RunBias_if_for_if_and_10_nl});
  assign PECore_RunBias_if_for_if_or_10_nl = MUX_v_20_2_2(PECore_RunBias_if_for_if_mux1h_5_nl,
      20'b11111111111111111111, or_dcpl_251);
  assign or_3882_nl = ((~ PECore_RunBias_if_for_12_operator_32_true_slc_operator_32_true_acc_13_svs)
      & (fsm_output[3])) | ((~ PECore_RunBias_if_for_14_operator_32_true_slc_operator_32_true_acc_13_svs)
      & (fsm_output[4]));
  assign mux_645_nl = MUX_v_20_2_2(PECore_RunBias_if_for_if_or_10_nl, z_out_45, or_3882_nl);
  assign nor_603_nl = ~((PECore_RunBias_if_for_12_operator_32_true_slc_operator_32_true_acc_13_svs
      & (fsm_output[3])) | (adpfloat_tmp_is_zero_land_11_lpi_1_dfm & (fsm_output[1]))
      | ((input_mem_banks_write_if_for_if_mux_cse[110:104]==7'b0000000) & (fsm_output[2]))
      | (PECore_RunBias_if_for_14_operator_32_true_slc_operator_32_true_acc_13_svs
      & (fsm_output[4])));
  assign and_5961_nl = MUX_v_20_2_2(20'b00000000000000000000, mux_645_nl, nor_603_nl);
  assign nl_z_out_30 = PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_11_sva
      + conv_s2u_20_32(and_5961_nl);
  assign z_out_30 = nl_z_out_30[31:0];
  assign PECore_RunBias_if_for_if_and_11_nl = (~(adpfloat_tmp_is_zero_land_6_lpi_1_dfm_st
      | (input_mem_banks_read_read_data_lpi_1[47]))) & (fsm_output[1]);
  assign adpfloat_tmp_to_fixed_20U_14U_and_10_nl = adpfloat_tmp_is_zero_land_6_lpi_1_dfm_st
      & (~ (input_mem_banks_read_read_data_lpi_1[47])) & (fsm_output[1]);
  assign PECore_RunBias_if_for_if_and_12_nl = (input_mem_banks_read_read_data_lpi_1[47])
      & (fsm_output[1]);
  assign PECore_RunBias_if_for_if_mux1h_6_nl = MUX1HOT_v_20_4_2(z_out_44, z_out_46,
      act_port_reg_data_asn_3_itm, z_out_20, {(fsm_output[2]) , PECore_RunBias_if_for_if_and_11_nl
      , adpfloat_tmp_to_fixed_20U_14U_and_10_nl , PECore_RunBias_if_for_if_and_12_nl});
  assign PECore_RunBias_if_for_if_or_11_nl = MUX_v_20_2_2(PECore_RunBias_if_for_if_mux1h_6_nl,
      20'b11111111111111111111, or_dcpl_251);
  assign or_3883_nl = ((~ PECore_RunBias_if_for_1_operator_32_true_slc_operator_32_true_acc_13_svs)
      & (fsm_output[3])) | ((~ PECore_RunBias_if_for_15_operator_32_true_slc_operator_32_true_acc_13_svs)
      & (fsm_output[4]));
  assign mux_646_nl = MUX_v_20_2_2(PECore_RunBias_if_for_if_or_11_nl, z_out_43, or_3883_nl);
  assign nor_607_nl = ~((PECore_RunBias_if_for_1_operator_32_true_slc_operator_32_true_acc_13_svs
      & (fsm_output[3])) | (adpfloat_tmp_is_zero_land_6_lpi_1_dfm & (fsm_output[1]))
      | ((input_mem_banks_write_if_for_if_mux_cse[118:112]==7'b0000000) & (fsm_output[2]))
      | (PECore_RunBias_if_for_15_operator_32_true_slc_operator_32_true_acc_13_svs
      & (fsm_output[4])));
  assign and_5968_nl = MUX_v_20_2_2(20'b00000000000000000000, mux_646_nl, nor_607_nl);
  assign nl_z_out_31 = PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_4_sva
      + conv_s2u_20_32(and_5968_nl);
  assign z_out_31 = nl_z_out_31[31:0];
  assign PECore_RunBias_if_for_if_and_13_nl = (~(adpfloat_tmp_is_zero_land_7_lpi_1_dfm_st
      | (input_mem_banks_read_read_data_lpi_1[55]))) & (fsm_output[1]);
  assign adpfloat_tmp_to_fixed_20U_14U_and_11_nl = adpfloat_tmp_is_zero_land_7_lpi_1_dfm_st
      & (~ (input_mem_banks_read_read_data_lpi_1[55])) & (fsm_output[1]);
  assign PECore_RunBias_if_for_if_and_14_nl = (input_mem_banks_read_read_data_lpi_1[55])
      & (fsm_output[1]);
  assign PECore_RunBias_if_for_if_mux1h_7_nl = MUX1HOT_v_20_4_2(z_out_45, z_out_47,
      act_port_reg_data_asn_itm, z_out_19, {(fsm_output[2]) , PECore_RunBias_if_for_if_and_13_nl
      , adpfloat_tmp_to_fixed_20U_14U_and_11_nl , PECore_RunBias_if_for_if_and_14_nl});
  assign PECore_RunBias_if_for_if_or_12_nl = MUX_v_20_2_2(PECore_RunBias_if_for_if_mux1h_7_nl,
      20'b11111111111111111111, or_dcpl_251);
  assign or_3884_nl = ((~ PECore_RunBias_if_for_2_operator_32_true_slc_operator_32_true_acc_13_svs)
      & (fsm_output[3])) | ((~ PECore_RunBias_if_for_16_operator_32_true_slc_operator_32_true_acc_13_svs)
      & (fsm_output[4]));
  assign mux_647_nl = MUX_v_20_2_2(PECore_RunBias_if_for_if_or_12_nl, z_out_44, or_3884_nl);
  assign nor_611_nl = ~((PECore_RunBias_if_for_2_operator_32_true_slc_operator_32_true_acc_13_svs
      & (fsm_output[3])) | (adpfloat_tmp_is_zero_land_7_lpi_1_dfm & (fsm_output[1]))
      | ((input_mem_banks_write_if_for_if_mux_cse[126:120]==7'b0000000) & (fsm_output[2]))
      | (PECore_RunBias_if_for_16_operator_32_true_slc_operator_32_true_acc_13_svs
      & (fsm_output[4])));
  assign and_5975_nl = MUX_v_20_2_2(20'b00000000000000000000, mux_647_nl, nor_611_nl);
  assign nl_z_out_32 = PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_5_sva
      + conv_s2u_20_32(and_5975_nl);
  assign z_out_32 = nl_z_out_32[31:0];
  assign PECore_RunBias_if_right_shift_mux_2_nl = MUX_v_3_2_2(pe_manager_adplfloat_bias_weight_0_sva,
      pe_manager_adplfloat_bias_weight_1_sva, pe_config_manager_counter_sva[0]);
  assign operator_3_false_mux_2_nl = MUX_v_3_2_2((~ PECore_RunBias_if_right_shift_mux_2_nl),
      (input_mem_banks_write_if_for_if_mux_cse[102:100]), fsm_output[2]);
  assign PECore_RunBias_if_right_shift_mux_3_nl = MUX_v_3_2_2(pe_manager_adplfloat_bias_input_0_sva,
      pe_manager_adplfloat_bias_input_1_sva, pe_config_manager_counter_sva[0]);
  assign operator_3_false_mux_3_nl = MUX_v_3_2_2((~ PECore_RunBias_if_right_shift_mux_3_nl),
      PECore_RunBias_if_for_if_bias_tmp2_mux_17, fsm_output[2]);
  assign nl_z_out_50 = conv_u2u_3_4(operator_3_false_mux_2_nl) + conv_u2u_3_4(operator_3_false_mux_3_nl);
  assign z_out_50 = nl_z_out_50[3:0];
  assign while_mux_440_cse = MUX_s_1_2_2(while_and_32_cse_1, while_and_30_itm_1,
      fsm_output[4]);
  assign and_5982_nl = PECore_UpdateFSM_switch_lp_nor_6_cse & (fsm_output[1]);
  assign PEManager_16U_GetInputAddr_1_PEManager_16U_GetInputAddr_1_mux_5_tmp = MUX_s_1_2_2((pe_config_manager_counter_sva[0]),
      (input_port_PopNB_mioi_idat_mxwt[128]), and_5982_nl);
  assign PEManager_16U_GetInputAddr_1_PEManager_16U_GetInputAddr_1_nor_nl = ~(or_tmp_3038
      | PEManager_16U_GetInputAddr_1_PEManager_16U_GetInputAddr_1_mux_5_tmp);
  assign PEManager_16U_GetInputAddr_1_and_1_nl = or_tmp_3038 & (~ PEManager_16U_GetInputAddr_1_PEManager_16U_GetInputAddr_1_mux_5_tmp);
  assign PEManager_16U_GetInputAddr_1_and_2_nl = (~ or_tmp_3038) & PEManager_16U_GetInputAddr_1_PEManager_16U_GetInputAddr_1_mux_5_tmp;
  assign PEManager_16U_GetInputAddr_1_and_3_nl = or_tmp_3038 & PEManager_16U_GetInputAddr_1_PEManager_16U_GetInputAddr_1_mux_5_tmp;
  assign z_out_41 = MUX1HOT_v_8_4_2((pe_manager_base_input_0_sva[7:0]), (pe_manager_base_bias_0_sva[7:0]),
      (pe_manager_base_input_1_sva[7:0]), (pe_manager_base_bias_1_sva[7:0]), {PEManager_16U_GetInputAddr_1_PEManager_16U_GetInputAddr_1_nor_nl
      , PEManager_16U_GetInputAddr_1_and_1_nl , PEManager_16U_GetInputAddr_1_and_2_nl
      , PEManager_16U_GetInputAddr_1_and_3_nl});
  assign adpfloat_tmp_to_fixed_20U_14U_mux1h_29_tmp = MUX1HOT_s_1_3_2((input_mem_banks_write_if_for_if_mux_cse[111]),
      (input_mem_banks_read_read_data_lpi_1[63]), (input_mem_banks_read_read_data_lpi_1[31]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])});
  assign adpfloat_tmp_to_fixed_20U_14U_adpfloat_tmp_to_fixed_20U_14U_nor_8_nl = ~((fsm_output[3])
      | adpfloat_tmp_to_fixed_20U_14U_mux1h_29_tmp);
  assign adpfloat_tmp_to_fixed_20U_14U_and_16_nl = (fsm_output[3]) & (~ adpfloat_tmp_to_fixed_20U_14U_mux1h_29_tmp);
  assign adpfloat_tmp_to_fixed_20U_14U_and_17_nl = (~ (fsm_output[4])) & adpfloat_tmp_to_fixed_20U_14U_mux1h_29_tmp;
  assign adpfloat_tmp_to_fixed_20U_14U_and_18_nl = (fsm_output[4]) & adpfloat_tmp_to_fixed_20U_14U_mux1h_29_tmp;
  assign z_out_43 = MUX1HOT_v_20_4_2(z_out_49, z_out_47, z_out_18, z_out_20, {adpfloat_tmp_to_fixed_20U_14U_adpfloat_tmp_to_fixed_20U_14U_nor_8_nl
      , adpfloat_tmp_to_fixed_20U_14U_and_16_nl , adpfloat_tmp_to_fixed_20U_14U_and_17_nl
      , adpfloat_tmp_to_fixed_20U_14U_and_18_nl});
  assign adpfloat_tmp_to_fixed_20U_14U_mux1h_30_tmp = MUX1HOT_s_1_3_2((input_mem_banks_write_if_for_if_mux_cse[119]),
      (input_mem_banks_read_read_data_lpi_1[71]), (input_mem_banks_read_read_data_lpi_1[39]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])});
  assign adpfloat_tmp_to_fixed_20U_14U_adpfloat_tmp_to_fixed_20U_14U_nor_nl = ~((fsm_output[4])
      | adpfloat_tmp_to_fixed_20U_14U_mux1h_30_tmp);
  assign adpfloat_tmp_to_fixed_20U_14U_and_20_nl = (fsm_output[4]) & (~ adpfloat_tmp_to_fixed_20U_14U_mux1h_30_tmp);
  assign adpfloat_tmp_to_fixed_20U_14U_and_21_nl = (~ (fsm_output[4])) & adpfloat_tmp_to_fixed_20U_14U_mux1h_30_tmp;
  assign adpfloat_tmp_to_fixed_20U_14U_and_22_nl = (fsm_output[4]) & adpfloat_tmp_to_fixed_20U_14U_mux1h_30_tmp;
  assign z_out_44 = MUX1HOT_v_20_4_2(z_out_48, z_out_46, z_out_19, z_out_17, {adpfloat_tmp_to_fixed_20U_14U_adpfloat_tmp_to_fixed_20U_14U_nor_nl
      , adpfloat_tmp_to_fixed_20U_14U_and_20_nl , adpfloat_tmp_to_fixed_20U_14U_and_21_nl
      , adpfloat_tmp_to_fixed_20U_14U_and_22_nl});
  assign adpfloat_tmp_to_fixed_20U_14U_mux1h_32_tmp = MUX1HOT_s_1_3_2((input_mem_banks_write_if_for_if_mux_cse[127]),
      (input_mem_banks_read_read_data_lpi_1[95]), (input_mem_banks_read_read_data_lpi_1[23]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])});
  assign adpfloat_tmp_to_fixed_20U_14U_and_23_nl = (fsm_output[2]) & (~ adpfloat_tmp_to_fixed_20U_14U_mux1h_32_tmp);
  assign adpfloat_tmp_to_fixed_20U_14U_and_24_nl = (fsm_output[3]) & (~ adpfloat_tmp_to_fixed_20U_14U_mux1h_32_tmp);
  assign adpfloat_tmp_to_fixed_20U_14U_and_25_nl = (fsm_output[4]) & (~ adpfloat_tmp_to_fixed_20U_14U_mux1h_32_tmp);
  assign adpfloat_tmp_to_fixed_20U_14U_and_26_nl = (~ (fsm_output[4])) & adpfloat_tmp_to_fixed_20U_14U_mux1h_32_tmp;
  assign adpfloat_tmp_to_fixed_20U_14U_and_27_nl = (fsm_output[4]) & adpfloat_tmp_to_fixed_20U_14U_mux1h_32_tmp;
  assign z_out_45 = MUX1HOT_v_20_5_2(z_out_47, z_out_49, z_out_48, z_out_20, z_out_19,
      {adpfloat_tmp_to_fixed_20U_14U_and_23_nl , adpfloat_tmp_to_fixed_20U_14U_and_24_nl
      , adpfloat_tmp_to_fixed_20U_14U_and_25_nl , adpfloat_tmp_to_fixed_20U_14U_and_26_nl
      , adpfloat_tmp_to_fixed_20U_14U_and_27_nl});

  function automatic  MUX1HOT_s_1_15_2;
    input  input_14;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [14:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    MUX1HOT_s_1_15_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_1_2;
    input  input_0;
    input  sel;
    reg  result;
  begin
    result = input_0 & sel;
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_5_2;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [4:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_8_2;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [7:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    MUX1HOT_s_1_8_2 = result;
  end
  endfunction


  function automatic [12:0] MUX1HOT_v_13_3_2;
    input [12:0] input_2;
    input [12:0] input_1;
    input [12:0] input_0;
    input [2:0] sel;
    reg [12:0] result;
  begin
    result = input_0 & {13{sel[0]}};
    result = result | (input_1 & {13{sel[1]}});
    result = result | (input_2 & {13{sel[2]}});
    MUX1HOT_v_13_3_2 = result;
  end
  endfunction


  function automatic [12:0] MUX1HOT_v_13_4_2;
    input [12:0] input_3;
    input [12:0] input_2;
    input [12:0] input_1;
    input [12:0] input_0;
    input [3:0] sel;
    reg [12:0] result;
  begin
    result = input_0 & {13{sel[0]}};
    result = result | (input_1 & {13{sel[1]}});
    result = result | (input_2 & {13{sel[2]}});
    result = result | (input_3 & {13{sel[3]}});
    MUX1HOT_v_13_4_2 = result;
  end
  endfunction


  function automatic [19:0] MUX1HOT_v_20_3_2;
    input [19:0] input_2;
    input [19:0] input_1;
    input [19:0] input_0;
    input [2:0] sel;
    reg [19:0] result;
  begin
    result = input_0 & {20{sel[0]}};
    result = result | (input_1 & {20{sel[1]}});
    result = result | (input_2 & {20{sel[2]}});
    MUX1HOT_v_20_3_2 = result;
  end
  endfunction


  function automatic [19:0] MUX1HOT_v_20_4_2;
    input [19:0] input_3;
    input [19:0] input_2;
    input [19:0] input_1;
    input [19:0] input_0;
    input [3:0] sel;
    reg [19:0] result;
  begin
    result = input_0 & {20{sel[0]}};
    result = result | (input_1 & {20{sel[1]}});
    result = result | (input_2 & {20{sel[2]}});
    result = result | (input_3 & {20{sel[3]}});
    MUX1HOT_v_20_4_2 = result;
  end
  endfunction


  function automatic [19:0] MUX1HOT_v_20_5_2;
    input [19:0] input_4;
    input [19:0] input_3;
    input [19:0] input_2;
    input [19:0] input_1;
    input [19:0] input_0;
    input [4:0] sel;
    reg [19:0] result;
  begin
    result = input_0 & {20{sel[0]}};
    result = result | (input_1 & {20{sel[1]}});
    result = result | (input_2 & {20{sel[2]}});
    result = result | (input_3 & {20{sel[3]}});
    result = result | (input_4 & {20{sel[4]}});
    MUX1HOT_v_20_5_2 = result;
  end
  endfunction


  function automatic [19:0] MUX1HOT_v_20_7_2;
    input [19:0] input_6;
    input [19:0] input_5;
    input [19:0] input_4;
    input [19:0] input_3;
    input [19:0] input_2;
    input [19:0] input_1;
    input [19:0] input_0;
    input [6:0] sel;
    reg [19:0] result;
  begin
    result = input_0 & {20{sel[0]}};
    result = result | (input_1 & {20{sel[1]}});
    result = result | (input_2 & {20{sel[2]}});
    result = result | (input_3 & {20{sel[3]}});
    result = result | (input_4 & {20{sel[4]}});
    result = result | (input_5 & {20{sel[5]}});
    result = result | (input_6 & {20{sel[6]}});
    MUX1HOT_v_20_7_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_3_2;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [2:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | (input_1 & {32{sel[1]}});
    result = result | (input_2 & {32{sel[2]}});
    MUX1HOT_v_32_3_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_4_2;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [3:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | (input_1 & {32{sel[1]}});
    result = result | (input_2 & {32{sel[2]}});
    result = result | (input_3 & {32{sel[3]}});
    MUX1HOT_v_32_4_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_5_2;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [4:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    MUX1HOT_v_4_5_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_7_2;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [6:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    MUX1HOT_v_4_7_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_3_2;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [2:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    MUX1HOT_v_5_3_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_4_2;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [3:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    MUX1HOT_v_5_4_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_5_2;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [4:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    MUX1HOT_v_5_5_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_3_2;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [2:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_4_2;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [3:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    MUX1HOT_v_7_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_4_2;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [3:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    MUX1HOT_v_8_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_5_2;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [4:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    MUX1HOT_v_8_5_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_6_2;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [5:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    MUX1HOT_v_8_6_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_16_2;
    input  input_0;
    input  input_1;
    input  input_2;
    input  input_3;
    input  input_4;
    input  input_5;
    input  input_6;
    input  input_7;
    input  input_8;
    input  input_9;
    input  input_10;
    input  input_11;
    input  input_12;
    input  input_13;
    input  input_14;
    input  input_15;
    input [3:0] sel;
    reg  result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_s_1_16_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_32_2;
    input  input_0;
    input  input_1;
    input  input_2;
    input  input_3;
    input  input_4;
    input  input_5;
    input  input_6;
    input  input_7;
    input  input_8;
    input  input_9;
    input  input_10;
    input  input_11;
    input  input_12;
    input  input_13;
    input  input_14;
    input  input_15;
    input  input_16;
    input  input_17;
    input  input_18;
    input  input_19;
    input  input_20;
    input  input_21;
    input  input_22;
    input  input_23;
    input  input_24;
    input  input_25;
    input  input_26;
    input  input_27;
    input  input_28;
    input  input_29;
    input  input_30;
    input  input_31;
    input [4:0] sel;
    reg  result;
  begin
    case (sel)
      5'b00000 : begin
        result = input_0;
      end
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      5'b10111 : begin
        result = input_23;
      end
      5'b11000 : begin
        result = input_24;
      end
      5'b11001 : begin
        result = input_25;
      end
      5'b11010 : begin
        result = input_26;
      end
      5'b11011 : begin
        result = input_27;
      end
      5'b11100 : begin
        result = input_28;
      end
      5'b11101 : begin
        result = input_29;
      end
      5'b11110 : begin
        result = input_30;
      end
      default : begin
        result = input_31;
      end
    endcase
    MUX_s_1_32_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input  sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_16_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input [11:0] input_2;
    input [11:0] input_3;
    input [11:0] input_4;
    input [11:0] input_5;
    input [11:0] input_6;
    input [11:0] input_7;
    input [11:0] input_8;
    input [11:0] input_9;
    input [11:0] input_10;
    input [11:0] input_11;
    input [11:0] input_12;
    input [11:0] input_13;
    input [11:0] input_14;
    input [11:0] input_15;
    input [3:0] sel;
    reg [11:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_12_16_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input  sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input  sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [14:0] MUX_v_15_2_2;
    input [14:0] input_0;
    input [14:0] input_1;
    input  sel;
    reg [14:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_15_2_2 = result;
  end
  endfunction


  function automatic [168:0] MUX_v_169_2_2;
    input [168:0] input_0;
    input [168:0] input_1;
    input  sel;
    reg [168:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_169_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input  sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_32_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [1:0] input_2;
    input [1:0] input_3;
    input [1:0] input_4;
    input [1:0] input_5;
    input [1:0] input_6;
    input [1:0] input_7;
    input [1:0] input_8;
    input [1:0] input_9;
    input [1:0] input_10;
    input [1:0] input_11;
    input [1:0] input_12;
    input [1:0] input_13;
    input [1:0] input_14;
    input [1:0] input_15;
    input [1:0] input_16;
    input [1:0] input_17;
    input [1:0] input_18;
    input [1:0] input_19;
    input [1:0] input_20;
    input [1:0] input_21;
    input [1:0] input_22;
    input [1:0] input_23;
    input [1:0] input_24;
    input [1:0] input_25;
    input [1:0] input_26;
    input [1:0] input_27;
    input [1:0] input_28;
    input [1:0] input_29;
    input [1:0] input_30;
    input [1:0] input_31;
    input [4:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      5'b00000 : begin
        result = input_0;
      end
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      5'b10111 : begin
        result = input_23;
      end
      5'b11000 : begin
        result = input_24;
      end
      5'b11001 : begin
        result = input_25;
      end
      5'b11010 : begin
        result = input_26;
      end
      5'b11011 : begin
        result = input_27;
      end
      5'b11100 : begin
        result = input_28;
      end
      5'b11101 : begin
        result = input_29;
      end
      5'b11110 : begin
        result = input_30;
      end
      default : begin
        result = input_31;
      end
    endcase
    MUX_v_2_32_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_4_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [31:0] input_3;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_32_4_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_32_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [2:0] input_2;
    input [2:0] input_3;
    input [2:0] input_4;
    input [2:0] input_5;
    input [2:0] input_6;
    input [2:0] input_7;
    input [2:0] input_8;
    input [2:0] input_9;
    input [2:0] input_10;
    input [2:0] input_11;
    input [2:0] input_12;
    input [2:0] input_13;
    input [2:0] input_14;
    input [2:0] input_15;
    input [2:0] input_16;
    input [2:0] input_17;
    input [2:0] input_18;
    input [2:0] input_19;
    input [2:0] input_20;
    input [2:0] input_21;
    input [2:0] input_22;
    input [2:0] input_23;
    input [2:0] input_24;
    input [2:0] input_25;
    input [2:0] input_26;
    input [2:0] input_27;
    input [2:0] input_28;
    input [2:0] input_29;
    input [2:0] input_30;
    input [2:0] input_31;
    input [4:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      5'b00000 : begin
        result = input_0;
      end
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      5'b10111 : begin
        result = input_23;
      end
      5'b11000 : begin
        result = input_24;
      end
      5'b11001 : begin
        result = input_25;
      end
      5'b11010 : begin
        result = input_26;
      end
      5'b11011 : begin
        result = input_27;
      end
      5'b11100 : begin
        result = input_28;
      end
      5'b11101 : begin
        result = input_29;
      end
      5'b11110 : begin
        result = input_30;
      end
      default : begin
        result = input_31;
      end
    endcase
    MUX_v_3_32_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_32_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [3:0] input_8;
    input [3:0] input_9;
    input [3:0] input_10;
    input [3:0] input_11;
    input [3:0] input_12;
    input [3:0] input_13;
    input [3:0] input_14;
    input [3:0] input_15;
    input [3:0] input_16;
    input [3:0] input_17;
    input [3:0] input_18;
    input [3:0] input_19;
    input [3:0] input_20;
    input [3:0] input_21;
    input [3:0] input_22;
    input [3:0] input_23;
    input [3:0] input_24;
    input [3:0] input_25;
    input [3:0] input_26;
    input [3:0] input_27;
    input [3:0] input_28;
    input [3:0] input_29;
    input [3:0] input_30;
    input [3:0] input_31;
    input [4:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      5'b00000 : begin
        result = input_0;
      end
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      5'b10111 : begin
        result = input_23;
      end
      5'b11000 : begin
        result = input_24;
      end
      5'b11001 : begin
        result = input_25;
      end
      5'b11010 : begin
        result = input_26;
      end
      5'b11011 : begin
        result = input_27;
      end
      5'b11100 : begin
        result = input_28;
      end
      5'b11101 : begin
        result = input_29;
      end
      5'b11110 : begin
        result = input_30;
      end
      default : begin
        result = input_31;
      end
    endcase
    MUX_v_4_32_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input  sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_32_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [4:0] input_2;
    input [4:0] input_3;
    input [4:0] input_4;
    input [4:0] input_5;
    input [4:0] input_6;
    input [4:0] input_7;
    input [4:0] input_8;
    input [4:0] input_9;
    input [4:0] input_10;
    input [4:0] input_11;
    input [4:0] input_12;
    input [4:0] input_13;
    input [4:0] input_14;
    input [4:0] input_15;
    input [4:0] input_16;
    input [4:0] input_17;
    input [4:0] input_18;
    input [4:0] input_19;
    input [4:0] input_20;
    input [4:0] input_21;
    input [4:0] input_22;
    input [4:0] input_23;
    input [4:0] input_24;
    input [4:0] input_25;
    input [4:0] input_26;
    input [4:0] input_27;
    input [4:0] input_28;
    input [4:0] input_29;
    input [4:0] input_30;
    input [4:0] input_31;
    input [4:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      5'b00000 : begin
        result = input_0;
      end
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      5'b10111 : begin
        result = input_23;
      end
      5'b11000 : begin
        result = input_24;
      end
      5'b11001 : begin
        result = input_25;
      end
      5'b11010 : begin
        result = input_26;
      end
      5'b11011 : begin
        result = input_27;
      end
      5'b11100 : begin
        result = input_28;
      end
      5'b11101 : begin
        result = input_29;
      end
      5'b11110 : begin
        result = input_30;
      end
      default : begin
        result = input_31;
      end
    endcase
    MUX_v_5_32_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_32_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [5:0] input_2;
    input [5:0] input_3;
    input [5:0] input_4;
    input [5:0] input_5;
    input [5:0] input_6;
    input [5:0] input_7;
    input [5:0] input_8;
    input [5:0] input_9;
    input [5:0] input_10;
    input [5:0] input_11;
    input [5:0] input_12;
    input [5:0] input_13;
    input [5:0] input_14;
    input [5:0] input_15;
    input [5:0] input_16;
    input [5:0] input_17;
    input [5:0] input_18;
    input [5:0] input_19;
    input [5:0] input_20;
    input [5:0] input_21;
    input [5:0] input_22;
    input [5:0] input_23;
    input [5:0] input_24;
    input [5:0] input_25;
    input [5:0] input_26;
    input [5:0] input_27;
    input [5:0] input_28;
    input [5:0] input_29;
    input [5:0] input_30;
    input [5:0] input_31;
    input [4:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      5'b00000 : begin
        result = input_0;
      end
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      5'b10111 : begin
        result = input_23;
      end
      5'b11000 : begin
        result = input_24;
      end
      5'b11001 : begin
        result = input_25;
      end
      5'b11010 : begin
        result = input_26;
      end
      5'b11011 : begin
        result = input_27;
      end
      5'b11100 : begin
        result = input_28;
      end
      5'b11101 : begin
        result = input_29;
      end
      5'b11110 : begin
        result = input_30;
      end
      default : begin
        result = input_31;
      end
    endcase
    MUX_v_6_32_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_32_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [6:0] input_2;
    input [6:0] input_3;
    input [6:0] input_4;
    input [6:0] input_5;
    input [6:0] input_6;
    input [6:0] input_7;
    input [6:0] input_8;
    input [6:0] input_9;
    input [6:0] input_10;
    input [6:0] input_11;
    input [6:0] input_12;
    input [6:0] input_13;
    input [6:0] input_14;
    input [6:0] input_15;
    input [6:0] input_16;
    input [6:0] input_17;
    input [6:0] input_18;
    input [6:0] input_19;
    input [6:0] input_20;
    input [6:0] input_21;
    input [6:0] input_22;
    input [6:0] input_23;
    input [6:0] input_24;
    input [6:0] input_25;
    input [6:0] input_26;
    input [6:0] input_27;
    input [6:0] input_28;
    input [6:0] input_29;
    input [6:0] input_30;
    input [6:0] input_31;
    input [4:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      5'b00000 : begin
        result = input_0;
      end
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      5'b10111 : begin
        result = input_23;
      end
      5'b11000 : begin
        result = input_24;
      end
      5'b11001 : begin
        result = input_25;
      end
      5'b11010 : begin
        result = input_26;
      end
      5'b11011 : begin
        result = input_27;
      end
      5'b11100 : begin
        result = input_28;
      end
      5'b11101 : begin
        result = input_29;
      end
      5'b11110 : begin
        result = input_30;
      end
      default : begin
        result = input_31;
      end
    endcase
    MUX_v_7_32_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_16_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [7:0] input_8;
    input [7:0] input_9;
    input [7:0] input_10;
    input [7:0] input_11;
    input [7:0] input_12;
    input [7:0] input_13;
    input [7:0] input_14;
    input [7:0] input_15;
    input [3:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_8_16_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_32_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [7:0] input_8;
    input [7:0] input_9;
    input [7:0] input_10;
    input [7:0] input_11;
    input [7:0] input_12;
    input [7:0] input_13;
    input [7:0] input_14;
    input [7:0] input_15;
    input [7:0] input_16;
    input [7:0] input_17;
    input [7:0] input_18;
    input [7:0] input_19;
    input [7:0] input_20;
    input [7:0] input_21;
    input [7:0] input_22;
    input [7:0] input_23;
    input [7:0] input_24;
    input [7:0] input_25;
    input [7:0] input_26;
    input [7:0] input_27;
    input [7:0] input_28;
    input [7:0] input_29;
    input [7:0] input_30;
    input [7:0] input_31;
    input [4:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      5'b00000 : begin
        result = input_0;
      end
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      5'b10111 : begin
        result = input_23;
      end
      5'b11000 : begin
        result = input_24;
      end
      5'b11001 : begin
        result = input_25;
      end
      5'b11010 : begin
        result = input_26;
      end
      5'b11011 : begin
        result = input_27;
      end
      5'b11100 : begin
        result = input_28;
      end
      5'b11101 : begin
        result = input_29;
      end
      5'b11110 : begin
        result = input_30;
      end
      default : begin
        result = input_31;
      end
    endcase
    MUX_v_8_32_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_14_1_13;
    input [13:0] vector;
    reg [13:0] tmp;
  begin
    tmp = vector >> 13;
    readslicef_14_1_13 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function automatic [12:0] signext_13_1;
    input  vector;
  begin
    signext_13_1= {{12{vector}}, vector};
  end
  endfunction


  function automatic [13:0] signext_14_1;
    input  vector;
  begin
    signext_14_1= {{13{vector}}, vector};
  end
  endfunction


  function automatic [14:0] signext_15_1;
    input  vector;
  begin
    signext_15_1= {{14{vector}}, vector};
  end
  endfunction


  function automatic [15:0] signext_16_1;
    input  vector;
  begin
    signext_16_1= {{15{vector}}, vector};
  end
  endfunction


  function automatic [2:0] signext_3_2;
    input [1:0] vector;
  begin
    signext_3_2= {{1{vector[1]}}, vector};
  end
  endfunction


  function automatic [3:0] signext_4_1;
    input  vector;
  begin
    signext_4_1= {{3{vector}}, vector};
  end
  endfunction


  function automatic [7:0] signext_8_1;
    input  vector;
  begin
    signext_8_1= {{7{vector}}, vector};
  end
  endfunction


  function automatic [4:0] conv_s2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_s2s_4_5 = {vector[3], vector};
  end
  endfunction


  function automatic [4:0] conv_s2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_s2u_4_5 = {vector[3], vector};
  end
  endfunction


  function automatic [13:0] conv_s2u_13_14 ;
    input [12:0]  vector ;
  begin
    conv_s2u_13_14 = {vector[12], vector};
  end
  endfunction


  function automatic [31:0] conv_s2u_20_32 ;
    input [19:0]  vector ;
  begin
    conv_s2u_20_32 = {{12{vector[19]}}, vector};
  end
  endfunction


  function automatic [32:0] conv_s2u_32_33 ;
    input [31:0]  vector ;
  begin
    conv_s2u_32_33 = {vector[31], vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_3_5 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_5 = {{2{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore
// ------------------------------------------------------------------


module PECore (
  clk, rst, start_val, start_rdy, start_msg, input_port_val, input_port_rdy, input_port_msg,
      rva_in_val, rva_in_rdy, rva_in_msg, rva_out_val, rva_out_rdy, rva_out_msg,
      act_port_val, act_port_rdy, act_port_msg, SC_SRAM_CONFIG
);
  input clk;
  input rst;
  input start_val;
  output start_rdy;
  input start_msg;
  input input_port_val;
  output input_port_rdy;
  input [137:0] input_port_msg;
  input rva_in_val;
  output rva_in_rdy;
  input [168:0] rva_in_msg;
  output rva_out_val;
  input rva_out_rdy;
  output [127:0] rva_out_msg;
  output act_port_val;
  input act_port_rdy;
  output [319:0] act_port_msg;
  input [31:0] SC_SRAM_CONFIG;


  // Interconnect Declarations
  wire weight_mem_banks_bank_array_impl_data0_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data0_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data0_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data0_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data1_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data1_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data1_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data1_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data1_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data2_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data2_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data2_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data2_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data2_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data3_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data3_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data3_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data3_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data3_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data4_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data4_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data4_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data4_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data4_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data5_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data5_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data5_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data5_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data5_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data6_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data6_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data6_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data6_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data6_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data7_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data7_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data7_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data7_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data7_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data8_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data8_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data8_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data8_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data8_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data9_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data9_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data9_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data9_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data9_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data10_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data10_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data10_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data10_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data10_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data11_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data11_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data11_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data11_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data11_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data12_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data12_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data12_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data12_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data12_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data13_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data13_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data13_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data13_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data13_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data14_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data14_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data14_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data14_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data14_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data15_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data15_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data15_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data15_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data15_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire input_mem_banks_bank_array_impl_data0_rsci_clken_d;
  wire [127:0] input_mem_banks_bank_array_impl_data0_rsci_d_d;
  wire [127:0] input_mem_banks_bank_array_impl_data0_rsci_q_d;
  wire [7:0] input_mem_banks_bank_array_impl_data0_rsci_radr_d;
  wire [7:0] input_mem_banks_bank_array_impl_data0_rsci_wadr_d;
  wire input_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data0_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data0_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data0_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data0_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data0_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data0_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data1_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data1_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data1_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data1_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data1_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data1_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data2_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data2_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data2_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data2_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data2_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data2_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data3_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data3_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data3_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data3_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data3_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data3_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data4_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data4_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data4_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data4_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data4_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data4_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data5_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data5_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data5_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data5_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data5_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data5_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data6_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data6_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data6_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data6_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data6_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data6_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data7_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data7_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data7_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data7_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data7_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data7_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data8_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data8_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data8_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data8_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data8_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data8_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data9_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data9_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data9_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data9_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data9_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data9_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data10_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data10_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data10_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data10_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data10_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data10_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data11_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data11_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data11_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data11_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data11_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data11_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data12_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data12_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data12_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data12_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data12_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data12_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data13_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data13_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data13_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data13_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data13_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data13_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data14_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data14_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data14_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data14_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data14_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data14_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data15_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data15_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data15_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data15_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data15_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data15_rsc_wadr;
  wire input_mem_banks_bank_array_impl_data0_rsc_clken;
  wire [127:0] input_mem_banks_bank_array_impl_data0_rsc_q;
  wire [7:0] input_mem_banks_bank_array_impl_data0_rsc_radr;
  wire input_mem_banks_bank_array_impl_data0_rsc_we;
  wire [127:0] input_mem_banks_bank_array_impl_data0_rsc_d;
  wire [7:0] input_mem_banks_bank_array_impl_data0_rsc_wadr;
  wire [11:0] weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_iff;
  wire weight_mem_banks_bank_array_impl_data0_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data1_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data2_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data3_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data4_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data5_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data6_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data7_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data8_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data9_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data10_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data11_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data12_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data13_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data14_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data15_rsci_we_d_iff;
  wire input_mem_banks_bank_array_impl_data0_rsci_we_d_iff;

  // Helper signals
  wire [2:0] state;
  assign state = {PECore_PECoreRun_inst.state_2_0_sva_2, PECore_PECoreRun_inst.state_2_0_sva_1, PECore_PECoreRun_inst.state_2_0_sva_0};

  wire is_start;
  assign is_start = PECore_PECoreRun_inst.is_start_sva;

  // PE_Config signals
  wire pe_config_is_valid = PECore_PECoreRun_inst.pe_config_is_valid_sva;
  wire pe_config_is_zero_first = PECore_PECoreRun_inst.pe_config_is_zero_first_sva;
  wire pe_config_is_cluster = PECore_PECoreRun_inst.pe_config_is_cluster_sva;
  wire pe_config_is_bias = PECore_PECoreRun_inst.pe_config_is_bias_sva;
  wire [3:0] pe_config_num_manager = PECore_PECoreRun_inst.pe_config_num_manager_sva;
  wire [7:0] pe_config_num_output = PECore_PECoreRun_inst.pe_config_num_output_sva;
  wire [3:0] pe_config_manager_counter = PECore_PECoreRun_inst.pe_config_manager_counter_sva;
  wire [7:0] pe_config_input_counter = PECore_PECoreRun_inst.pe_config_input_counter_sva;
  wire [7:0] pe_config_output_counter = PECore_PECoreRun_inst.pe_config_output_counter_sva;

  // RVA_IN Decode
  wire rva_in_rw = rva_in_msg[168];
  wire [15:0] rva_in_wstrb = rva_in_msg[167:152];
  wire [23:0] rva_in_addr = rva_in_msg[151:128];
  wire [127:0] rva_in_data = rva_in_msg[127:0];

  // Interconnect Declarations for Component Instantiations 
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1)) weight_mem_banks_bank_array_impl_data0_rsc_comp (
      .clk(clk),
      .clken(weight_mem_banks_bank_array_impl_data0_rsc_clken),
      .d(weight_mem_banks_bank_array_impl_data0_rsc_d),
      .q(weight_mem_banks_bank_array_impl_data0_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data0_rsc_radr),
      .wadr(weight_mem_banks_bank_array_impl_data0_rsc_wadr),
      .we(weight_mem_banks_bank_array_impl_data0_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1)) weight_mem_banks_bank_array_impl_data1_rsc_comp (
      .clk(clk),
      .clken(weight_mem_banks_bank_array_impl_data1_rsc_clken),
      .d(weight_mem_banks_bank_array_impl_data1_rsc_d),
      .q(weight_mem_banks_bank_array_impl_data1_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data1_rsc_radr),
      .wadr(weight_mem_banks_bank_array_impl_data1_rsc_wadr),
      .we(weight_mem_banks_bank_array_impl_data1_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1)) weight_mem_banks_bank_array_impl_data2_rsc_comp (
      .clk(clk),
      .clken(weight_mem_banks_bank_array_impl_data2_rsc_clken),
      .d(weight_mem_banks_bank_array_impl_data2_rsc_d),
      .q(weight_mem_banks_bank_array_impl_data2_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data2_rsc_radr),
      .wadr(weight_mem_banks_bank_array_impl_data2_rsc_wadr),
      .we(weight_mem_banks_bank_array_impl_data2_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1)) weight_mem_banks_bank_array_impl_data3_rsc_comp (
      .clk(clk),
      .clken(weight_mem_banks_bank_array_impl_data3_rsc_clken),
      .d(weight_mem_banks_bank_array_impl_data3_rsc_d),
      .q(weight_mem_banks_bank_array_impl_data3_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data3_rsc_radr),
      .wadr(weight_mem_banks_bank_array_impl_data3_rsc_wadr),
      .we(weight_mem_banks_bank_array_impl_data3_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1)) weight_mem_banks_bank_array_impl_data4_rsc_comp (
      .clk(clk),
      .clken(weight_mem_banks_bank_array_impl_data4_rsc_clken),
      .d(weight_mem_banks_bank_array_impl_data4_rsc_d),
      .q(weight_mem_banks_bank_array_impl_data4_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data4_rsc_radr),
      .wadr(weight_mem_banks_bank_array_impl_data4_rsc_wadr),
      .we(weight_mem_banks_bank_array_impl_data4_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1)) weight_mem_banks_bank_array_impl_data5_rsc_comp (
      .clk(clk),
      .clken(weight_mem_banks_bank_array_impl_data5_rsc_clken),
      .d(weight_mem_banks_bank_array_impl_data5_rsc_d),
      .q(weight_mem_banks_bank_array_impl_data5_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data5_rsc_radr),
      .wadr(weight_mem_banks_bank_array_impl_data5_rsc_wadr),
      .we(weight_mem_banks_bank_array_impl_data5_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1)) weight_mem_banks_bank_array_impl_data6_rsc_comp (
      .clk(clk),
      .clken(weight_mem_banks_bank_array_impl_data6_rsc_clken),
      .d(weight_mem_banks_bank_array_impl_data6_rsc_d),
      .q(weight_mem_banks_bank_array_impl_data6_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data6_rsc_radr),
      .wadr(weight_mem_banks_bank_array_impl_data6_rsc_wadr),
      .we(weight_mem_banks_bank_array_impl_data6_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1)) weight_mem_banks_bank_array_impl_data7_rsc_comp (
      .clk(clk),
      .clken(weight_mem_banks_bank_array_impl_data7_rsc_clken),
      .d(weight_mem_banks_bank_array_impl_data7_rsc_d),
      .q(weight_mem_banks_bank_array_impl_data7_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data7_rsc_radr),
      .wadr(weight_mem_banks_bank_array_impl_data7_rsc_wadr),
      .we(weight_mem_banks_bank_array_impl_data7_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1)) weight_mem_banks_bank_array_impl_data8_rsc_comp (
      .clk(clk),
      .clken(weight_mem_banks_bank_array_impl_data8_rsc_clken),
      .d(weight_mem_banks_bank_array_impl_data8_rsc_d),
      .q(weight_mem_banks_bank_array_impl_data8_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data8_rsc_radr),
      .wadr(weight_mem_banks_bank_array_impl_data8_rsc_wadr),
      .we(weight_mem_banks_bank_array_impl_data8_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1)) weight_mem_banks_bank_array_impl_data9_rsc_comp (
      .clk(clk),
      .clken(weight_mem_banks_bank_array_impl_data9_rsc_clken),
      .d(weight_mem_banks_bank_array_impl_data9_rsc_d),
      .q(weight_mem_banks_bank_array_impl_data9_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data9_rsc_radr),
      .wadr(weight_mem_banks_bank_array_impl_data9_rsc_wadr),
      .we(weight_mem_banks_bank_array_impl_data9_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1)) weight_mem_banks_bank_array_impl_data10_rsc_comp (
      .clk(clk),
      .clken(weight_mem_banks_bank_array_impl_data10_rsc_clken),
      .d(weight_mem_banks_bank_array_impl_data10_rsc_d),
      .q(weight_mem_banks_bank_array_impl_data10_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data10_rsc_radr),
      .wadr(weight_mem_banks_bank_array_impl_data10_rsc_wadr),
      .we(weight_mem_banks_bank_array_impl_data10_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1)) weight_mem_banks_bank_array_impl_data11_rsc_comp (
      .clk(clk),
      .clken(weight_mem_banks_bank_array_impl_data11_rsc_clken),
      .d(weight_mem_banks_bank_array_impl_data11_rsc_d),
      .q(weight_mem_banks_bank_array_impl_data11_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data11_rsc_radr),
      .wadr(weight_mem_banks_bank_array_impl_data11_rsc_wadr),
      .we(weight_mem_banks_bank_array_impl_data11_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1)) weight_mem_banks_bank_array_impl_data12_rsc_comp (
      .clk(clk),
      .clken(weight_mem_banks_bank_array_impl_data12_rsc_clken),
      .d(weight_mem_banks_bank_array_impl_data12_rsc_d),
      .q(weight_mem_banks_bank_array_impl_data12_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data12_rsc_radr),
      .wadr(weight_mem_banks_bank_array_impl_data12_rsc_wadr),
      .we(weight_mem_banks_bank_array_impl_data12_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1)) weight_mem_banks_bank_array_impl_data13_rsc_comp (
      .clk(clk),
      .clken(weight_mem_banks_bank_array_impl_data13_rsc_clken),
      .d(weight_mem_banks_bank_array_impl_data13_rsc_d),
      .q(weight_mem_banks_bank_array_impl_data13_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data13_rsc_radr),
      .wadr(weight_mem_banks_bank_array_impl_data13_rsc_wadr),
      .we(weight_mem_banks_bank_array_impl_data13_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1)) weight_mem_banks_bank_array_impl_data14_rsc_comp (
      .clk(clk),
      .clken(weight_mem_banks_bank_array_impl_data14_rsc_clken),
      .d(weight_mem_banks_bank_array_impl_data14_rsc_d),
      .q(weight_mem_banks_bank_array_impl_data14_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data14_rsc_radr),
      .wadr(weight_mem_banks_bank_array_impl_data14_rsc_wadr),
      .we(weight_mem_banks_bank_array_impl_data14_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1)) weight_mem_banks_bank_array_impl_data15_rsc_comp (
      .clk(clk),
      .clken(weight_mem_banks_bank_array_impl_data15_rsc_clken),
      .d(weight_mem_banks_bank_array_impl_data15_rsc_d),
      .q(weight_mem_banks_bank_array_impl_data15_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data15_rsc_radr),
      .wadr(weight_mem_banks_bank_array_impl_data15_rsc_wadr),
      .we(weight_mem_banks_bank_array_impl_data15_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd8),
  .data_width(32'sd128),
  .depth(32'sd256),
  .latency(32'sd1)) input_mem_banks_bank_array_impl_data0_rsc_comp (
      .clk(clk),
      .clken(input_mem_banks_bank_array_impl_data0_rsc_clken),
      .d(input_mem_banks_bank_array_impl_data0_rsc_d),
      .q(input_mem_banks_bank_array_impl_data0_rsc_q),
      .radr(input_mem_banks_bank_array_impl_data0_rsc_radr),
      .wadr(input_mem_banks_bank_array_impl_data0_rsc_wadr),
      .we(input_mem_banks_bank_array_impl_data0_rsc_we)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_108_12_128_4096_4096_128_1_gen
      weight_mem_banks_bank_array_impl_data0_rsci (
      .clken(weight_mem_banks_bank_array_impl_data0_rsc_clken),
      .q(weight_mem_banks_bank_array_impl_data0_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data0_rsc_radr),
      .we(weight_mem_banks_bank_array_impl_data0_rsc_we),
      .d(weight_mem_banks_bank_array_impl_data0_rsc_d),
      .wadr(weight_mem_banks_bank_array_impl_data0_rsc_wadr),
      .clken_d(weight_mem_banks_bank_array_impl_data0_rsci_clken_d),
      .d_d(weight_mem_banks_bank_array_impl_data0_rsci_d_d),
      .q_d(weight_mem_banks_bank_array_impl_data0_rsci_q_d),
      .radr_d(weight_mem_banks_bank_array_impl_data0_rsci_radr_d),
      .wadr_d(weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_array_impl_data0_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_array_impl_data0_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_109_12_128_4096_4096_128_1_gen
      weight_mem_banks_bank_array_impl_data1_rsci (
      .clken(weight_mem_banks_bank_array_impl_data1_rsc_clken),
      .q(weight_mem_banks_bank_array_impl_data1_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data1_rsc_radr),
      .we(weight_mem_banks_bank_array_impl_data1_rsc_we),
      .d(weight_mem_banks_bank_array_impl_data1_rsc_d),
      .wadr(weight_mem_banks_bank_array_impl_data1_rsc_wadr),
      .clken_d(weight_mem_banks_bank_array_impl_data1_rsci_clken_d),
      .d_d(weight_mem_banks_bank_array_impl_data1_rsci_d_d),
      .q_d(weight_mem_banks_bank_array_impl_data1_rsci_q_d),
      .radr_d(weight_mem_banks_bank_array_impl_data1_rsci_radr_d),
      .wadr_d(weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_array_impl_data1_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_array_impl_data1_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data1_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_110_12_128_4096_4096_128_1_gen
      weight_mem_banks_bank_array_impl_data2_rsci (
      .clken(weight_mem_banks_bank_array_impl_data2_rsc_clken),
      .q(weight_mem_banks_bank_array_impl_data2_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data2_rsc_radr),
      .we(weight_mem_banks_bank_array_impl_data2_rsc_we),
      .d(weight_mem_banks_bank_array_impl_data2_rsc_d),
      .wadr(weight_mem_banks_bank_array_impl_data2_rsc_wadr),
      .clken_d(weight_mem_banks_bank_array_impl_data2_rsci_clken_d),
      .d_d(weight_mem_banks_bank_array_impl_data2_rsci_d_d),
      .q_d(weight_mem_banks_bank_array_impl_data2_rsci_q_d),
      .radr_d(weight_mem_banks_bank_array_impl_data2_rsci_radr_d),
      .wadr_d(weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_array_impl_data2_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_array_impl_data2_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data2_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_111_12_128_4096_4096_128_1_gen
      weight_mem_banks_bank_array_impl_data3_rsci (
      .clken(weight_mem_banks_bank_array_impl_data3_rsc_clken),
      .q(weight_mem_banks_bank_array_impl_data3_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data3_rsc_radr),
      .we(weight_mem_banks_bank_array_impl_data3_rsc_we),
      .d(weight_mem_banks_bank_array_impl_data3_rsc_d),
      .wadr(weight_mem_banks_bank_array_impl_data3_rsc_wadr),
      .clken_d(weight_mem_banks_bank_array_impl_data3_rsci_clken_d),
      .d_d(weight_mem_banks_bank_array_impl_data3_rsci_d_d),
      .q_d(weight_mem_banks_bank_array_impl_data3_rsci_q_d),
      .radr_d(weight_mem_banks_bank_array_impl_data3_rsci_radr_d),
      .wadr_d(weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_array_impl_data3_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_array_impl_data3_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data3_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_112_12_128_4096_4096_128_1_gen
      weight_mem_banks_bank_array_impl_data4_rsci (
      .clken(weight_mem_banks_bank_array_impl_data4_rsc_clken),
      .q(weight_mem_banks_bank_array_impl_data4_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data4_rsc_radr),
      .we(weight_mem_banks_bank_array_impl_data4_rsc_we),
      .d(weight_mem_banks_bank_array_impl_data4_rsc_d),
      .wadr(weight_mem_banks_bank_array_impl_data4_rsc_wadr),
      .clken_d(weight_mem_banks_bank_array_impl_data4_rsci_clken_d),
      .d_d(weight_mem_banks_bank_array_impl_data4_rsci_d_d),
      .q_d(weight_mem_banks_bank_array_impl_data4_rsci_q_d),
      .radr_d(weight_mem_banks_bank_array_impl_data4_rsci_radr_d),
      .wadr_d(weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_array_impl_data4_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_array_impl_data4_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data4_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_113_12_128_4096_4096_128_1_gen
      weight_mem_banks_bank_array_impl_data5_rsci (
      .clken(weight_mem_banks_bank_array_impl_data5_rsc_clken),
      .q(weight_mem_banks_bank_array_impl_data5_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data5_rsc_radr),
      .we(weight_mem_banks_bank_array_impl_data5_rsc_we),
      .d(weight_mem_banks_bank_array_impl_data5_rsc_d),
      .wadr(weight_mem_banks_bank_array_impl_data5_rsc_wadr),
      .clken_d(weight_mem_banks_bank_array_impl_data5_rsci_clken_d),
      .d_d(weight_mem_banks_bank_array_impl_data5_rsci_d_d),
      .q_d(weight_mem_banks_bank_array_impl_data5_rsci_q_d),
      .radr_d(weight_mem_banks_bank_array_impl_data5_rsci_radr_d),
      .wadr_d(weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_array_impl_data5_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_array_impl_data5_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data5_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_114_12_128_4096_4096_128_1_gen
      weight_mem_banks_bank_array_impl_data6_rsci (
      .clken(weight_mem_banks_bank_array_impl_data6_rsc_clken),
      .q(weight_mem_banks_bank_array_impl_data6_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data6_rsc_radr),
      .we(weight_mem_banks_bank_array_impl_data6_rsc_we),
      .d(weight_mem_banks_bank_array_impl_data6_rsc_d),
      .wadr(weight_mem_banks_bank_array_impl_data6_rsc_wadr),
      .clken_d(weight_mem_banks_bank_array_impl_data6_rsci_clken_d),
      .d_d(weight_mem_banks_bank_array_impl_data6_rsci_d_d),
      .q_d(weight_mem_banks_bank_array_impl_data6_rsci_q_d),
      .radr_d(weight_mem_banks_bank_array_impl_data6_rsci_radr_d),
      .wadr_d(weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_array_impl_data6_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_array_impl_data6_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data6_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_115_12_128_4096_4096_128_1_gen
      weight_mem_banks_bank_array_impl_data7_rsci (
      .clken(weight_mem_banks_bank_array_impl_data7_rsc_clken),
      .q(weight_mem_banks_bank_array_impl_data7_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data7_rsc_radr),
      .we(weight_mem_banks_bank_array_impl_data7_rsc_we),
      .d(weight_mem_banks_bank_array_impl_data7_rsc_d),
      .wadr(weight_mem_banks_bank_array_impl_data7_rsc_wadr),
      .clken_d(weight_mem_banks_bank_array_impl_data7_rsci_clken_d),
      .d_d(weight_mem_banks_bank_array_impl_data7_rsci_d_d),
      .q_d(weight_mem_banks_bank_array_impl_data7_rsci_q_d),
      .radr_d(weight_mem_banks_bank_array_impl_data7_rsci_radr_d),
      .wadr_d(weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_array_impl_data7_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_array_impl_data7_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data7_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_116_12_128_4096_4096_128_1_gen
      weight_mem_banks_bank_array_impl_data8_rsci (
      .clken(weight_mem_banks_bank_array_impl_data8_rsc_clken),
      .q(weight_mem_banks_bank_array_impl_data8_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data8_rsc_radr),
      .we(weight_mem_banks_bank_array_impl_data8_rsc_we),
      .d(weight_mem_banks_bank_array_impl_data8_rsc_d),
      .wadr(weight_mem_banks_bank_array_impl_data8_rsc_wadr),
      .clken_d(weight_mem_banks_bank_array_impl_data8_rsci_clken_d),
      .d_d(weight_mem_banks_bank_array_impl_data8_rsci_d_d),
      .q_d(weight_mem_banks_bank_array_impl_data8_rsci_q_d),
      .radr_d(weight_mem_banks_bank_array_impl_data8_rsci_radr_d),
      .wadr_d(weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_array_impl_data8_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_array_impl_data8_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data8_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_117_12_128_4096_4096_128_1_gen
      weight_mem_banks_bank_array_impl_data9_rsci (
      .clken(weight_mem_banks_bank_array_impl_data9_rsc_clken),
      .q(weight_mem_banks_bank_array_impl_data9_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data9_rsc_radr),
      .we(weight_mem_banks_bank_array_impl_data9_rsc_we),
      .d(weight_mem_banks_bank_array_impl_data9_rsc_d),
      .wadr(weight_mem_banks_bank_array_impl_data9_rsc_wadr),
      .clken_d(weight_mem_banks_bank_array_impl_data9_rsci_clken_d),
      .d_d(weight_mem_banks_bank_array_impl_data9_rsci_d_d),
      .q_d(weight_mem_banks_bank_array_impl_data9_rsci_q_d),
      .radr_d(weight_mem_banks_bank_array_impl_data9_rsci_radr_d),
      .wadr_d(weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_array_impl_data9_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_array_impl_data9_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data9_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_118_12_128_4096_4096_128_1_gen
      weight_mem_banks_bank_array_impl_data10_rsci (
      .clken(weight_mem_banks_bank_array_impl_data10_rsc_clken),
      .q(weight_mem_banks_bank_array_impl_data10_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data10_rsc_radr),
      .we(weight_mem_banks_bank_array_impl_data10_rsc_we),
      .d(weight_mem_banks_bank_array_impl_data10_rsc_d),
      .wadr(weight_mem_banks_bank_array_impl_data10_rsc_wadr),
      .clken_d(weight_mem_banks_bank_array_impl_data10_rsci_clken_d),
      .d_d(weight_mem_banks_bank_array_impl_data10_rsci_d_d),
      .q_d(weight_mem_banks_bank_array_impl_data10_rsci_q_d),
      .radr_d(weight_mem_banks_bank_array_impl_data10_rsci_radr_d),
      .wadr_d(weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_array_impl_data10_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_array_impl_data10_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data10_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_119_12_128_4096_4096_128_1_gen
      weight_mem_banks_bank_array_impl_data11_rsci (
      .clken(weight_mem_banks_bank_array_impl_data11_rsc_clken),
      .q(weight_mem_banks_bank_array_impl_data11_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data11_rsc_radr),
      .we(weight_mem_banks_bank_array_impl_data11_rsc_we),
      .d(weight_mem_banks_bank_array_impl_data11_rsc_d),
      .wadr(weight_mem_banks_bank_array_impl_data11_rsc_wadr),
      .clken_d(weight_mem_banks_bank_array_impl_data11_rsci_clken_d),
      .d_d(weight_mem_banks_bank_array_impl_data11_rsci_d_d),
      .q_d(weight_mem_banks_bank_array_impl_data11_rsci_q_d),
      .radr_d(weight_mem_banks_bank_array_impl_data11_rsci_radr_d),
      .wadr_d(weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_array_impl_data11_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_array_impl_data11_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data11_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_120_12_128_4096_4096_128_1_gen
      weight_mem_banks_bank_array_impl_data12_rsci (
      .clken(weight_mem_banks_bank_array_impl_data12_rsc_clken),
      .q(weight_mem_banks_bank_array_impl_data12_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data12_rsc_radr),
      .we(weight_mem_banks_bank_array_impl_data12_rsc_we),
      .d(weight_mem_banks_bank_array_impl_data12_rsc_d),
      .wadr(weight_mem_banks_bank_array_impl_data12_rsc_wadr),
      .clken_d(weight_mem_banks_bank_array_impl_data12_rsci_clken_d),
      .d_d(weight_mem_banks_bank_array_impl_data12_rsci_d_d),
      .q_d(weight_mem_banks_bank_array_impl_data12_rsci_q_d),
      .radr_d(weight_mem_banks_bank_array_impl_data12_rsci_radr_d),
      .wadr_d(weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_array_impl_data12_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_array_impl_data12_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data12_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_121_12_128_4096_4096_128_1_gen
      weight_mem_banks_bank_array_impl_data13_rsci (
      .clken(weight_mem_banks_bank_array_impl_data13_rsc_clken),
      .q(weight_mem_banks_bank_array_impl_data13_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data13_rsc_radr),
      .we(weight_mem_banks_bank_array_impl_data13_rsc_we),
      .d(weight_mem_banks_bank_array_impl_data13_rsc_d),
      .wadr(weight_mem_banks_bank_array_impl_data13_rsc_wadr),
      .clken_d(weight_mem_banks_bank_array_impl_data13_rsci_clken_d),
      .d_d(weight_mem_banks_bank_array_impl_data13_rsci_d_d),
      .q_d(weight_mem_banks_bank_array_impl_data13_rsci_q_d),
      .radr_d(weight_mem_banks_bank_array_impl_data13_rsci_radr_d),
      .wadr_d(weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_array_impl_data13_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_array_impl_data13_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data13_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_122_12_128_4096_4096_128_1_gen
      weight_mem_banks_bank_array_impl_data14_rsci (
      .clken(weight_mem_banks_bank_array_impl_data14_rsc_clken),
      .q(weight_mem_banks_bank_array_impl_data14_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data14_rsc_radr),
      .we(weight_mem_banks_bank_array_impl_data14_rsc_we),
      .d(weight_mem_banks_bank_array_impl_data14_rsc_d),
      .wadr(weight_mem_banks_bank_array_impl_data14_rsc_wadr),
      .clken_d(weight_mem_banks_bank_array_impl_data14_rsci_clken_d),
      .d_d(weight_mem_banks_bank_array_impl_data14_rsci_d_d),
      .q_d(weight_mem_banks_bank_array_impl_data14_rsci_q_d),
      .radr_d(weight_mem_banks_bank_array_impl_data14_rsci_radr_d),
      .wadr_d(weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_array_impl_data14_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_array_impl_data14_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data14_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_123_12_128_4096_4096_128_1_gen
      weight_mem_banks_bank_array_impl_data15_rsci (
      .clken(weight_mem_banks_bank_array_impl_data15_rsc_clken),
      .q(weight_mem_banks_bank_array_impl_data15_rsc_q),
      .radr(weight_mem_banks_bank_array_impl_data15_rsc_radr),
      .we(weight_mem_banks_bank_array_impl_data15_rsc_we),
      .d(weight_mem_banks_bank_array_impl_data15_rsc_d),
      .wadr(weight_mem_banks_bank_array_impl_data15_rsc_wadr),
      .clken_d(weight_mem_banks_bank_array_impl_data15_rsci_clken_d),
      .d_d(weight_mem_banks_bank_array_impl_data15_rsci_d_d),
      .q_d(weight_mem_banks_bank_array_impl_data15_rsci_q_d),
      .radr_d(weight_mem_banks_bank_array_impl_data15_rsci_radr_d),
      .wadr_d(weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_array_impl_data15_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_array_impl_data15_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data15_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_125_8_128_256_256_128_1_gen
      input_mem_banks_bank_array_impl_data0_rsci (
      .clken(input_mem_banks_bank_array_impl_data0_rsc_clken),
      .q(input_mem_banks_bank_array_impl_data0_rsc_q),
      .radr(input_mem_banks_bank_array_impl_data0_rsc_radr),
      .we(input_mem_banks_bank_array_impl_data0_rsc_we),
      .d(input_mem_banks_bank_array_impl_data0_rsc_d),
      .wadr(input_mem_banks_bank_array_impl_data0_rsc_wadr),
      .clken_d(input_mem_banks_bank_array_impl_data0_rsci_clken_d),
      .d_d(input_mem_banks_bank_array_impl_data0_rsci_d_d),
      .q_d(input_mem_banks_bank_array_impl_data0_rsci_q_d),
      .radr_d(input_mem_banks_bank_array_impl_data0_rsci_radr_d),
      .wadr_d(input_mem_banks_bank_array_impl_data0_rsci_wadr_d),
      .we_d(input_mem_banks_bank_array_impl_data0_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(input_mem_banks_bank_array_impl_data0_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(input_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  PECore_PECore_PECoreRun PECore_PECoreRun_inst (
      .clk(clk),
      .rst(rst),
      .start_val(start_val),
      .start_rdy(start_rdy),
      .start_msg(start_msg),
      .input_port_val(input_port_val),
      .input_port_rdy(input_port_rdy),
      .input_port_msg(input_port_msg),
      .rva_in_val(rva_in_val),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_msg(rva_in_msg),
      .rva_out_val(rva_out_val),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_msg(rva_out_msg),
      .act_port_val(act_port_val),
      .act_port_rdy(act_port_rdy),
      .act_port_msg(act_port_msg),
      .SC_SRAM_CONFIG(SC_SRAM_CONFIG),
      .weight_mem_banks_bank_array_impl_data0_rsci_clken_d(weight_mem_banks_bank_array_impl_data0_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data0_rsci_d_d(weight_mem_banks_bank_array_impl_data0_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data0_rsci_q_d(weight_mem_banks_bank_array_impl_data0_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data0_rsci_radr_d(weight_mem_banks_bank_array_impl_data0_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data1_rsci_clken_d(weight_mem_banks_bank_array_impl_data1_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data1_rsci_d_d(weight_mem_banks_bank_array_impl_data1_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data1_rsci_q_d(weight_mem_banks_bank_array_impl_data1_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data1_rsci_radr_d(weight_mem_banks_bank_array_impl_data1_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data1_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data1_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data2_rsci_clken_d(weight_mem_banks_bank_array_impl_data2_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data2_rsci_d_d(weight_mem_banks_bank_array_impl_data2_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data2_rsci_q_d(weight_mem_banks_bank_array_impl_data2_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data2_rsci_radr_d(weight_mem_banks_bank_array_impl_data2_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data2_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data2_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data3_rsci_clken_d(weight_mem_banks_bank_array_impl_data3_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data3_rsci_d_d(weight_mem_banks_bank_array_impl_data3_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data3_rsci_q_d(weight_mem_banks_bank_array_impl_data3_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data3_rsci_radr_d(weight_mem_banks_bank_array_impl_data3_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data3_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data3_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data4_rsci_clken_d(weight_mem_banks_bank_array_impl_data4_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data4_rsci_d_d(weight_mem_banks_bank_array_impl_data4_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data4_rsci_q_d(weight_mem_banks_bank_array_impl_data4_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data4_rsci_radr_d(weight_mem_banks_bank_array_impl_data4_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data4_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data4_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data5_rsci_clken_d(weight_mem_banks_bank_array_impl_data5_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data5_rsci_d_d(weight_mem_banks_bank_array_impl_data5_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data5_rsci_q_d(weight_mem_banks_bank_array_impl_data5_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data5_rsci_radr_d(weight_mem_banks_bank_array_impl_data5_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data5_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data5_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data6_rsci_clken_d(weight_mem_banks_bank_array_impl_data6_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data6_rsci_d_d(weight_mem_banks_bank_array_impl_data6_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data6_rsci_q_d(weight_mem_banks_bank_array_impl_data6_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data6_rsci_radr_d(weight_mem_banks_bank_array_impl_data6_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data6_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data6_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data7_rsci_clken_d(weight_mem_banks_bank_array_impl_data7_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data7_rsci_d_d(weight_mem_banks_bank_array_impl_data7_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data7_rsci_q_d(weight_mem_banks_bank_array_impl_data7_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data7_rsci_radr_d(weight_mem_banks_bank_array_impl_data7_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data7_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data7_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data8_rsci_clken_d(weight_mem_banks_bank_array_impl_data8_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data8_rsci_d_d(weight_mem_banks_bank_array_impl_data8_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data8_rsci_q_d(weight_mem_banks_bank_array_impl_data8_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data8_rsci_radr_d(weight_mem_banks_bank_array_impl_data8_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data8_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data8_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data9_rsci_clken_d(weight_mem_banks_bank_array_impl_data9_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data9_rsci_d_d(weight_mem_banks_bank_array_impl_data9_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data9_rsci_q_d(weight_mem_banks_bank_array_impl_data9_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data9_rsci_radr_d(weight_mem_banks_bank_array_impl_data9_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data9_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data9_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data10_rsci_clken_d(weight_mem_banks_bank_array_impl_data10_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data10_rsci_d_d(weight_mem_banks_bank_array_impl_data10_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data10_rsci_q_d(weight_mem_banks_bank_array_impl_data10_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data10_rsci_radr_d(weight_mem_banks_bank_array_impl_data10_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data10_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data10_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data11_rsci_clken_d(weight_mem_banks_bank_array_impl_data11_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data11_rsci_d_d(weight_mem_banks_bank_array_impl_data11_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data11_rsci_q_d(weight_mem_banks_bank_array_impl_data11_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data11_rsci_radr_d(weight_mem_banks_bank_array_impl_data11_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data11_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data11_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data12_rsci_clken_d(weight_mem_banks_bank_array_impl_data12_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data12_rsci_d_d(weight_mem_banks_bank_array_impl_data12_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data12_rsci_q_d(weight_mem_banks_bank_array_impl_data12_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data12_rsci_radr_d(weight_mem_banks_bank_array_impl_data12_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data12_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data12_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data13_rsci_clken_d(weight_mem_banks_bank_array_impl_data13_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data13_rsci_d_d(weight_mem_banks_bank_array_impl_data13_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data13_rsci_q_d(weight_mem_banks_bank_array_impl_data13_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data13_rsci_radr_d(weight_mem_banks_bank_array_impl_data13_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data13_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data13_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data14_rsci_clken_d(weight_mem_banks_bank_array_impl_data14_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data14_rsci_d_d(weight_mem_banks_bank_array_impl_data14_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data14_rsci_q_d(weight_mem_banks_bank_array_impl_data14_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data14_rsci_radr_d(weight_mem_banks_bank_array_impl_data14_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data14_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data14_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data15_rsci_clken_d(weight_mem_banks_bank_array_impl_data15_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data15_rsci_d_d(weight_mem_banks_bank_array_impl_data15_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data15_rsci_q_d(weight_mem_banks_bank_array_impl_data15_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data15_rsci_radr_d(weight_mem_banks_bank_array_impl_data15_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data15_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data15_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .input_mem_banks_bank_array_impl_data0_rsci_clken_d(input_mem_banks_bank_array_impl_data0_rsci_clken_d),
      .input_mem_banks_bank_array_impl_data0_rsci_d_d(input_mem_banks_bank_array_impl_data0_rsci_d_d),
      .input_mem_banks_bank_array_impl_data0_rsci_q_d(input_mem_banks_bank_array_impl_data0_rsci_q_d),
      .input_mem_banks_bank_array_impl_data0_rsci_radr_d(input_mem_banks_bank_array_impl_data0_rsci_radr_d),
      .input_mem_banks_bank_array_impl_data0_rsci_wadr_d(input_mem_banks_bank_array_impl_data0_rsci_wadr_d),
      .input_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d(input_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_pff(weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_iff),
      .weight_mem_banks_bank_array_impl_data0_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data0_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data1_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data1_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data2_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data2_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data3_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data3_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data4_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data4_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data5_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data5_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data6_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data6_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data7_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data7_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data8_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data8_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data9_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data9_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data10_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data10_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data11_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data11_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data12_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data12_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data13_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data13_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data14_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data14_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data15_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data15_rsci_we_d_iff),
      .input_mem_banks_bank_array_impl_data0_rsci_we_d_pff(input_mem_banks_bank_array_impl_data0_rsci_we_d_iff)
    );
endmodule
