// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun (
  clk, rst, start_val, start_rdy, start_msg, input_port_val, input_port_rdy, input_port_msg,
      rva_in_val, rva_in_rdy, rva_in_msg, rva_out_val, rva_out_rdy, rva_out_msg,
      act_port_val, act_port_rdy, act_port_msg, SC_SRAM_CONFIG, weight_mem_banks_bank_array_impl_data0_rsci_clken_d,
      weight_mem_banks_bank_array_impl_data0_rsci_d_d, weight_mem_banks_bank_array_impl_data0_rsci_q_d,
      weight_mem_banks_bank_array_impl_data0_rsci_radr_d, weight_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data1_rsci_clken_d, weight_mem_banks_bank_array_impl_data1_rsci_d_d,
      weight_mem_banks_bank_array_impl_data1_rsci_q_d, weight_mem_banks_bank_array_impl_data1_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data1_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data2_rsci_clken_d, weight_mem_banks_bank_array_impl_data2_rsci_d_d,
      weight_mem_banks_bank_array_impl_data2_rsci_q_d, weight_mem_banks_bank_array_impl_data2_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data2_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data3_rsci_clken_d, weight_mem_banks_bank_array_impl_data3_rsci_d_d,
      weight_mem_banks_bank_array_impl_data3_rsci_q_d, weight_mem_banks_bank_array_impl_data3_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data3_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data4_rsci_clken_d, weight_mem_banks_bank_array_impl_data4_rsci_d_d,
      weight_mem_banks_bank_array_impl_data4_rsci_q_d, weight_mem_banks_bank_array_impl_data4_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data4_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data5_rsci_clken_d, weight_mem_banks_bank_array_impl_data5_rsci_d_d,
      weight_mem_banks_bank_array_impl_data5_rsci_q_d, weight_mem_banks_bank_array_impl_data5_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data5_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data6_rsci_clken_d, weight_mem_banks_bank_array_impl_data6_rsci_d_d,
      weight_mem_banks_bank_array_impl_data6_rsci_q_d, weight_mem_banks_bank_array_impl_data6_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data6_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data7_rsci_clken_d, weight_mem_banks_bank_array_impl_data7_rsci_d_d,
      weight_mem_banks_bank_array_impl_data7_rsci_q_d, weight_mem_banks_bank_array_impl_data7_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data7_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data8_rsci_clken_d, weight_mem_banks_bank_array_impl_data8_rsci_d_d,
      weight_mem_banks_bank_array_impl_data8_rsci_q_d, weight_mem_banks_bank_array_impl_data8_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data8_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data9_rsci_clken_d, weight_mem_banks_bank_array_impl_data9_rsci_d_d,
      weight_mem_banks_bank_array_impl_data9_rsci_q_d, weight_mem_banks_bank_array_impl_data9_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data9_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data10_rsci_clken_d, weight_mem_banks_bank_array_impl_data10_rsci_d_d,
      weight_mem_banks_bank_array_impl_data10_rsci_q_d, weight_mem_banks_bank_array_impl_data10_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data10_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data11_rsci_clken_d, weight_mem_banks_bank_array_impl_data11_rsci_d_d,
      weight_mem_banks_bank_array_impl_data11_rsci_q_d, weight_mem_banks_bank_array_impl_data11_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data11_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data12_rsci_clken_d, weight_mem_banks_bank_array_impl_data12_rsci_d_d,
      weight_mem_banks_bank_array_impl_data12_rsci_q_d, weight_mem_banks_bank_array_impl_data12_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data12_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data13_rsci_clken_d, weight_mem_banks_bank_array_impl_data13_rsci_d_d,
      weight_mem_banks_bank_array_impl_data13_rsci_q_d, weight_mem_banks_bank_array_impl_data13_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data13_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data14_rsci_clken_d, weight_mem_banks_bank_array_impl_data14_rsci_d_d,
      weight_mem_banks_bank_array_impl_data14_rsci_q_d, weight_mem_banks_bank_array_impl_data14_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data14_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data15_rsci_clken_d, weight_mem_banks_bank_array_impl_data15_rsci_d_d,
      weight_mem_banks_bank_array_impl_data15_rsci_q_d, weight_mem_banks_bank_array_impl_data15_rsci_radr_d,
      weight_mem_banks_bank_array_impl_data15_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      input_mem_banks_bank_array_impl_data0_rsci_clken_d, input_mem_banks_bank_array_impl_data0_rsci_d_d,
      input_mem_banks_bank_array_impl_data0_rsci_q_d, input_mem_banks_bank_array_impl_data0_rsci_radr_d,
      input_mem_banks_bank_array_impl_data0_rsci_wadr_d, input_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_pff, weight_mem_banks_bank_array_impl_data0_rsci_we_d_pff,
      weight_mem_banks_bank_array_impl_data1_rsci_we_d_pff, weight_mem_banks_bank_array_impl_data2_rsci_we_d_pff,
      weight_mem_banks_bank_array_impl_data3_rsci_we_d_pff, weight_mem_banks_bank_array_impl_data4_rsci_we_d_pff,
      weight_mem_banks_bank_array_impl_data5_rsci_we_d_pff, weight_mem_banks_bank_array_impl_data6_rsci_we_d_pff,
      weight_mem_banks_bank_array_impl_data7_rsci_we_d_pff, weight_mem_banks_bank_array_impl_data8_rsci_we_d_pff,
      weight_mem_banks_bank_array_impl_data9_rsci_we_d_pff, weight_mem_banks_bank_array_impl_data10_rsci_we_d_pff,
      weight_mem_banks_bank_array_impl_data11_rsci_we_d_pff, weight_mem_banks_bank_array_impl_data12_rsci_we_d_pff,
      weight_mem_banks_bank_array_impl_data13_rsci_we_d_pff, weight_mem_banks_bank_array_impl_data14_rsci_we_d_pff,
      weight_mem_banks_bank_array_impl_data15_rsci_we_d_pff, input_mem_banks_bank_array_impl_data0_rsci_we_d_pff
);
  input clk;
  input rst;
  input start_val;
  output start_rdy;
  input start_msg;
  input input_port_val;
  output input_port_rdy;
  input [137:0] input_port_msg;
  input rva_in_val;
  output rva_in_rdy;
  input [168:0] rva_in_msg;
  output rva_out_val;
  input rva_out_rdy;
  output [127:0] rva_out_msg;
  output act_port_val;
  input act_port_rdy;
  output [319:0] act_port_msg;
  input [31:0] SC_SRAM_CONFIG;
  output weight_mem_banks_bank_array_impl_data0_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data0_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data0_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data0_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data1_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data1_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data1_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data1_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data1_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data2_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data2_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data2_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data2_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data2_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data3_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data3_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data3_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data3_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data3_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data4_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data4_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data4_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data4_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data4_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data5_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data5_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data5_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data5_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data5_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data6_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data6_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data6_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data6_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data6_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data7_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data7_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data7_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data7_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data7_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data8_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data8_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data8_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data8_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data8_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data9_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data9_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data9_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data9_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data9_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data10_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data10_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data10_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data10_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data10_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data11_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data11_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data11_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data11_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data11_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data12_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data12_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data12_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data12_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data12_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data13_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data13_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data13_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data13_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data13_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data14_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data14_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data14_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data14_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data14_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output weight_mem_banks_bank_array_impl_data15_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_array_impl_data15_rsci_d_d;
  input [127:0] weight_mem_banks_bank_array_impl_data15_rsci_q_d;
  output [11:0] weight_mem_banks_bank_array_impl_data15_rsci_radr_d;
  output weight_mem_banks_bank_array_impl_data15_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output input_mem_banks_bank_array_impl_data0_rsci_clken_d;
  output [127:0] input_mem_banks_bank_array_impl_data0_rsci_d_d;
  input [127:0] input_mem_banks_bank_array_impl_data0_rsci_q_d;
  output [7:0] input_mem_banks_bank_array_impl_data0_rsci_radr_d;
  output [7:0] input_mem_banks_bank_array_impl_data0_rsci_wadr_d;
  output input_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output [11:0] weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_pff;
  output weight_mem_banks_bank_array_impl_data0_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data1_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data2_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data3_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data4_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data5_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data6_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data7_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data8_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data9_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data10_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data11_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data12_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data13_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data14_rsci_we_d_pff;
  output weight_mem_banks_bank_array_impl_data15_rsci_we_d_pff;
  output input_mem_banks_bank_array_impl_data0_rsci_we_d_pff;


  // Interconnect Declarations
  wire PECoreRun_wen;
  wire PECoreRun_wten;
  wire [136:0] input_port_PopNB_mioi_idat_mxwt;
  wire input_port_PopNB_mioi_ivld_mxwt;
  wire [168:0] rva_in_PopNB_mioi_idat_mxwt;
  wire rva_in_PopNB_mioi_ivld_mxwt;
  wire act_port_Push_mioi_wen_comp;
  wire rva_out_Push_mioi_wen_comp;
  wire start_PopNB_mioi_idat_mxwt;
  wire start_PopNB_mioi_ivld_mxwt;
  wire [31:0] Datapath_for_1_ProductSum_cmp_out_rsc_z;
  wire Datapath_for_1_ProductSum_cmp_ccs_ccore_en;
  wire [31:0] Datapath_for_1_ProductSum_cmp_1_out_rsc_z;
  wire [31:0] Datapath_for_1_ProductSum_cmp_2_out_rsc_z;
  wire [31:0] Datapath_for_1_ProductSum_cmp_3_out_rsc_z;
  wire [12:0] PEManager_16U_GetWeightAddr_if_acc_4_cmp_z;
  reg [19:0] act_port_Push_mioi_idat_319_300;
  reg [19:0] act_port_Push_mioi_idat_299_280;
  reg [19:0] act_port_Push_mioi_idat_279_260;
  reg [19:0] act_port_Push_mioi_idat_259_240;
  reg [19:0] act_port_Push_mioi_idat_239_220;
  reg [19:0] act_port_Push_mioi_idat_219_200;
  reg [19:0] act_port_Push_mioi_idat_199_180;
  reg [19:0] act_port_Push_mioi_idat_179_160;
  reg [19:0] act_port_Push_mioi_idat_159_140;
  reg [19:0] act_port_Push_mioi_idat_139_120;
  reg [19:0] act_port_Push_mioi_idat_119_100;
  reg [19:0] act_port_Push_mioi_idat_99_80;
  reg [19:0] act_port_Push_mioi_idat_79_60;
  reg [19:0] act_port_Push_mioi_idat_59_40;
  reg [19:0] act_port_Push_mioi_idat_39_20;
  reg [19:0] act_port_Push_mioi_idat_19_0;
  reg [7:0] rva_out_Push_mioi_idat_127_120;
  reg [7:0] rva_out_Push_mioi_idat_119_112;
  reg [7:0] rva_out_Push_mioi_idat_111_104;
  reg [7:0] rva_out_Push_mioi_idat_103_96;
  reg [7:0] rva_out_Push_mioi_idat_95_88;
  reg [7:0] rva_out_Push_mioi_idat_87_80;
  reg [7:0] rva_out_Push_mioi_idat_79_72;
  reg [7:0] rva_out_Push_mioi_idat_71_64;
  reg [7:0] rva_out_Push_mioi_idat_63_56;
  reg [7:0] rva_out_Push_mioi_idat_55_48;
  reg [7:0] rva_out_Push_mioi_idat_47_40;
  reg [3:0] rva_out_Push_mioi_idat_39_36;
  reg [3:0] rva_out_Push_mioi_idat_35_32;
  reg [4:0] rva_out_Push_mioi_idat_31_27;
  reg [1:0] rva_out_Push_mioi_idat_26_25;
  reg rva_out_Push_mioi_idat_24;
  reg [4:0] rva_out_Push_mioi_idat_23_19;
  reg [1:0] rva_out_Push_mioi_idat_18_17;
  reg rva_out_Push_mioi_idat_16;
  reg [4:0] rva_out_Push_mioi_idat_15_11;
  reg [1:0] rva_out_Push_mioi_idat_10_9;
  reg rva_out_Push_mioi_idat_8;
  reg [6:0] rva_out_Push_mioi_idat_7_1;
  reg rva_out_Push_mioi_idat_0;
  wire [4:0] fsm_output;
  wire [8:0] operator_16_false_acc_tmp;
  wire [9:0] nl_operator_16_false_acc_tmp;
  wire [8:0] operator_8_false_acc_tmp;
  wire [9:0] nl_operator_8_false_acc_tmp;
  wire [4:0] operator_4_false_acc_tmp;
  wire [5:0] nl_operator_4_false_acc_tmp;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_239_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_238_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_237_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_236_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_235_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_234_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_232_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_231_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_230_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_229_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_228_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_227_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_226_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_225_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_224_tmp;
  wire [15:0] weight_mem_write_arbxbar_xbar_for_lshift_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_16_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_16_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_15_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_15_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_15_Arbiter_16U_Roundrobin_pick_priority_and_4_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_14_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_14_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_14_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_13_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_13_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_13_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_12_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_12_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_12_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_11_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_11_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_11_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_10_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_10_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_10_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_9_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_9_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_9_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_8_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_8_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_8_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_7_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_7_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_7_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_6_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_6_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_6_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_5_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_5_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_5_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_4_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_4_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_4_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_Arbiter_16U_Roundrobin_pick_or_3_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_3_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_3_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_2_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_2_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_1_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_for_3_1_operator_15_false_operator_15_false_operator_15_false_or_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_16_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_2_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_15_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_3_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_14_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_4_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_13_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_5_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_12_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_6_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_11_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_7_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_10_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_8_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_9_lshift_tmp;
  wire [15:0] weight_mem_read_arbxbar_xbar_for_1_lshift_tmp;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_nor_7_tmp;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_nor_9_tmp;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_nor_11_tmp;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_nor_13_tmp;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_nor_15_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_and_233_tmp;
  wire or_tmp_18;
  wire or_tmp_20;
  wire or_dcpl;
  wire or_dcpl_34;
  wire and_dcpl_135;
  wire and_dcpl_210;
  wire and_dcpl_211;
  wire or_tmp_545;
  wire or_dcpl_247;
  wire and_dcpl_414;
  wire or_dcpl_251;
  wire or_tmp_1286;
  wire or_dcpl_285;
  wire or_dcpl_286;
  wire and_dcpl_437;
  wire and_dcpl_439;
  wire or_dcpl_295;
  wire and_dcpl_440;
  wire or_dcpl_300;
  wire or_dcpl_301;
  wire or_dcpl_302;
  wire or_dcpl_306;
  wire or_dcpl_310;
  wire or_dcpl_313;
  wire or_dcpl_327;
  wire or_dcpl_334;
  wire or_dcpl_362;
  wire or_dcpl_363;
  wire or_dcpl_364;
  wire or_dcpl_365;
  wire or_dcpl_369;
  wire and_dcpl_700;
  wire and_dcpl_702;
  wire or_dcpl_370;
  wire and_dcpl_704;
  wire and_dcpl_705;
  wire and_dcpl_706;
  wire and_dcpl_707;
  wire and_dcpl_708;
  wire and_dcpl_709;
  wire or_dcpl_374;
  wire or_dcpl_375;
  wire or_dcpl_378;
  wire and_dcpl_725;
  wire and_dcpl_726;
  wire and_dcpl_733;
  wire and_dcpl_748;
  wire and_dcpl_749;
  wire and_dcpl_756;
  wire and_dcpl_771;
  wire and_dcpl_772;
  wire and_dcpl_779;
  wire and_dcpl_794;
  wire and_dcpl_795;
  wire and_dcpl_802;
  wire and_dcpl_817;
  wire and_dcpl_818;
  wire and_dcpl_825;
  wire and_dcpl_840;
  wire and_dcpl_841;
  wire and_dcpl_848;
  wire and_dcpl_863;
  wire and_dcpl_864;
  wire and_dcpl_871;
  wire and_dcpl_886;
  wire and_dcpl_887;
  wire and_dcpl_894;
  wire and_dcpl_909;
  wire and_dcpl_910;
  wire and_dcpl_917;
  wire and_dcpl_932;
  wire and_dcpl_933;
  wire and_dcpl_939;
  wire and_dcpl_954;
  wire and_dcpl_955;
  wire and_dcpl_962;
  wire and_dcpl_977;
  wire and_dcpl_978;
  wire and_dcpl_985;
  wire and_dcpl_1000;
  wire and_dcpl_1001;
  wire and_dcpl_1008;
  wire and_dcpl_1023;
  wire and_dcpl_1024;
  wire and_dcpl_1029;
  wire and_dcpl_1043;
  wire and_dcpl_1044;
  wire and_dcpl_1051;
  wire and_dcpl_1066;
  wire and_dcpl_1067;
  wire and_dcpl_1074;
  wire or_tmp_1334;
  wire or_tmp_1655;
  wire or_tmp_2232;
  wire or_tmp_2557;
  wire PECore_RunMac_PECore_RunMac_and_2_cse;
  wire PECore_UpdateFSM_switch_lp_nor_6_cse;
  wire and_2164_cse;
  wire and_2907_cse;
  wire and_4616_cse;
  reg PECore_RunMac_nor_tmp;
  reg pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_pe_config_UpdateInputCounter_if_nor_svs;
  reg PECore_RunFSM_switch_lp_equal_tmp;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_1;
  reg PECore_RunFSM_switch_lp_equal_tmp_1;
  reg PECore_RunFSM_switch_lp_equal_tmp_2;
  reg state_2_0_sva_2;
  reg pe_config_is_valid_sva;
  reg is_start_sva;
  reg input_mem_banks_load_store_for_else_and_cse;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_1_lpi_1_dfm;
  reg PECore_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva;
  reg PECore_CheckStart_start_reg_sva;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp;
  reg [168:0] rva_in_PopNB_mio_mrgout_dat_sva;
  reg PECore_DecodeAxiRead_switch_lp_nor_2_itm;
  reg state_2_0_sva_0;
  reg state_2_0_sva_1;
  wire input_mem_banks_load_store_for_else_and_cse_1;
  reg input_read_req_valid_lpi_1_dfm_5;
  reg input_write_req_valid_lpi_1_dfm_5;
  wire pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1;
  wire pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_nor_svs_1;
  wire pe_config_is_zero_first_sva_dfm_4_mx0;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
  wire PECore_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_mx1;
  wire weight_read_ack_15_lpi_1_dfm_15_mx0;
  wire weight_read_ack_14_lpi_1_dfm_15_mx0;
  wire weight_read_ack_13_lpi_1_dfm_15_mx0;
  wire weight_read_ack_12_lpi_1_dfm_15_mx0;
  wire weight_read_ack_11_lpi_1_dfm_15_mx0;
  wire weight_read_ack_10_lpi_1_dfm_15_mx0;
  wire weight_read_ack_8_lpi_1_dfm_15_mx0;
  wire weight_read_ack_7_lpi_1_dfm_15_mx0;
  wire weight_read_ack_6_lpi_1_dfm_15_mx0;
  wire weight_read_ack_5_lpi_1_dfm_15_mx0;
  wire weight_read_ack_4_lpi_1_dfm_15_mx0;
  wire weight_read_ack_3_lpi_1_dfm_15_mx0;
  wire weight_read_ack_2_lpi_1_dfm_15_mx0;
  wire weight_read_ack_1_lpi_1_dfm_15_mx0;
  wire weight_read_ack_0_lpi_1_dfm_15_mx0;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_15_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_2_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_15_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_15_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_15_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_15_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_15_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_15_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_15_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_15_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_15_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_15_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_15_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_2_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_2_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_2_1_sva_1;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_15_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_15_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_15_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_15_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_15_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_15_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_14_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_14_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_14_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_14_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_14_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_14_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_13_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_13_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_13_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_13_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_13_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_13_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_12_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_12_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_12_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_12_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_12_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_12_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_11_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_11_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_11_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_11_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_11_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_11_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_10_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_10_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_10_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_10_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_10_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_10_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_9_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_9_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_9_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_9_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_9_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_9_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_8_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_8_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_8_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_8_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_8_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_8_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_7_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_7_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_7_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_7_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_7_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_7_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_6_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_6_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_6_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_6_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_6_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_6_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_5_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_5_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_5_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_5_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_5_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_5_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_4_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_4_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_4_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_4_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_4_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_4_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_3_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_3_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_3_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_2_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_2_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_2_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_1_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_7_sva;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_3_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_2_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_1_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_31U_Arbiter_16U_Roundrobin_UnrolledMask_nvhls_nvhls_t_5U_nvuint_t_idx_0_1_lpi_1_dfm_mx0;
  wire Arbiter_16U_Roundrobin_pick_priority_27_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_26_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_30_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_29_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_28_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_23_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_22_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_19_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_18_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_21_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_20_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_25_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_24_1_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_0_15_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_14_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_13_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_12_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_11_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_10_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_8_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_7_sva;
  wire [168:0] rva_in_PopNB_mio_mrgout_dat_sva_1;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_6;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_7;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_8;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_5;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_nor_tmp_1;
  wire PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_5;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_31;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_4;
  wire PECore_DecodeAxiRead_switch_lp_nor_tmp_mx0w0;
  wire PECore_RunFSM_switch_lp_equal_tmp_3;
  reg pe_config_is_bias_sva;
  wire PECore_RunFSM_switch_lp_nor_3_cse_1;
  wire PECore_RunFSM_switch_lp_equal_tmp_5;
  wire PECore_RunFSM_switch_lp_equal_tmp_4;
  wire PECore_RunBias_if_for_11_operator_32_true_slc_operator_32_true_acc_13_svs_mx0;
  reg while_and_46_tmp_1;
  wire PECore_RunBias_if_for_10_operator_32_true_slc_operator_32_true_acc_13_svs_mx0;
  wire PECore_RunBias_if_for_7_operator_32_true_slc_operator_32_true_acc_13_svs_mx0;
  wire PECore_RunBias_if_for_6_operator_32_true_slc_operator_32_true_acc_13_svs_mx0;
  wire PECore_RunBias_if_for_2_operator_32_true_slc_operator_32_true_acc_13_svs_mx2;
  wire PECore_RunBias_if_for_12_operator_32_true_slc_operator_32_true_acc_13_svs_mx2;
  wire PECore_RunBias_if_for_1_operator_32_true_slc_operator_32_true_acc_13_svs_mx2;
  wire PECore_RunBias_if_for_16_operator_32_true_slc_operator_32_true_acc_13_svs_mx1;
  wire while_and_48_tmp_1;
  wire PECore_RunBias_if_for_15_operator_32_true_slc_operator_32_true_acc_13_svs_mx1;
  wire PECore_RunBias_if_for_14_operator_32_true_slc_operator_32_true_acc_13_svs_mx1;
  wire PECore_RunBias_if_for_13_operator_32_true_slc_operator_32_true_acc_13_svs_mx1;
  wire weight_read_ack_9_lpi_1_dfm_15_mx0;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_12_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_11_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_10_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_9_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_8_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_7_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_6_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_5_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_4_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_3_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_2_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  reg while_stage_0_2;
  reg while_asn_41_itm_1;
  reg adpfloat_tmp_is_zero_land_11_lpi_1_dfm;
  reg adpfloat_tmp_is_zero_land_11_lpi_1_dfm_st;
  reg adpfloat_tmp_is_zero_land_10_lpi_1_dfm;
  reg adpfloat_tmp_is_zero_land_10_lpi_1_dfm_st;
  reg PECore_UpdateFSM_case_4_is_output_end_pe_config_UpdateManagerCounter_nand_itm;
  reg PECore_UpdateFSM_switch_lp_unequal_tmp;
  reg [127:0] input_mem_banks_read_read_data_lpi_1;
  reg adpfloat_tmp_is_zero_land_7_lpi_1_dfm;
  reg adpfloat_tmp_is_zero_land_7_lpi_1_dfm_st;
  reg adpfloat_tmp_is_zero_land_6_lpi_1_dfm;
  reg adpfloat_tmp_is_zero_land_6_lpi_1_dfm_st;
  reg while_and_29_itm_1;
  reg while_and_30_itm_1;
  reg PECore_RunBias_if_for_14_operator_32_true_slc_operator_32_true_acc_13_svs;
  reg PECore_RunBias_if_for_15_operator_32_true_slc_operator_32_true_acc_13_svs;
  reg PECore_RunBias_if_for_13_operator_32_true_slc_operator_32_true_acc_13_svs;
  reg PECore_RunBias_if_for_16_operator_32_true_slc_operator_32_true_acc_13_svs;
  reg PECore_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva;
  reg w_axi_rsp_lpi_1_dfm_1;
  reg pe_config_is_zero_first_sva;
  reg pe_manager_zero_active_1_sva;
  reg pe_manager_zero_active_0_sva;
  reg pe_config_is_cluster_sva;
  reg [3:0] pe_config_manager_counter_sva;
  reg [15:0] weight_mem_write_arbxbar_xbar_for_empty_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_16_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_15_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_14_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_13_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_12_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_11_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_10_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_9_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_8_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_7_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_6_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_5_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_4_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_3_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_2_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_1_weight_mem_read_arbxbar_xbar_for_3_if_1_operator_16_false_1_or_mdf_sva;
  reg PECore_DecodeAxiRead_case_4_switch_lp_and_2_itm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_15_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_14_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_13_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_12_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_9_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_8_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_7_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_6_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_5_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_4_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_3_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_2_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_for_land_11_lpi_1_dfm;
  wire [31:0] PECore_RunBias_if_accum_vector_out_data_11_lpi_1_dfm_mx2;
  wire [31:0] PECore_RunBias_if_accum_vector_out_data_10_lpi_1_dfm_mx2;
  wire [31:0] PECore_RunBias_if_accum_vector_out_data_7_lpi_1_dfm_mx2;
  wire [31:0] PECore_RunBias_if_accum_vector_out_data_6_lpi_1_dfm_mx2;
  wire pe_config_manager_counter_sva_dfm_4_mx0_0;
  reg PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva;
  wire while_and_71_m1c;
  wire while_and_73_m1c;
  wire while_and_65_m1c;
  wire while_and_79_m1c;
  wire while_and_63_m1c;
  wire while_and_61_m1c;
  wire while_and_59_m1c;
  wire while_and_57_m1c;
  wire while_and_87_m1c;
  wire while_and_85_m1c;
  wire while_and_83_m1c;
  wire while_and_81_m1c;
  reg [19:0] reg_PECore_RunBias_if_accum_vector_out_data_11_lpi_1_dfm_ftd_12;
  reg [19:0] reg_PECore_RunBias_if_accum_vector_out_data_10_lpi_1_dfm_ftd_12;
  reg [19:0] reg_PECore_RunBias_if_accum_vector_out_data_7_lpi_1_dfm_ftd_12;
  reg [19:0] reg_PECore_RunBias_if_accum_vector_out_data_6_lpi_1_dfm_ftd_12;
  wire while_and_67_m1c;
  wire while_and_69_m1c;
  wire while_and_75_m1c;
  wire while_and_77_m1c;
  wire weight_mem_banks_write_if_for_if_mux_cse;
  wire weight_mem_banks_write_if_for_if_mux_1_cse;
  wire weight_mem_banks_read_for_mux_cse;
  wire weight_mem_banks_read_for_mux_1_cse;
  wire weight_mem_banks_write_if_for_if_mux_4_cse;
  wire weight_mem_banks_write_if_for_if_mux_5_cse;
  wire weight_mem_banks_read_for_mux_4_cse;
  wire weight_mem_banks_read_for_mux_5_cse;
  wire weight_mem_banks_write_if_for_if_mux_8_cse;
  wire weight_mem_banks_write_if_for_if_mux_9_cse;
  wire weight_mem_banks_read_for_mux_8_cse;
  wire weight_mem_banks_read_for_mux_9_cse;
  wire weight_mem_banks_write_if_for_if_mux_12_cse;
  wire weight_mem_banks_write_if_for_if_mux_13_cse;
  wire weight_mem_banks_read_for_mux_12_cse;
  wire weight_mem_banks_read_for_mux_13_cse;
  wire weight_mem_banks_write_if_for_if_mux_16_cse;
  wire weight_mem_banks_write_if_for_if_mux_17_cse;
  wire weight_mem_banks_read_for_mux_16_cse;
  wire weight_mem_banks_read_for_mux_17_cse;
  wire weight_mem_banks_write_if_for_if_mux_20_cse;
  wire weight_mem_banks_write_if_for_if_mux_21_cse;
  wire weight_mem_banks_read_for_mux_20_cse;
  wire weight_mem_banks_read_for_mux_21_cse;
  wire weight_mem_banks_write_if_for_if_mux_24_cse;
  wire weight_mem_banks_write_if_for_if_mux_25_cse;
  wire weight_mem_banks_read_for_mux_24_cse;
  wire weight_mem_banks_read_for_mux_25_cse;
  wire weight_mem_banks_write_if_for_if_mux_28_cse;
  wire weight_mem_banks_write_if_for_if_mux_29_cse;
  wire weight_mem_banks_read_for_mux_28_cse;
  wire weight_mem_banks_read_for_mux_29_cse;
  wire weight_mem_banks_write_if_for_if_mux_32_cse;
  wire weight_mem_banks_write_if_for_if_mux_33_cse;
  wire weight_mem_banks_read_for_mux_32_cse;
  wire weight_mem_banks_read_for_mux_33_cse;
  wire weight_mem_banks_write_if_for_if_mux_36_cse;
  wire weight_mem_banks_write_if_for_if_mux_37_cse;
  wire weight_mem_banks_read_for_mux_36_cse;
  wire weight_mem_banks_read_for_mux_37_cse;
  wire weight_mem_banks_write_if_for_if_mux_40_cse;
  wire weight_mem_banks_write_if_for_if_mux_41_cse;
  wire weight_mem_banks_read_for_mux_40_cse;
  wire weight_mem_banks_read_for_mux_41_cse;
  wire weight_mem_banks_write_if_for_if_mux_44_cse;
  wire weight_mem_banks_write_if_for_if_mux_45_cse;
  wire weight_mem_banks_read_for_mux_44_cse;
  wire weight_mem_banks_read_for_mux_45_cse;
  wire weight_mem_banks_write_if_for_if_mux_48_cse;
  wire weight_mem_banks_write_if_for_if_mux_49_cse;
  wire weight_mem_banks_read_for_mux_48_cse;
  wire weight_mem_banks_read_for_mux_49_cse;
  wire weight_mem_banks_write_if_for_if_mux_52_cse;
  wire weight_mem_banks_write_if_for_if_mux_53_cse;
  wire weight_mem_banks_read_for_mux_52_cse;
  wire weight_mem_banks_read_for_mux_53_cse;
  wire weight_mem_banks_write_if_for_if_mux_56_cse;
  wire weight_mem_banks_write_if_for_if_mux_57_cse;
  wire weight_mem_banks_read_for_mux_56_cse;
  wire weight_mem_banks_read_for_mux_57_cse;
  wire weight_mem_banks_write_if_for_if_mux_60_cse;
  wire weight_mem_banks_write_if_for_if_mux_61_cse;
  wire weight_mem_banks_read_for_mux_60_cse;
  wire weight_mem_banks_read_for_mux_61_cse;
  wire input_mem_banks_write_if_for_if_mux_1_cse;
  wire input_mem_banks_write_if_for_if_mux_2_cse;
  wire input_mem_banks_read_for_mux_cse;
  wire input_mem_banks_read_for_mux_1_cse;
  reg reg_input_port_PopNB_mioi_oswt_cse;
  reg reg_rva_in_PopNB_mioi_oswt_cse;
  wire PECore_RunMac_if_and_208_cse;
  wire PECore_RunMac_if_and_209_cse;
  wire PECore_RunMac_if_and_176_cse;
  wire PECore_RunMac_if_and_177_cse;
  wire PECore_RunMac_if_and_144_cse;
  wire PECore_RunMac_if_and_145_cse;
  wire PECore_RunMac_if_and_112_cse;
  wire PECore_RunMac_if_and_113_cse;
  wire PECore_PushAxiRsp_if_and_cse;
  wire PECore_PushAxiRsp_if_and_10_cse;
  wire PECore_PushOutput_if_and_cse;
  reg reg_Datapath_for_1_ProductSum_cmp_cgo_ir_3_cse;
  reg reg_input_mem_banks_bank_array_impl_data0_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data15_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data14_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data13_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data12_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data11_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data10_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data9_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data8_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data7_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data6_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data5_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data4_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data3_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data2_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data1_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_array_impl_data0_rsci_cgo_ir_cse;
  reg reg_start_PopNB_mioi_iswt0_cse;
  reg reg_rva_out_Push_mioi_iswt0_cse;
  reg reg_act_port_Push_mioi_iswt0_cse;
  wire pe_manager_adplfloat_bias_weight_and_cse;
  wire pe_manager_adplfloat_bias_weight_and_1_cse;
  wire pe_manager_cluster_lut_data_and_cse;
  wire pe_manager_cluster_lut_data_and_1_cse;
  wire pe_config_num_output_and_cse;
  wire and_5345_cse;
  wire PECore_RunMac_if_and_12_cse;
  wire PECore_RunMac_if_and_13_cse;
  wire PECore_RunMac_if_and_10_cse;
  wire PECore_RunMac_if_and_11_cse;
  wire or_1405_cse;
  wire or_1409_cse;
  wire or_1413_cse;
  wire or_1417_cse;
  wire or_1421_cse;
  wire or_1425_cse;
  wire or_1429_cse;
  wire or_1433_cse;
  wire or_1437_cse;
  wire or_1441_cse;
  wire or_1445_cse;
  wire or_1449_cse;
  wire or_1453_cse;
  wire or_1457_cse;
  wire or_1461_cse;
  wire or_1465_cse;
  wire or_1183_cse;
  wire [127:0] input_mem_banks_write_if_for_if_mux_cse;
  wire or_500_cse;
  wire and_cse;
  wire and_3039_cse;
  wire and_3035_cse;
  wire and_3031_cse;
  wire and_3027_cse;
  wire and_3023_cse;
  wire and_3019_cse;
  wire and_3015_cse;
  wire and_3011_cse;
  wire and_3007_cse;
  wire and_3003_cse;
  wire and_2999_cse;
  wire and_2995_cse;
  wire and_2991_cse;
  wire and_2987_cse;
  wire and_2983_cse;
  wire and_2979_cse;
  wire nor_499_cse;
  wire and_5335_cse;
  wire or_55_cse;
  wire nand_199_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_450_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_452_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_453_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_454_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_455_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_456_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_457_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_420_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_422_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_423_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_424_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_425_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_426_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_427_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_390_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_392_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_393_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_394_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_395_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_396_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_397_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_360_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_362_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_363_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_364_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_365_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_366_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_367_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_330_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_332_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_333_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_334_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_335_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_336_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_337_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_300_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_302_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_303_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_304_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_305_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_306_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_307_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_270_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_272_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_273_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_274_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_275_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_276_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_277_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_240_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_242_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_243_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_244_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_245_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_246_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_247_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_210_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_212_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_213_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_214_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_215_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_216_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_217_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_180_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_182_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_183_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_184_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_185_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_186_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_187_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_150_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_152_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_153_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_154_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_155_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_156_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_157_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_120_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_122_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_123_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_124_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_125_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_126_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_127_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_90_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_92_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_93_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_94_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_95_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_96_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_97_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_60_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_62_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_63_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_64_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_65_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_66_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_67_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_30_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_32_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_33_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_34_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_35_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_36_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_37_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_2_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_3_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_4_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_5_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_6_cse;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_7_cse;
  wire PECore_PushAxiRsp_if_and_45_cse;
  wire pe_config_is_valid_and_cse;
  wire or_1584_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_1_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_2_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_3_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_4_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_5_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_6_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_7_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_8_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_9_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_10_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_11_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_12_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_13_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_14_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_15_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_16_operator_7_false_operator_7_false_operator_7_false_or_cse;
  wire and_2973_cse;
  wire rva_out_reg_data_and_2_cse;
  wire [7:0] weight_write_data_data_mux1h_14_rmff;
  wire [7:0] weight_write_data_data_mux1h_13_rmff;
  wire [7:0] weight_write_data_data_mux1h_12_rmff;
  wire [7:0] weight_write_data_data_mux1h_11_rmff;
  wire [7:0] weight_write_data_data_mux1h_10_rmff;
  wire [7:0] weight_write_data_data_mux1h_9_rmff;
  wire [7:0] weight_write_data_data_mux1h_8_rmff;
  wire [7:0] weight_write_data_data_mux1h_7_rmff;
  wire [7:0] weight_write_data_data_mux1h_6_rmff;
  wire [7:0] weight_write_data_data_mux1h_5_rmff;
  wire [7:0] weight_write_data_data_mux1h_4_rmff;
  wire [7:0] weight_write_data_data_mux1h_3_rmff;
  wire [7:0] weight_write_data_data_mux1h_2_rmff;
  wire [7:0] weight_write_data_data_mux1h_1_rmff;
  wire [7:0] weight_write_data_data_mux1h_rmff;
  wire [127:0] input_mem_banks_read_read_data_mux_rmff;
  wire or_2419_rmff;
  wire or_2438_rmff;
  wire or_2437_rmff;
  wire or_2436_rmff;
  wire or_2435_rmff;
  wire or_2434_rmff;
  wire or_2433_rmff;
  wire or_2432_rmff;
  wire or_2431_rmff;
  wire or_2430_rmff;
  wire or_2429_rmff;
  wire or_2428_rmff;
  wire or_2427_rmff;
  wire or_2426_rmff;
  wire or_2425_rmff;
  wire or_2424_rmff;
  wire or_2423_rmff;
  wire or_2422_rmff;
  wire or_2421_rmff;
  reg [7:0] pe_config_output_counter_sva;
  reg [7:0] pe_manager_num_input_0_sva;
  reg [7:0] pe_manager_num_input_1_sva;
  reg [7:0] pe_config_input_counter_sva;
  reg [7:0] PECore_RunMac_if_mux_175_itm;
  reg [7:0] pe_manager_cluster_lut_data_0_0_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_1_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_2_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_3_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_4_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_5_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_6_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_7_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_8_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_9_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_10_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_11_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_12_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_13_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_14_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_0_15_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_0_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_1_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_2_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_3_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_4_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_5_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_6_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_7_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_8_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_9_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_10_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_11_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_12_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_13_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_14_sva_dfm_4;
  reg [7:0] pe_manager_cluster_lut_data_1_15_sva_dfm_4;
  wire [7:0] weight_port_read_out_data_7_15_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_15_15_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_15_itm;
  reg [7:0] PECore_RunMac_if_mux_174_itm;
  reg [7:0] weight_port_read_out_data_15_14_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_173_itm;
  wire [7:0] weight_port_read_out_data_7_14_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_15_13_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_13_itm;
  reg [7:0] PECore_RunMac_if_mux_172_itm;
  reg [7:0] weight_port_read_out_data_15_12_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_13_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] rva_out_reg_data_79_72_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_171_itm;
  wire [7:0] weight_port_read_out_data_7_13_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_15_11_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_12_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_170_itm;
  reg [7:0] weight_port_read_out_data_15_10_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_11_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_169_itm;
  wire [7:0] weight_port_read_out_data_7_12_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_15_9_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_10_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_9_itm;
  reg [7:0] PECore_RunMac_if_mux_168_itm;
  reg [7:0] weight_port_read_out_data_15_8_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_9_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_8_itm;
  reg [7:0] PECore_RunMac_if_mux_167_itm;
  wire [7:0] weight_port_read_out_data_7_11_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_15_7_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_8_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_7_itm;
  reg [7:0] PECore_RunMac_if_mux_166_itm;
  reg [7:0] weight_port_read_out_data_15_6_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_7_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_6_itm;
  reg [7:0] PECore_RunMac_if_mux_165_itm;
  wire [7:0] weight_port_read_out_data_7_10_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_15_5_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_6_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_5_itm;
  reg [7:0] PECore_RunMac_if_mux_164_itm;
  reg [7:0] weight_port_read_out_data_15_4_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_5_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_4_itm;
  reg [7:0] PECore_RunMac_if_mux_163_itm;
  wire [7:0] weight_port_read_out_data_7_9_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_15_3_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_4_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_3_itm;
  reg [7:0] PECore_RunMac_if_mux_162_itm;
  reg [7:0] weight_port_read_out_data_15_2_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_3_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_2_itm;
  reg [7:0] PECore_RunMac_if_mux_161_itm;
  wire [7:0] weight_port_read_out_data_7_8_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_15_1_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_2_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_160_itm;
  reg [7:0] weight_port_read_out_data_15_0_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_16_data_in_tmp_operator_for_1_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_itm;
  reg [7:0] PECore_RunMac_if_mux_95_itm;
  wire [7:0] weight_port_read_out_data_6_15_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_13_15_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_191_itm;
  reg [7:0] PECore_RunMac_if_mux_79_itm;
  reg [7:0] PECore_RunMac_if_mux_94_itm;
  reg [7:0] weight_port_read_out_data_13_14_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_190_itm;
  reg [7:0] PECore_RunMac_if_mux_78_itm;
  reg [7:0] PECore_RunMac_if_mux_93_itm;
  wire [7:0] weight_port_read_out_data_6_14_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_13_13_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_15;
  reg [7:0] PECore_RunMac_if_mux_189_itm;
  reg [7:0] PECore_RunMac_if_mux_77_itm;
  reg [7:0] PECore_RunMac_if_mux_92_itm;
  reg [7:0] weight_port_read_out_data_13_12_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_17;
  reg [7:0] PECore_RunMac_if_mux_188_itm;
  reg [7:0] PECore_RunMac_if_mux_76_itm;
  reg [7:0] PECore_RunMac_if_mux_91_itm;
  wire [7:0] weight_port_read_out_data_6_13_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_13_11_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_19;
  reg [7:0] PECore_RunMac_if_mux_187_itm;
  reg [7:0] PECore_RunMac_if_mux_75_itm;
  reg [7:0] PECore_RunMac_if_mux_90_itm;
  reg [7:0] weight_port_read_out_data_13_10_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_21;
  reg [7:0] PECore_RunMac_if_mux_186_itm;
  reg [7:0] PECore_RunMac_if_mux_74_itm;
  reg [7:0] PECore_RunMac_if_mux_89_itm;
  wire [7:0] weight_port_read_out_data_6_12_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_13_9_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_23;
  reg [7:0] PECore_RunMac_if_mux_185_itm;
  reg [7:0] PECore_RunMac_if_mux_73_itm;
  reg [7:0] PECore_RunMac_if_mux_88_itm;
  reg [7:0] weight_port_read_out_data_13_8_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_25;
  reg [7:0] PECore_RunMac_if_mux_184_itm;
  reg [7:0] PECore_RunMac_if_mux_72_itm;
  reg [7:0] PECore_RunMac_if_mux_87_itm;
  wire [7:0] weight_port_read_out_data_6_11_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_13_7_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_27;
  reg [7:0] PECore_RunMac_if_mux_183_itm;
  reg [7:0] PECore_RunMac_if_mux_71_itm;
  reg [7:0] PECore_RunMac_if_mux_86_itm;
  reg [7:0] weight_port_read_out_data_13_6_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_29;
  reg [7:0] PECore_RunMac_if_mux_182_itm;
  reg [7:0] PECore_RunMac_if_mux_70_itm;
  reg [7:0] PECore_RunMac_if_mux_85_itm;
  wire [7:0] weight_port_read_out_data_6_10_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_13_5_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_31;
  reg [7:0] PECore_RunMac_if_mux_181_itm;
  reg [7:0] PECore_RunMac_if_mux_69_itm;
  reg [7:0] PECore_RunMac_if_mux_84_itm;
  reg [7:0] weight_port_read_out_data_13_4_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_33;
  reg [7:0] PECore_RunMac_if_mux_180_itm;
  reg [7:0] PECore_RunMac_if_mux_68_itm;
  reg [7:0] PECore_RunMac_if_mux_83_itm;
  wire [7:0] weight_port_read_out_data_6_9_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_13_3_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_35;
  reg [7:0] PECore_RunMac_if_mux_179_itm;
  reg [7:0] PECore_RunMac_if_mux_67_itm;
  reg [7:0] PECore_RunMac_if_mux_82_itm;
  reg [7:0] weight_port_read_out_data_13_2_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_37;
  reg [7:0] PECore_RunMac_if_mux_178_itm;
  reg [7:0] PECore_RunMac_if_mux_66_itm;
  reg [7:0] PECore_RunMac_if_mux_81_itm;
  wire [7:0] weight_port_read_out_data_6_8_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_13_1_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_39;
  reg [7:0] PECore_RunMac_if_mux_177_itm;
  reg [7:0] PECore_RunMac_if_mux_65_itm;
  reg [7:0] PECore_RunMac_if_mux_80_itm;
  reg [7:0] weight_port_read_out_data_13_0_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_14_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_41;
  reg [7:0] PECore_RunMac_if_mux_176_itm;
  reg [7:0] PECore_RunMac_if_mux_64_itm;
  reg [7:0] PECore_RunMac_if_mux_111_itm;
  wire [7:0] weight_port_read_out_data_7_7_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_14_15_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_63_itm;
  reg [7:0] PECore_RunMac_if_mux_110_itm;
  reg [7:0] weight_port_read_out_data_14_14_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_62_itm;
  reg [7:0] PECore_RunMac_if_mux_109_itm;
  wire [7:0] weight_port_read_out_data_7_6_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_14_13_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_14_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_61_itm;
  reg [7:0] PECore_RunMac_if_mux_108_itm;
  reg [7:0] weight_port_read_out_data_14_12_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_13_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_60_itm;
  reg [7:0] PECore_RunMac_if_mux_107_itm;
  wire [7:0] weight_port_read_out_data_7_5_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_14_11_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_12_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_59_itm;
  reg [7:0] PECore_RunMac_if_mux_106_itm;
  reg [7:0] weight_port_read_out_data_14_10_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_11_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_58_itm;
  reg [7:0] PECore_RunMac_if_mux_105_itm;
  wire [7:0] weight_port_read_out_data_7_4_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_14_9_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_10_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_57_itm;
  reg [7:0] weight_port_read_out_data_14_8_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_9_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_136_itm;
  reg [7:0] PECore_RunMac_if_mux_56_itm;
  wire [7:0] weight_port_read_out_data_7_3_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_14_7_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_8_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_135_itm;
  reg [7:0] PECore_RunMac_if_mux_55_itm;
  reg [7:0] weight_port_read_out_data_14_6_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_7_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_134_itm;
  reg [7:0] PECore_RunMac_if_mux_54_itm;
  wire [7:0] weight_port_read_out_data_7_2_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_14_5_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_6_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_133_itm;
  reg [7:0] PECore_RunMac_if_mux_53_itm;
  reg [7:0] weight_port_read_out_data_14_4_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_5_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_132_itm;
  reg [7:0] PECore_RunMac_if_mux_52_itm;
  reg [7:0] PECore_RunMac_if_mux_99_itm;
  wire [7:0] weight_port_read_out_data_7_1_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_14_3_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_4_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_131_itm;
  reg [7:0] PECore_RunMac_if_mux_51_itm;
  reg [7:0] PECore_RunMac_if_mux_98_itm;
  reg [7:0] weight_port_read_out_data_14_2_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_3_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_130_itm;
  reg [7:0] PECore_RunMac_if_mux_50_itm;
  reg [7:0] PECore_RunMac_if_mux_97_itm;
  wire [7:0] weight_port_read_out_data_7_0_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_14_1_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_2_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_49_itm;
  reg [7:0] PECore_RunMac_if_mux_96_itm;
  reg [7:0] weight_port_read_out_data_14_0_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_15_data_in_tmp_operator_for_1_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  reg [7:0] PECore_RunMac_if_mux_48_itm;
  reg [7:0] PECore_RunMac_if_mux_159_itm;
  wire [7:0] weight_port_read_out_data_6_7_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_12_15_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1;
  reg [7:0] PECore_RunMac_if_mux_47_itm;
  reg [7:0] PECore_RunMac_if_mux_158_itm;
  reg [7:0] weight_port_read_out_data_12_14_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1;
  reg [7:0] PECore_RunMac_if_mux_46_itm;
  reg [7:0] PECore_RunMac_if_mux_157_itm;
  wire [7:0] weight_port_read_out_data_6_6_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_12_13_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1;
  reg [7:0] PECore_RunMac_if_mux_45_itm;
  reg [7:0] PECore_RunMac_if_mux_156_itm;
  reg [7:0] weight_port_read_out_data_12_12_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1;
  reg [7:0] PECore_RunMac_if_mux_44_itm;
  reg [7:0] PECore_RunMac_if_mux_155_itm;
  wire [7:0] weight_port_read_out_data_6_5_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_12_11_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1;
  reg [7:0] PECore_RunMac_if_mux_43_itm;
  reg [7:0] PECore_RunMac_if_mux_154_itm;
  reg [7:0] weight_port_read_out_data_12_10_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1;
  reg [7:0] PECore_RunMac_if_mux_42_itm;
  reg [7:0] PECore_RunMac_if_mux_153_itm;
  wire [7:0] weight_port_read_out_data_6_4_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_12_9_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1;
  reg [7:0] rva_out_reg_data_95_88_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_41_itm;
  reg [7:0] PECore_RunMac_if_mux_152_itm;
  reg [7:0] weight_port_read_out_data_12_8_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1;
  reg [7:0] rva_out_reg_data_87_80_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_40_itm;
  reg [7:0] PECore_RunMac_if_mux_151_itm;
  wire [7:0] weight_port_read_out_data_6_3_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_12_7_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1;
  reg [7:0] rva_out_reg_data_71_64_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_39_itm;
  reg [7:0] PECore_RunMac_if_mux_150_itm;
  reg [7:0] weight_port_read_out_data_12_6_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1;
  reg [7:0] rva_out_reg_data_63_56_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_38_itm;
  reg [7:0] PECore_RunMac_if_mux_149_itm;
  wire [7:0] weight_port_read_out_data_6_2_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_12_5_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_37_itm;
  reg [7:0] PECore_RunMac_if_mux_148_itm;
  reg [7:0] weight_port_read_out_data_12_4_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1;
  reg [7:0] rva_out_reg_data_47_40_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_36_itm;
  reg [7:0] PECore_RunMac_if_mux_147_itm;
  wire [7:0] weight_port_read_out_data_6_1_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_12_3_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1;
  reg [7:0] rva_out_reg_data_127_120_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_35_itm;
  reg [7:0] PECore_RunMac_if_mux_146_itm;
  reg [7:0] weight_port_read_out_data_12_2_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1;
  reg [7:0] rva_out_reg_data_119_112_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_34_itm;
  reg [7:0] PECore_RunMac_if_mux_145_itm;
  wire [7:0] weight_port_read_out_data_6_0_sva_dfm_mx1;
  reg [7:0] weight_port_read_out_data_12_1_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1;
  reg [7:0] rva_out_reg_data_111_104_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_33_itm;
  reg [7:0] PECore_RunMac_if_mux_144_itm;
  reg [7:0] weight_port_read_out_data_12_0_sva_dfm;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_13_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1;
  reg [7:0] rva_out_reg_data_103_96_sva_dfm_4;
  reg [7:0] PECore_RunMac_if_mux_32_itm;
  wire while_and_127_cse_1;
  wire [11:0] weight_read_addrs_0_15_4_lpi_1_dfm_5_mx0;
  wire [15:0] weight_read_addrs_1_lpi_1_dfm_2;
  wire [14:0] weight_read_addrs_2_15_1_lpi_1_dfm_2;
  wire [15:0] weight_read_addrs_3_lpi_1_dfm_2;
  wire [13:0] weight_read_addrs_4_15_2_lpi_1_dfm_2;
  wire [15:0] weight_read_addrs_5_lpi_1_dfm_2;
  wire [14:0] weight_read_addrs_6_15_1_lpi_1_dfm_2;
  wire [15:0] weight_read_addrs_7_lpi_1_dfm_2;
  wire [12:0] weight_read_addrs_8_15_3_lpi_1_dfm_3;
  wire [15:0] weight_read_addrs_9_lpi_1_dfm_3;
  wire [14:0] weight_read_addrs_10_15_1_lpi_1_dfm_3;
  wire [15:0] weight_read_addrs_11_lpi_1_dfm_3;
  wire [13:0] weight_read_addrs_12_15_2_lpi_1_dfm_3;
  wire [15:0] weight_read_addrs_13_lpi_1_dfm_3;
  wire [14:0] weight_read_addrs_14_15_1_lpi_1_dfm_3;
  wire [15:0] weight_read_addrs_15_lpi_1_dfm_3;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_3_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_3_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_3_0_sva_1;
  wire [15:0] weight_write_addrs_lpi_1_dfm_6;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_4_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_4_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_4_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_5_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_5_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_5_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_6_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_6_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_6_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_7_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_7_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_7_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_8_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_8_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_8_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_9_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_9_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_9_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_10_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_10_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_10_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_11_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_11_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_11_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_12_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_12_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_12_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_13_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_13_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_13_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_14_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_14_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_14_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_15_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_15_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_15_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_16_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_16_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_16_0_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_17_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_17_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_17_0_sva_1;
  reg [15:0] pe_manager_base_input_0_sva;
  reg [15:0] pe_manager_base_input_1_sva;
  reg [15:0] pe_manager_base_bias_0_sva;
  reg [15:0] pe_manager_base_bias_1_sva;
  wire or_dcpl_717;
  wire or_dcpl_718;
  wire or_dcpl_724;
  reg [31:0] PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_11_sva;
  reg [31:0] PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_1_sva;
  reg [31:0] PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_5_sva;
  reg [31:0] PECore_RunBias_if_for_PECore_RunBias_if_for_rshift_1_cse_4_sva;
  wire PECore_DecodeAxiRead_switch_lp_nor_10_cse_1;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_5;
  reg [7:0] weight_port_read_out_data_0_0_sva_dfm;
  reg [31:0] accum_vector_data_4_sva;
  reg [31:0] accum_vector_data_3_sva;
  reg [31:0] accum_vector_data_2_sva;
  reg [19:0] act_port_reg_data_10_sva;
  reg [19:0] act_port_reg_data_9_sva;
  reg [19:0] act_port_reg_data_6_sva;
  reg [19:0] act_port_reg_data_5_sva;
  reg [31:0] accum_vector_data_9_sva;
  reg [31:0] accum_vector_data_6_sva;
  reg [31:0] accum_vector_data_5_sva;
  reg [31:0] PECore_RunBias_if_accum_vector_out_data_14_lpi_1_dfm;
  reg [31:0] PECore_RunBias_if_accum_vector_out_data_15_lpi_1_dfm;
  wire and_tmp;
  wire PECore_PushAxiRsp_if_asn_70;
  wire and_5501_cse;
  wire and_5502_cse;
  wire or_1593_cse;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_or_6_cse_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_6_sva_1;
  wire [7:0] while_while_and_18_itm;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_3;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_4;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_5;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_6;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_7;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_8;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_9;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_10;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_11;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_12;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_13;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_14;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_2_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_6_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_14_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_1_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_5_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_13_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_0_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_4_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_12_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_1_3_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_3_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_11_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_2_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_10_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_1_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_9_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_0_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_8_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_2_7_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_7_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_6_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_5_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_4_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_3_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_2_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_1_15;
  wire Arbiter_16U_Roundrobin_pick_if_1_and_stg_3_0_15;
  wire [4:0] z_out_4;
  wire [5:0] nl_z_out_4;
  wire [7:0] z_out_5;
  wire [8:0] nl_z_out_5;
  wire [19:0] z_out_17;
  wire [20:0] nl_z_out_17;
  wire [19:0] z_out_18;
  wire [20:0] nl_z_out_18;
  wire [19:0] z_out_19;
  wire [20:0] nl_z_out_19;
  wire [19:0] z_out_20;
  wire [20:0] nl_z_out_20;
  wire [31:0] z_out_25;
  wire [32:0] nl_z_out_25;
  wire [31:0] z_out_26;
  wire [32:0] nl_z_out_26;
  wire [31:0] z_out_27;
  wire [32:0] nl_z_out_27;
  wire [31:0] z_out_28;
  wire [32:0] nl_z_out_28;
  wire [31:0] z_out_29;
  wire [32:0] nl_z_out_29;
  wire [31:0] z_out_30;
  wire [32:0] nl_z_out_30;
  wire [31:0] z_out_31;
  wire [32:0] nl_z_out_31;
  wire [31:0] z_out_32;
  wire [32:0] nl_z_out_32;
  wire [31:0] z_out_37;
  wire [31:0] z_out_38;
  wire [31:0] z_out_39;
  wire [31:0] z_out_40;
  wire or_tmp_3038;
  wire [7:0] z_out_41;
  wire [19:0] z_out_43;
  wire [19:0] z_out_44;
  wire [19:0] z_out_45;
  wire [19:0] z_out_46;
  wire [19:0] z_out_47;
  wire [19:0] z_out_48;
  wire [19:0] z_out_49;
  wire [3:0] z_out_50;
  wire [4:0] nl_z_out_50;
  reg weight_mem_read_arbxbar_arbiters_next_7_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_8_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_9_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_10_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_11_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_12_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_13_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_9_sva;
  reg weight_mem_read_arbxbar_arbiters_next_14_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_15_1_sva;
  reg [2:0] pe_manager_adplfloat_bias_weight_0_sva;
  reg [2:0] pe_manager_adplfloat_bias_weight_1_sva;
  reg [2:0] pe_manager_adplfloat_bias_bias_0_sva;
  reg [2:0] pe_manager_adplfloat_bias_bias_1_sva;
  reg [2:0] pe_manager_adplfloat_bias_input_0_sva;
  reg [2:0] pe_manager_adplfloat_bias_input_1_sva;
  reg [15:0] pe_manager_base_weight_0_sva;
  reg [15:0] pe_manager_base_weight_1_sva;
  reg [3:0] pe_config_num_manager_sva;
  reg [7:0] pe_config_num_output_sva;
  reg [31:0] accum_vector_data_0_sva;
  reg [31:0] accum_vector_data_1_sva;
  reg [31:0] accum_vector_data_10_sva;
  reg [31:0] accum_vector_data_11_sva;
  reg [31:0] accum_vector_data_7_sva;
  reg [31:0] accum_vector_data_8_sva;
  reg [31:0] accum_vector_data_12_sva;
  reg [31:0] accum_vector_data_13_sva;
  reg [31:0] accum_vector_data_14_sva;
  reg [31:0] accum_vector_data_15_sva;
  reg [19:0] act_port_reg_data_7_sva;
  reg [19:0] act_port_reg_data_8_sva;
  reg [19:0] act_port_reg_data_4_sva;
  reg [19:0] act_port_reg_data_11_sva;
  reg [19:0] act_port_reg_data_3_sva;
  reg [19:0] act_port_reg_data_12_sva;
  reg [19:0] act_port_reg_data_2_sva;
  reg [19:0] act_port_reg_data_13_sva;
  reg [19:0] act_port_reg_data_1_sva;
  reg [19:0] act_port_reg_data_14_sva;
  reg [19:0] act_port_reg_data_0_sva;
  reg [19:0] act_port_reg_data_15_sva;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm;
  reg weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm;
  reg crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm;
  reg [7:0] weight_port_read_out_data_0_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_0_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_1_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_2_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_3_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_4_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_5_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_6_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_7_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_8_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_9_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_10_15_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_0_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_1_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_2_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_3_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_4_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_5_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_6_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_7_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_8_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_9_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_10_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_11_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_12_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_13_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_14_sva_dfm;
  reg [7:0] weight_port_read_out_data_11_15_sva_dfm;
  reg PECore_RunBias_if_for_1_operator_32_true_slc_operator_32_true_acc_13_svs;
  reg PECore_RunBias_if_for_2_operator_32_true_slc_operator_32_true_acc_13_svs;
  reg PECore_RunBias_if_for_12_operator_32_true_slc_operator_32_true_acc_13_svs;
  reg [31:0] PECore_RunBias_if_accum_vector_out_data_13_lpi_1_dfm;
  reg [31:0] PECore_RunBias_if_accum_vector_out_data_lpi_1_dfm;
  reg PECore_DecodeAxiRead_case_4_switch_lp_and_itm;
  reg PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm;
  reg PECore_DecodeAxiRead_case_4_switch_lp_and_5_itm;
  reg [7:0] PECore_RunMac_if_mux_31_itm;
  reg [7:0] PECore_RunMac_if_mux_30_itm;
  reg [7:0] PECore_RunMac_if_mux_29_itm;
  reg [7:0] PECore_RunMac_if_mux_28_itm;
  reg [7:0] PECore_RunMac_if_mux_27_itm;
  reg [7:0] PECore_RunMac_if_mux_26_itm;
  reg [7:0] PECore_RunMac_if_mux_25_itm;
  reg [7:0] PECore_RunMac_if_mux_24_itm;
  reg [7:0] PECore_RunMac_if_mux_23_itm;
  reg [7:0] PECore_RunMac_if_mux_22_itm;
  reg [7:0] PECore_RunMac_if_mux_21_itm;
  reg [7:0] PECore_RunMac_if_mux_20_itm;
  reg [7:0] PECore_RunMac_if_mux_19_itm;
  reg [7:0] PECore_RunMac_if_mux_18_itm;
  reg [7:0] PECore_RunMac_if_mux_17_itm;
  reg [7:0] PECore_RunMac_if_mux_16_itm;
  reg PECore_RunBias_if_for_6_operator_4_false_slc_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_0_itm;
  reg PECore_RunBias_if_for_7_operator_4_false_slc_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_0_itm;
  reg PECore_RunBias_if_for_10_operator_4_false_slc_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_0_itm;
  reg PECore_RunBias_if_for_11_operator_4_false_slc_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_0_itm;
  reg [19:0] act_port_reg_data_asn_itm;
  reg [19:0] act_port_reg_data_asn_1_itm;
  reg [19:0] act_port_reg_data_asn_2_itm;
  reg [19:0] act_port_reg_data_asn_3_itm;
  reg pe_manager_cluster_lut_data_1_0_sva_0;
  reg pe_manager_cluster_lut_data_1_1_sva_0;
  reg pe_manager_cluster_lut_data_1_2_sva_0;
  reg pe_manager_cluster_lut_data_1_3_sva_0;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  wire [7:0] weight_port_read_out_data_5_8_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_9_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_10_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_11_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_12_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_13_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_14_sva_dfm_mx1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  wire [7:0] weight_port_read_out_data_5_15_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_0_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_1_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_2_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_3_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_4_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_5_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_6_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_7_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_8_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_9_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_10_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_11_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_12_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_13_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_14_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_4_15_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_8_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_9_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_10_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_11_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_12_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_13_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_14_sva_dfm_mx1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  wire [7:0] weight_port_read_out_data_3_15_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_0_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_1_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_2_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_3_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_4_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_5_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_6_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_3_7_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_0_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_1_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_2_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_3_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_4_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_5_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_6_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_7_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_8_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_9_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_10_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_11_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_12_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_13_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_14_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_2_15_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_8_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_9_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_10_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_11_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_12_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_13_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_14_sva_dfm_mx1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  wire [7:0] weight_port_read_out_data_1_15_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_0_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_1_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_2_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_3_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_4_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_5_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_6_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_1_7_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_8_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_9_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_10_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_11_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_12_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_13_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_14_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_15_sva_dfm_mx1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_1_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  wire [7:0] weight_port_read_out_data_0_0_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_1_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_2_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_3_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_4_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_5_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_6_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_0_7_sva_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_3_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_4_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_5_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_6_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_7_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_8_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_9_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_10_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_11_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_12_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_13_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_14_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_15_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_16_3_lpi_1_dfm_mx1;
  wire weight_mem_read_arbxbar_xbar_for_3_source_local_17_3_lpi_1_dfm_mx1;
  wire adpfloat_tmp_is_zero_land_11_lpi_1_dfm_mx1w0;
  wire adpfloat_tmp_is_zero_land_10_lpi_1_dfm_mx1w0;
  wire adpfloat_tmp_is_zero_land_7_lpi_1_dfm_mx1w0;
  wire adpfloat_tmp_is_zero_land_6_lpi_1_dfm_mx1w0;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_mx0w1;
  wire [7:0] weight_port_read_out_data_5_0_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_1_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_2_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_3_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_4_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_5_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_6_sva_dfm_mx1;
  wire [7:0] weight_port_read_out_data_5_7_sva_dfm_mx1;
  wire while_and_32_cse_1;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_0_lpi_1_dfm_1;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_0_lpi_1_dfm_1;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_0_lpi_1_dfm_1;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_3_lpi_1_dfm_1;
  wire input_read_req_valid_lpi_1_dfm_6;
  wire PECore_DecodeAxiRead_switch_lp_nor_2_itm_mx0w0;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_13_cse_1;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_12_cse_1;
  wire PECore_DecodeAxiRead_switch_lp_nor_14_cse_1;
  wire [12:0] PEManager_16U_GetWeightAddr_if_acc_2_psp_sva_1;
  wire [13:0] nl_PEManager_16U_GetWeightAddr_if_acc_2_psp_sva_1;
  wire [15:0] PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx1;
  wire [11:0] PEManager_16U_GetWeightAddr_1_else_acc_2_psp_sva_1;
  wire [12:0] nl_PEManager_16U_GetWeightAddr_1_else_acc_2_psp_sva_1;
  wire [2:0] weight_read_addrs_8_2_0_lpi_1_dfm_1;
  wire [3:0] while_asn_294_mx0w0;
  wire [3:0] pe_config_manager_counter_sva_dfm_4_mx1;
  wire [7:0] pe_config_input_counter_sva_dfm_4_mx0;
  wire [7:0] pe_config_output_counter_sva_dfm_4_mx0;
  wire [1:0] weight_read_addrs_4_1_0_lpi_1_dfm_1;
  wire weight_read_addrs_0_2_0_lpi_1_dfm_4_2_mx0;
  wire weight_read_addrs_0_2_0_lpi_1_dfm_4_1_mx0;
  wire weight_read_addrs_0_2_0_lpi_1_dfm_4_0_mx0;
  wire weight_read_addrs_0_3_lpi_1_dfm_6;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_0_14_sva_1;
  wire weight_read_addrs_0_3_lpi_1_dfm_5_mx0;
  wire weight_mem_run_1_if_for_land_1_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_2_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_3_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_4_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_5_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_6_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_7_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_8_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_9_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_10_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_11_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_12_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_13_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_14_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_land_15_lpi_1_dfm_1;
  wire weight_read_req_valid_0_lpi_1_dfm_4_mx0;
  wire Arbiter_16U_Roundrobin_pick_return_0_1_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_2_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_3_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_4_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_5_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_6_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_7_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_8_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_9_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_10_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_11_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_12_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_13_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_14_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_15_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_return_0_lpi_1_dfm_2;
  wire input_write_req_valid_lpi_1_dfm_6;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_1_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_1_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_1_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_1_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_1_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_1_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_1_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_1_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_2_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_2_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_2_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_2_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_2_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_2_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_2_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_2_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_3_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_3_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_3_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_3_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_3_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_3_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_3_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_3_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_4_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_4_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_4_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_4_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_4_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_4_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_4_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_4_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_5_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_5_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_5_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_5_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_5_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_5_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_5_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_5_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_6_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_6_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_6_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_6_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_6_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_6_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_6_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_7_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_7_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_7_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_7_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_7_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_7_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_7_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_7_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_8_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_8_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_8_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_8_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_8_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_8_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_8_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_8_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_8_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_8_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_8_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_9_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_9_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_9_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_9_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_9_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_9_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_9_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_9_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_9_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_9_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_9_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_10_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_10_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_10_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_10_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_10_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_10_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_10_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_10_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_10_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_10_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_10_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_11_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_11_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_11_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_11_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_11_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_11_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_11_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_11_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_11_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_11_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_11_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_12_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_12_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_12_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_12_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_12_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_12_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_12_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_12_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_12_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_12_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_12_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_13_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_13_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_13_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_13_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_13_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_13_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_13_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_13_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_13_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_13_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_13_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_14_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_14_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_14_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_14_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_14_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_14_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_14_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_14_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_14_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_14_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_14_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_15_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_15_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_15_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_15_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_15_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_15_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_15_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_15_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_15_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_15_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_15_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_sva_1;
  wire operator_3_false_operator_3_false_operator_3_false_or_mdf_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_sva_1;
  wire Arbiter_16U_Roundrobin_pick_priority_17_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_sva_1;
  wire operator_4_false_operator_4_false_operator_4_false_or_mdf_sva_1;
  wire operator_2_false_3_operator_2_false_3_operator_2_false_3_or_mdf_sva_1;
  wire operator_2_false_4_operator_2_false_4_operator_2_false_4_or_mdf_sva_1;
  wire operator_4_false_1_operator_4_false_1_operator_4_false_1_or_mdf_sva_1;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_mdf_sva_1;
  wire operator_2_false_6_operator_2_false_6_operator_2_false_6_or_mdf_sva_1;
  wire operator_4_false_2_operator_4_false_2_operator_4_false_2_or_mdf_sva_1;
  wire [3:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_lpi_1_dfm_1;
  wire [3:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_14_lpi_1_dfm_1;
  wire [1:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_13_3_2_lpi_1_dfm_1;
  wire [1:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_13_1_0_lpi_1_dfm_1;
  wire [3:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_12_lpi_1_dfm_1;
  wire [2:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_11_3_1_lpi_1_dfm_1;
  wire [2:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_9_2_0_lpi_1_dfm_1;
  wire [3:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_8_lpi_1_dfm_1;
  wire [2:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_7_3_1_lpi_1_dfm_1;
  wire [3:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_6_lpi_1_dfm_1;
  wire [1:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_5_3_2_lpi_1_dfm_1;
  wire [1:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_5_1_0_lpi_1_dfm_1;
  wire [3:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_4_lpi_1_dfm_1;
  wire [2:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_3_3_1_lpi_1_dfm_1;
  wire [3:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_2_lpi_1_dfm_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_1_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_2_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_3_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_4_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_5_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_6_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_7_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_8_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_9_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_10_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_11_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_12_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_13_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_1_14_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_2_14_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_3_14_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_4_14_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_5_14_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_6_14_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_2_7_14_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_0_14_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_1_14_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_2_14_sva_1;
  wire weight_mem_run_1_if_for_if_and_stg_1_3_14_sva_1;
  wire pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_pe_config_UpdateInputCounter_if_nor_svs_1;
  wire PECore_UpdateFSM_switch_lp_unequal_tmp_1;
  wire weight_read_req_valid_8_lpi_1_dfm_1;
  wire weight_read_addrs_10_0_lpi_1_dfm_2;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_8_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_9_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_10_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_11_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_12_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_13_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_14_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_15_sva_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_if_for_13_Arbiter_16U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire [3:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_10_lpi_1_dfm_1;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_241;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_243;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_245;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_247;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_249;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_251;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_253;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_255;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_257;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_259;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_261;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_263;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_265;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_267;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_269;
  wire Arbiter_16U_Roundrobin_pick_if_1_not_271;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_1_sva_mx0w2;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_1_sva_mx0w2;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_12_sva_mx0w1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_12_sva_mx0w1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_2_sva_mx0w1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_2_sva_mx0w1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_3_sva_mx0w1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_3_sva_mx0w1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_4_sva_mx0w1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_4_sva_mx0w1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_5_sva_mx0w1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_5_sva_mx0w1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_8_sva_mx0w1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_8_sva_mx0w1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_9_sva_mx0w1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_9_sva_mx0w1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_12_mx1w2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_11_mx1w2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_13_mx1w2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_3_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_0_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_0_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_1_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_1_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_2_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_2_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_3_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_3_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_4_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_4_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_5_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_5_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_6_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_6_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_7_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_7_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_8_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_8_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_9_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_9_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_10_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_10_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_11_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_11_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_12_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_12_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_13_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_13_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_14_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_14_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_0_15_lpi_1_dfm_2;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_1_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_2_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_3_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_4_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_5_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_6_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_7_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_8_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_9_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_10_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_11_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_12_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_13_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_14_15_lpi_1_dfm_3;
  wire [7:0] weight_mem_run_1_bankread_rsp_rdata_data_15_15_lpi_1_dfm_3;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_5_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_7_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_9_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1;
  wire [3:0] operator_4_false_acc_psp_1_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_1_sva_1;
  wire [3:0] operator_4_false_acc_psp_2_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_2_sva_1;
  wire [3:0] operator_4_false_acc_psp_3_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_3_sva_1;
  wire [3:0] operator_4_false_acc_psp_4_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_4_sva_1;
  wire [3:0] operator_4_false_acc_psp_5_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_5_sva_1;
  wire [3:0] operator_4_false_acc_psp_8_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_8_sva_1;
  wire [3:0] operator_4_false_acc_psp_9_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_9_sva_1;
  wire [3:0] operator_4_false_acc_psp_12_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_12_sva_1;
  wire [3:0] operator_4_false_acc_psp_13_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_13_sva_1;
  wire [3:0] operator_4_false_acc_psp_14_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_14_sva_1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_14_sva_1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_14_sva_1;
  wire [3:0] operator_4_false_acc_psp_15_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_15_sva_1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_15_sva_1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_15_sva_1;
  wire [3:0] operator_4_false_acc_psp_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_sva_1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_sva_1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_sva_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_1_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_12_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_8_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_4_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_2_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_7_0_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_15_8_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_23_16_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_31_24_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_39_32_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_47_40_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_55_48_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_63_56_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_71_64_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_79_72_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_87_80_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_95_88_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_103_96_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_111_104_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_15_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_sdt_119_112_lpi_1_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_11_data_in_tmp_operator_for_16_data_in_tmp_operator_for_slc_drf_data_in_8_7_0_1_pmx_sva_1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_6_sva_1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_6_sva_1;
  wire [3:0] operator_4_false_acc_psp_6_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_6_sva_1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_7_sva_1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_7_sva_1;
  wire [3:0] operator_4_false_acc_psp_7_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_7_sva_1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_10_sva_1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_10_sva_1;
  wire [3:0] operator_4_false_acc_psp_10_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_10_sva_1;
  wire [3:0] adpfloat_tmp_to_fixed_20U_14U_acc_sdt_11_sva_1;
  wire [4:0] nl_adpfloat_tmp_to_fixed_20U_14U_acc_sdt_11_sva_1;
  wire [3:0] operator_4_false_acc_psp_11_sva_1;
  wire [4:0] nl_operator_4_false_acc_psp_11_sva_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_16;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_18;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_20;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_22;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_24;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_26;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_28;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_10_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_30;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_32;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_34;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_36;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_38;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_40;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_42;
  wire [7:0] crossbar_spec_PE_Weight_WordType_16U_16U_for_6_data_in_tmp_operator_for_15_data_in_tmp_operator_for_data_in_tmp_operator_for_mux_44;
  wire [2:0] PECore_RunBias_if_for_if_bias_tmp2_mux_17;
  wire PECore_PushAxiRsp_if_asn_66;
  wire PECore_PushAxiRsp_if_asn_68;
  wire [3:0] PEManager_16U_GetWeightAddr_if_slc_pe_manager_base_weight_16_15_0_ncse_sva_mx0_3_0;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1_3;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1_2;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1_1;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1_0;
  wire [2:0] crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_15_lpi_1_dfm_1_3_1;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_15_lpi_1_dfm_1_0;
  reg [7:0] reg_Datapath_for_conc_4_ftd;
  reg [7:0] reg_Datapath_for_conc_4_ftd_1;
  reg [7:0] reg_Datapath_for_conc_4_ftd_2;
  reg [7:0] reg_Datapath_for_conc_4_ftd_3;
  reg [7:0] reg_Datapath_for_conc_4_ftd_4;
  reg [7:0] reg_Datapath_for_conc_4_ftd_5;
  reg [7:0] reg_Datapath_for_conc_4_ftd_6;
  reg [7:0] reg_Datapath_for_conc_4_ftd_7;
  reg [7:0] reg_Datapath_for_conc_4_ftd_8;
  reg [7:0] reg_Datapath_for_conc_4_ftd_9;
  reg [7:0] reg_Datapath_for_conc_4_ftd_10;
  reg [7:0] reg_Datapath_for_conc_4_ftd_11;
  reg [7:0] reg_Datapath_for_conc_4_ftd_12;
  reg [7:0] reg_Datapath_for_conc_4_ftd_13;
  reg [7:0] reg_Datapath_for_conc_4_ftd_14;
  reg [7:0] reg_Datapath_for_conc_4_ftd_15;
  reg reg_PECore_RunMac_if_mux_143_ftd;
  reg [6:0] reg_PECore_RunMac_if_mux_143_ftd_1;
  reg [3:0] reg_PECore_RunMac_if_mux_142_ftd;
  reg [3:0] reg_PECore_RunMac_if_mux_142_ftd_1;
  reg [2:0] reg_PECore_RunMac_if_mux_141_ftd;
  reg [4:0] reg_PECore_RunMac_if_mux_141_ftd_1;
  reg [5:0] reg_PECore_RunMac_if_mux_140_ftd;
  reg [1:0] reg_PECore_RunMac_if_mux_140_ftd_1;
  reg [2:0] reg_PECore_RunMac_if_mux_14_ftd;
  reg [4:0] reg_PECore_RunMac_if_mux_14_ftd_1;
  reg [5:0] reg_PECore_RunMac_if_mux_139_ftd;
  reg [1:0] reg_PECore_RunMac_if_mux_139_ftd_1;
  reg [2:0] reg_PECore_RunMac_if_mux_138_ftd;
  reg [4:0] reg_PECore_RunMac_if_mux_138_ftd_1;
  reg [5:0] reg_PECore_RunMac_if_mux_137_ftd;
  reg [1:0] reg_PECore_RunMac_if_mux_137_ftd_1;
  reg [3:0] reg_PECore_RunMac_if_mux_129_ftd;
  reg [3:0] reg_PECore_RunMac_if_mux_129_ftd_1;
  reg [3:0] reg_PECore_RunMac_if_mux_128_ftd;
  reg [3:0] reg_PECore_RunMac_if_mux_128_ftd_1;
  reg [3:0] reg_PECore_RunMac_if_mux_127_ftd;
  reg [3:0] reg_PECore_RunMac_if_mux_127_ftd_1;
  reg [3:0] reg_PECore_RunMac_if_mux_126_ftd;
  reg [3:0] reg_PECore_RunMac_if_mux_126_ftd_1;
  reg [3:0] reg_PECore_RunMac_if_mux_125_ftd;
  reg [3:0] reg_PECore_RunMac_if_mux_125_ftd_1;
  reg [3:0] reg_PECore_RunMac_if_mux_124_ftd;
  reg [3:0] reg_PECore_RunMac_if_mux_124_ftd_1;
  reg [3:0] reg_PECore_RunMac_if_mux_123_ftd;
  reg [3:0] reg_PECore_RunMac_if_mux_123_ftd_1;
  reg [3:0] reg_PECore_RunMac_if_mux_11_ftd;
  reg [3:0] reg_PECore_RunMac_if_mux_11_ftd_1;
  reg [3:0] reg_PECore_RunMac_if_mux_122_ftd;
  reg [3:0] reg_PECore_RunMac_if_mux_122_ftd_1;
  wire PECore_RunBias_if_for_or_m1c_5;
  wire and_4031_m1c;
  wire PECore_RunMac_if_or_5_m1c;
  wire PECore_DecodeAxiRead_switch_lp_and_3_rgt;
  wire operator_32_true_and_6_rgt;
  wire PECore_RunBias_if_for_and_50_rgt;
  wire operator_32_true_and_2_rgt;
  wire PECore_RunMac_if_nand_56_rgt;
  wire PECore_RunMac_if_and_674_rgt;
  wire PECore_RunMac_if_and_675_rgt;
  wire PECore_RunMac_if_and_676_rgt;
  wire PECore_RunMac_if_and_627_rgt;
  wire PECore_RunMac_if_and_628_rgt;
  wire PECore_RunMac_if_and_580_rgt;
  wire PECore_RunMac_if_and_569_rgt;
  wire PECore_RunMac_if_and_570_rgt;
  wire PECore_RunMac_if_and_571_rgt;
  wire PECore_RunBias_if_for_and_45_rgt;
  wire PECore_RunBias_if_for_and_34_rgt;
  wire rva_out_reg_data_and_87_rgt;
  wire rva_out_reg_data_and_88_rgt;
  wire PECore_RunMac_if_and_346_rgt;
  reg reg_PECore_RunMac_asn_15_itm_1_ftd;
  reg reg_PECore_RunMac_asn_15_itm_1_ftd_1;
  reg reg_PECore_RunMac_asn_15_itm_1_ftd_2;
  wire PECore_RunMac_if_and_721_ssc;
  reg [2:0] reg_PECore_RunMac_if_mux_100_ftd;
  reg [4:0] reg_PECore_RunMac_if_mux_100_ftd_1;
  reg [2:0] reg_PECore_RunMac_if_mux_101_ftd;
  reg [4:0] reg_PECore_RunMac_if_mux_101_ftd_1;
  wire PECore_RunMac_if_and_723_ssc;
  reg [2:0] reg_PECore_RunMac_if_mux_102_ftd;
  reg [4:0] reg_PECore_RunMac_if_mux_102_ftd_1;
  reg [2:0] reg_PECore_RunMac_if_mux_103_ftd;
  reg [4:0] reg_PECore_RunMac_if_mux_103_ftd_1;
  reg [2:0] reg_PECore_RunMac_if_mux_104_ftd;
  reg [4:0] reg_PECore_RunMac_if_mux_104_ftd_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_7;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_3;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_1;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_sva_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_1_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_2_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_3_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_4_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_5_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_6_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_7_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_8_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_9_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_10_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_11_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_12_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_13_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_14_ssc;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_14;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_13;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_12;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_11;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_10;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_9;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_8;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_7;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_6;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_5;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_4;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_3;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_1;
  reg nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_0;
  wire weight_mem_read_arbxbar_xbar_for_3_1_operator_31_false_operator_31_false_operator_31_false_or_seb;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_1_lpi_1_dfm_3_0;
  wire weight_mem_read_arbxbar_xbar_for_3_2_operator_31_false_operator_31_false_operator_31_false_or_seb;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_2_lpi_1_dfm_3_0;
  wire weight_mem_read_arbxbar_xbar_for_3_3_operator_31_false_operator_31_false_operator_31_false_or_seb;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_3_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_4_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_5_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_6_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_7_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_8_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_9_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_10_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_11_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_12_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_13_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_14_lpi_1_dfm_3_0;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_15_lpi_1_dfm_3_0;
  wire is_start_and_cse;
  wire [31:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_15_cse;
  wire [31:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_14_cse;
  wire [19:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_25_cse;
  wire [19:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_26_cse;
  wire [19:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_21_cse;
  wire [19:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_22_cse;
  wire pe_config_manager_counter_and_cse;
  wire [31:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_2_cse;
  wire [31:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_3_cse;
  wire [31:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_4_cse;
  wire [31:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_12_cse;
  wire [31:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_1_cse;
  wire [31:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_13_cse;
  wire PECore_RunMac_if_and_572_cse;
  wire PECore_RunMac_if_and_cse;
  wire [31:0] PECore_RunBias_if_accum_vector_out_data_mux_5_cse;
  wire [31:0] PECore_RunBias_if_accum_vector_out_data_mux_9_cse;
  wire [31:0] PECore_RunBias_if_accum_vector_out_data_mux_11_cse;
  wire [31:0] PECore_RunBias_if_accum_vector_out_data_mux_7_cse;
  wire PECore_RunMac_if_and_434_cse;
  wire PECore_RunMac_if_and_433_cse;
  wire and_5541_cse;
  wire or_796_cse;
  wire or_3399_cse;
  wire PECore_RunMac_if_and_470_cse;
  wire PECore_RunMac_if_and_444_cse;
  wire PECore_RunMac_if_and_445_cse;
  wire PECore_RunMac_if_and_398_cse;
  wire PECore_RunMac_if_and_399_cse;
  wire PECore_RunMac_if_and_390_cse;
  wire PECore_RunMac_if_and_391_cse;
  wire while_and_74_cse;
  wire while_and_66_cse;
  reg [2:0] reg_PECore_RunMac_if_mux_10_ftd;
  reg [4:0] reg_PECore_RunMac_if_mux_10_ftd_1;
  reg [2:0] reg_PECore_RunMac_if_mux_1_ftd;
  reg [4:0] reg_PECore_RunMac_if_mux_1_ftd_1;
  wire PECore_RunMac_if_or_140_m1c;
  wire PECore_RunMac_if_or_143_m1c;
  wire PECore_RunMac_if_or_145_m1c;
  wire PECore_RunBias_if_accum_vector_out_data_and_15_rgt;
  wire PECore_RunMac_if_and_817_rgt;
  wire PECore_RunMac_if_and_472_rgt;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_1_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_2_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_3_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_4_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_5_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_6_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_7_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_8_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_9_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_10_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_11_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_12_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_13_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_14_lpi_1_dfm_1_mx1_2;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_15_lpi_1_dfm_1_mx1_2;
  wire accum_vector_data_and_6_cse;
  wire act_port_reg_data_and_8_cse;
  wire weight_port_read_out_data_and_cse;
  wire weight_port_read_out_data_and_16_cse;
  wire weight_port_read_out_data_and_32_cse;
  wire weight_port_read_out_data_and_48_cse;
  wire weight_port_read_out_data_and_64_cse;
  wire weight_port_read_out_data_and_80_cse;
  wire weight_port_read_out_data_and_96_cse;
  wire weight_port_read_out_data_and_112_cse;
  wire weight_port_read_out_data_and_128_cse;
  wire weight_port_read_out_data_and_136_cse;
  wire weight_port_read_out_data_and_152_cse;
  wire weight_port_read_out_data_and_168_cse;
  wire weight_port_read_out_data_and_184_cse;
  wire weight_port_read_out_data_and_200_cse;
  wire accum_vector_data_and_9_cse;
  wire PECore_DecodeAxi_if_and_3_cse;
  wire or_1534_cse;
  wire PECore_CheckStart_start_reg_and_cse;
  wire operator_4_false_and_cse;
  wire adpfloat_tmp_is_zero_aelse_and_cse;
  wire operator_32_true_and_12_cse;
  wire weight_port_read_out_data_and_216_cse;
  wire weight_port_read_out_data_and_232_cse;
  wire adpfloat_tmp_is_zero_aelse_and_4_cse;
  wire accum_vector_data_and_15_cse;
  wire adpfloat_tmp_is_zero_aelse_and_6_cse;
  wire PECore_RunMac_if_and_685_cse;
  wire PECore_RunMac_if_and_701_cse;
  wire PECore_RunMac_if_and_717_cse;
  wire PECore_RunMac_if_and_726_cse;
  wire while_and_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_2_cse;
  wire PECore_RunBias_if_for_and_47_cse;
  wire PECore_RunBias_if_for_and_48_cse;
  wire and_2966_cse;
  wire act_port_reg_data_and_24_cse;
  wire rva_out_reg_data_and_91_cse;
  wire pe_config_UpdateInputCounter_if_and_cse;
  wire PECore_RunBias_if_for_and_42_cse;
  wire or_1521_cse;
  wire PECore_RunBias_if_for_and_cse;
  wire PECore_RunMac_if_and_359_cse;
  wire PECore_RunMac_if_and_360_cse;
  wire PECore_RunMac_if_and_361_cse;
  wire PECore_RunMac_if_and_834_rgt;
  wire PECore_RunMac_if_and_820_rgt;
  wire PECore_RunMac_if_and_430_cse;
  wire PECore_RunMac_if_and_431_cse;
  wire PECore_RunBias_if_accum_vector_out_data_and_17_cse;
  wire PECore_RunMac_if_and_859_cse;
  wire PECore_RunMac_if_and_867_cse;
  wire PECore_RunMac_if_and_872_cse;
  wire pe_config_UpdateManagerCounter_if_unequal_tmp;
  wire and_5872_cse;
  wire and_5844_cse;
  wire and_5871_cse;
  reg reg_PECore_RunMac_if_mux_123_1_enexo;
  reg reg_PECore_RunMac_if_mux_142_1_enexo;
  reg reg_rva_out_reg_data_47_40_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_63_56_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_71_64_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_79_72_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_87_80_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_95_88_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_103_96_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_111_104_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_119_112_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_127_120_sva_dfm_4_enexo;
  reg reg_act_port_reg_data_0_enexo;
  reg reg_act_port_reg_data_1_enexo;
  reg reg_act_port_reg_data_2_enexo;
  reg reg_act_port_reg_data_3_enexo;
  reg reg_act_port_reg_data_4_enexo;
  reg reg_act_port_reg_data_5_enexo;
  reg reg_act_port_reg_data_6_enexo;
  reg reg_act_port_reg_data_9_enexo;
  reg reg_act_port_reg_data_10_enexo;
  reg reg_act_port_reg_data_asn_3_enexo;
  reg reg_act_port_reg_data_asn_2_enexo;
  reg reg_act_port_reg_data_asn_1_enexo;
  reg reg_act_port_reg_data_asn_enexo;
  reg reg_act_port_reg_data_14_enexo;
  reg reg_act_port_reg_data_13_enexo;
  reg reg_act_port_reg_data_12_enexo;
  reg reg_act_port_reg_data_15_enexo;
  reg reg_PECore_RunMac_if_mux_31_enexo;
  wire PECore_PushAxiRsp_if_and_47_enex5;
  wire PECore_PushAxiRsp_if_and_48_enex5;
  wire PECore_PushAxiRsp_if_and_49_enex5;
  wire PECore_PushAxiRsp_if_and_50_enex5;
  wire PECore_PushAxiRsp_if_and_51_enex5;
  wire PECore_PushAxiRsp_if_and_52_enex5;
  wire PECore_PushAxiRsp_if_and_53_enex5;
  wire PECore_PushAxiRsp_if_and_54_enex5;
  wire PECore_PushAxiRsp_if_and_55_enex5;
  wire PECore_PushAxiRsp_if_and_56_enex5;
  wire PECore_PushAxiRsp_if_and_57_enex5;
  wire PECore_PushAxiRsp_if_and_58_enex5;
  wire PECore_PushAxiRsp_if_and_59_enex5;
  wire PECore_PushOutput_if_and_16_enex5;
  wire PECore_PushOutput_if_and_17_enex5;
  wire PECore_PushOutput_if_and_18_enex5;
  wire PECore_PushOutput_if_and_19_enex5;
  wire PECore_PushOutput_if_and_20_enex5;
  wire PECore_PushOutput_if_and_21_enex5;
  wire PECore_PushOutput_if_and_22_enex5;
  wire PECore_PushOutput_if_and_25_enex5;
  wire PECore_PushOutput_if_and_26_enex5;
  wire PECore_PushOutput_if_and_28_enex5;
  wire PECore_PushOutput_if_and_29_enex5;
  wire PECore_PushOutput_if_and_30_enex5;
  wire PECore_PushOutput_if_and_31_enex5;
  wire act_port_reg_data_and_enex5;
  wire act_port_reg_data_and_28_enex5;
  wire act_port_reg_data_and_29_enex5;
  wire act_port_reg_data_and_30_enex5;
  wire Datapath_for_and_enex5;
  wire PECore_RunMac_if_and_854_tmp;
  wire PECore_RunMac_if_and_865_tmp;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_and_15_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_16_operator_31_false_operator_31_false_operator_31_false_or_cse;
  wire PECore_RunMac_if_and_860_cse;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_1_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_2_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_3_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_4_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_5_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_6_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_7_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_8_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_9_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_10_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_11_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_12_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_13_itm;
  wire weight_mem_read_arbxbar_xbar_for_3_16_Arbiter_16U_Roundrobin_pick_if_1_temp2_or_14_itm;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_1;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_2;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_3;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_4;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_5;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_6;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_7;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_8;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_9;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_10;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_11;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_12;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_13;
  reg reg_nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_ftd_14;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_14;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_13;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_12;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_11;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_10;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_9;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_8;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_7;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_6;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_5;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_4;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_3;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_2;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_1;
  wire Arbiter_16U_Roundrobin_pick_mux_2460_tmp_0;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_14;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_13;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_12;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_11;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_10;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_9;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_8;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_6;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_5;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_4;
  wire nvhls_set_slc_Arbiter_16U_Roundrobin_Mask_nvhls_nvhls_t_15U_nvuint_t_X_temp_15_1_lpi_1_dfm_1_mx1_2;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_14;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_13;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_12;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_11;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_10;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_9;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_8;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_7;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_6;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_5;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_4;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_3;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_2;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_1;
  wire Arbiter_16U_Roundrobin_pick_return_15_1_lpi_1_dfm_3_0;
  wire [11:0] operator_16_false_1_mux_10_cse;
  wire operator_16_false_1_mux_14_cse;
  wire z_out_10_13;
  wire z_out_11_13;
  wire z_out_12_13;
  wire z_out_13_13;
  wire z_out_21_32;
  wire z_out_22_32;
  wire z_out_23_32;
  wire z_out_24_32;
  wire [15:0] operator_16_false_1_mux_16_cse;
  wire while_mux_440_cse;
  wire adpfloat_tmp_to_fixed_20U_14U_mux1h_28_tmp;
  wire or_3880_tmp;
  wire while_while_mux_15_m1c;
  wire while_mux1h_62_m1c;
  wire while_while_mux_13_m1c;
  wire while_mux1h_57_m1c;
  wire while_while_mux_11_m1c;
  wire while_mux1h_52_m1c;
  wire while_while_mux_9_m1c;
  wire while_mux1h_47_m1c;
  wire PEManager_16U_GetInputAddr_1_PEManager_16U_GetInputAddr_1_mux_5_tmp;
  wire adpfloat_tmp_to_fixed_20U_14U_mux1h_29_tmp;
  wire adpfloat_tmp_to_fixed_20U_14U_mux1h_30_tmp;
  wire adpfloat_tmp_to_fixed_20U_14U_mux1h_32_tmp;
  wire while_while_nor_cse;
  wire while_and_268_cse;

  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_10;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_10;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_11;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_12;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_12;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_13;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_28;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_28;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_28;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_28;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_14;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_14;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_29;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_29;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_29;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_29;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_30;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_30;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_30;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_30;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_15;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_31;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_31;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_31;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_31;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_32;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_32;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_32;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_32;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_16;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_16;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_33;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_33;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_33;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_33;
  wire PECore_PushAxiRsp_if_else_mux_14_nl;
  wire PECore_DecodeAxi_mux_139_nl;
  wire PECore_DecodeAxi_if_mux_74_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_19_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_11_nl;
  wire[6:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_18_nl;
  wire PECore_PushAxiRsp_if_else_mux_15_nl;
  wire PECore_DecodeAxi_mux_141_nl;
  wire PECore_DecodeAxi_if_mux_126_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_17_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_8_nl;
  wire[1:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl;
  wire[4:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_15_nl;
  wire PECore_PushAxiRsp_if_else_mux_16_nl;
  wire PECore_DecodeAxi_mux_143_nl;
  wire PECore_DecodeAxi_if_mux_127_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_13_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_5_nl;
  wire[1:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_12_nl;
  wire[4:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_10_nl;
  wire PECore_PushAxiRsp_if_else_mux_17_nl;
  wire PECore_DecodeAxi_mux_145_nl;
  wire PECore_DecodeAxi_if_mux_128_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_12_nl;
  wire[1:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_9_nl;
  wire[4:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl;
  wire input_mem_banks_read_read_data_and_nl;
  wire mux_594_nl;
  wire or_1536_nl;
  wire mux_593_nl;
  wire mux_592_nl;
  wire mux_591_nl;
  wire nor_244_nl;
  wire or_1531_nl;
  wire or_1530_nl;
  wire mux_596_nl;
  wire mux_595_nl;
  wire nor_242_nl;
  wire nor_243_nl;
  wire mux_600_nl;
  wire mux_599_nl;
  wire mux_598_nl;
  wire nor_241_nl;
  wire mux_597_nl;
  wire PECore_UpdateFSM_switch_lp_mux_6_nl;
  wire PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_7_nl;
  wire and_3383_nl;
  wire PECore_UpdateFSM_switch_lp_mux1h_42_nl;
  wire PECore_UpdateFSM_switch_lp_not_47_nl;
  wire PECore_UpdateFSM_switch_lp_not_48_nl;
  wire PECore_UpdateFSM_switch_lp_not_49_nl;
  wire while_and_221_nl;
  wire while_and_225_nl;
  wire while_and_226_nl;
  wire while_and_227_nl;
  wire[19:0] mux1h_12_nl;
  wire while_or_11_nl;
  wire while_and_288_nl;
  wire while_and_289_nl;
  wire while_mux1h_46_nl;
  wire while_and_222_nl;
  wire while_and_223_nl;
  wire while_and_224_nl;
  wire while_and_290_nl;
  wire while_mux1h_48_nl;
  wire PECore_RunBias_if_for_and_55_nl;
  wire PECore_RunBias_if_for_and_56_nl;
  wire PECore_RunBias_if_for_and_57_nl;
  wire while_mux1h_49_nl;
  wire while_and_228_nl;
  wire while_and_229_nl;
  wire while_and_230_nl;
  wire PECore_UpdateFSM_switch_lp_not_65_nl;
  wire while_and_231_nl;
  wire while_and_235_nl;
  wire while_and_236_nl;
  wire while_and_237_nl;
  wire[19:0] mux1h_13_nl;
  wire while_or_10_nl;
  wire while_and_283_nl;
  wire while_and_284_nl;
  wire while_mux1h_51_nl;
  wire while_and_232_nl;
  wire while_and_233_nl;
  wire while_and_234_nl;
  wire while_and_285_nl;
  wire while_mux1h_53_nl;
  wire PECore_RunBias_if_for_and_58_nl;
  wire PECore_RunBias_if_for_and_59_nl;
  wire PECore_RunBias_if_for_and_60_nl;
  wire while_mux1h_54_nl;
  wire while_and_238_nl;
  wire while_and_239_nl;
  wire while_and_240_nl;
  wire PECore_UpdateFSM_switch_lp_not_66_nl;
  wire while_and_241_nl;
  wire while_and_245_nl;
  wire while_and_246_nl;
  wire while_and_247_nl;
  wire[19:0] mux1h_14_nl;
  wire while_or_9_nl;
  wire while_and_278_nl;
  wire while_and_279_nl;
  wire while_mux1h_56_nl;
  wire while_and_242_nl;
  wire while_and_243_nl;
  wire while_and_244_nl;
  wire while_and_280_nl;
  wire while_mux1h_58_nl;
  wire PECore_RunBias_if_for_and_61_nl;
  wire PECore_RunBias_if_for_and_62_nl;
  wire PECore_RunBias_if_for_and_63_nl;
  wire while_mux1h_59_nl;
  wire while_and_248_nl;
  wire PECore_UpdateFSM_switch_lp_not_67_nl;
  wire while_and_249_nl;
  wire while_and_253_nl;
  wire while_and_254_nl;
  wire while_and_255_nl;
  wire[19:0] mux1h_15_nl;
  wire while_or_nl;
  wire while_and_273_nl;
  wire while_and_274_nl;
  wire while_mux1h_61_nl;
  wire while_and_250_nl;
  wire while_and_251_nl;
  wire while_and_252_nl;
  wire while_and_275_nl;
  wire while_mux1h_63_nl;
  wire PECore_RunBias_if_for_and_64_nl;
  wire PECore_RunBias_if_for_and_65_nl;
  wire PECore_RunBias_if_for_and_66_nl;
  wire while_mux1h_64_nl;
  wire while_and_256_nl;
  wire PECore_UpdateFSM_switch_lp_not_38_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_if_1_crossbar_spec_PE_Weight_WordType_16U_16U_for_if_1_crossbar_spec_PE_Weight_WordType_16U_16U_for_if_1_nor_5_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_252_nl;
  wire[3:0] pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_and_1_nl;
  wire pe_config_UpdateManagerCounter_if_not_7_nl;
  wire and_3501_nl;
  wire[31:0] while_mux1h_67_nl;
  wire while_and_269_nl;
  wire while_and_270_nl;
  wire PECore_UpdateFSM_switch_lp_not_55_nl;
  wire[31:0] while_mux_nl;
  wire PECore_UpdateFSM_switch_lp_not_56_nl;
  wire[31:0] while_mux1h_65_nl;
  wire PECore_UpdateFSM_switch_lp_not_57_nl;
  wire[31:0] while_mux_449_nl;
  wire PECore_UpdateFSM_switch_lp_not_58_nl;
  wire[19:0] while_while_mux1h_12_nl;
  wire while_and_202_nl;
  wire while_and_203_nl;
  wire while_and_204_nl;
  wire PECore_RunBias_if_for_and_25_nl;
  wire while_and_82_nl;
  wire PECore_UpdateFSM_switch_lp_not_36_nl;
  wire[19:0] while_while_mux1h_13_nl;
  wire while_and_199_nl;
  wire while_and_200_nl;
  wire while_and_201_nl;
  wire PECore_RunBias_if_for_and_27_nl;
  wire while_and_84_nl;
  wire PECore_UpdateFSM_switch_lp_not_64_nl;
  wire[19:0] while_while_mux1h_14_nl;
  wire while_and_196_nl;
  wire while_and_197_nl;
  wire while_and_198_nl;
  wire PECore_RunBias_if_for_and_29_nl;
  wire while_and_86_nl;
  wire PECore_UpdateFSM_switch_lp_not_63_nl;
  wire[19:0] while_while_mux1h_15_nl;
  wire while_and_193_nl;
  wire while_and_194_nl;
  wire while_and_195_nl;
  wire PECore_RunBias_if_for_and_31_nl;
  wire while_and_88_nl;
  wire PECore_UpdateFSM_switch_lp_not_62_nl;
  wire PECore_UpdateFSM_switch_lp_mux_7_nl;
  wire pe_config_UpdateManagerCounter_mux_1_nl;
  wire pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl;
  wire and_3991_nl;
  wire[7:0] pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl;
  wire pe_config_UpdateInputCounter_if_not_2_nl;
  wire PECore_UpdateFSM_switch_lp_and_nl;
  wire[7:0] pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl;
  wire pe_config_UpdateManagerCounter_if_not_9_nl;
  wire and_4037_nl;
  wire PECore_UpdateFSM_switch_lp_not_50_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_94_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_92_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_90_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_88_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_86_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_84_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_82_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_80_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_81_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_83_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_85_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_87_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_89_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_91_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_93_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_95_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_78_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_76_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_74_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_72_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_70_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_68_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_66_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_64_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_65_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_67_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_69_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_71_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_73_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_75_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_77_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_79_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_62_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_60_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_58_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_56_nl;
  wire[2:0] PEManager_16U_ClusterLookup_for_mux_54_nl;
  wire[4:0] PECore_RunBias_if_for_10_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_10_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_10_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_10_operator_33_true_acc_nl;
  wire[4:0] PEManager_16U_ClusterLookup_for_mux_139_nl;
  wire[2:0] PEManager_16U_ClusterLookup_for_mux_52_nl;
  wire[4:0] PECore_RunBias_if_for_11_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_11_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_11_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_11_operator_33_true_acc_nl;
  wire[4:0] PEManager_16U_ClusterLookup_for_mux_140_nl;
  wire[2:0] PEManager_16U_ClusterLookup_for_mux_50_nl;
  wire[4:0] PEManager_16U_ClusterLookup_for_mux_141_nl;
  wire[4:0] PECore_RunBias_if_for_5_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_5_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_5_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_5_operator_33_true_acc_nl;
  wire PECore_RunMac_if_and_829_nl;
  wire[2:0] PEManager_16U_ClusterLookup_for_mux_48_nl;
  wire[4:0] PECore_RunBias_if_for_6_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_6_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_6_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_6_operator_33_true_acc_nl;
  wire[4:0] PEManager_16U_ClusterLookup_for_mux_142_nl;
  wire[2:0] PEManager_16U_ClusterLookup_for_mux_49_nl;
  wire[4:0] PECore_RunBias_if_for_7_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_7_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_7_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_7_operator_33_true_acc_nl;
  wire[4:0] PEManager_16U_ClusterLookup_for_mux_143_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_51_nl;
  wire[4:0] PECore_RunBias_if_for_8_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_8_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_8_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_8_operator_33_true_acc_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_53_nl;
  wire[4:0] PECore_RunBias_if_for_9_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_9_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_9_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_9_operator_33_true_acc_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_55_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_57_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_59_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_61_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_63_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_46_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_44_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_42_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_40_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_38_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_36_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_34_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_32_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_33_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_35_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_37_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_39_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_41_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_43_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_45_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_47_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_2_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux1h_6_nl;
  wire PECore_RunBias_if_for_and_49_nl;
  wire PECore_RunBias_if_for_and_40_nl;
  wire PECore_RunBias_if_for_and_36_nl;
  wire PECore_DecodeAxi_mux_133_nl;
  wire PECore_DecodeAxi_if_mux_67_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_or_1_nl;
  wire adpfloat_tmp_is_zero_if_adpfloat_tmp_is_zero_if_nor_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_29_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_7_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_62_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_28_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_8_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_60_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_27_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_9_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_58_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_26_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_10_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_56_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_25_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_19_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_49_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_18_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_51_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_20_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_48_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_21_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_4_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_22_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_52_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_20_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_23_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_50_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_and_3_nl;
  wire[7:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_9_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_11_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_54_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux1h_13_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux1h_11_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux1h_16_nl;
  wire PECore_DecodeAxi_mux_138_nl;
  wire PECore_DecodeAxi_if_mux_125_nl;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_or_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_258_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_257_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_256_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_255_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_254_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_251_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_250_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_249_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_248_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_247_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_246_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_245_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_244_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_for_mux_253_nl;
  wire PECore_RunMac_nor_nl;
  wire PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl;
  wire PECore_UpdateFSM_case_1_if_mux_nl;
  wire pe_manager_zero_active_mux_nl;
  wire PECore_DecodeAxi_mux_127_nl;
  wire PECore_DecodeAxi_if_mux_57_nl;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_34_nl;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_32_nl;
  wire pe_manager_zero_active_mux_1_nl;
  wire PECore_DecodeAxi_mux_125_nl;
  wire PECore_DecodeAxi_if_mux_55_nl;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_35_nl;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_33_nl;
  wire[2:0] PEManager_16U_ClusterLookup_for_mux_15_nl;
  wire[4:0] PEManager_16U_ClusterLookup_for_mux_145_nl;
  wire[4:0] PECore_RunBias_if_for_3_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_3_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_3_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_3_operator_33_true_acc_nl;
  wire[2:0] PEManager_16U_ClusterLookup_for_mux_6_nl;
  wire[4:0] PEManager_16U_ClusterLookup_for_mux_144_nl;
  wire[4:0] PECore_RunBias_if_for_4_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_4_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_4_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_4_operator_33_true_acc_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_3_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_74_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_72_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_70_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_68_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_66_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_64_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_65_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_30_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_94_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_31_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_92_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_32_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_90_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_33_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_88_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_34_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_86_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_35_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_84_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_36_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_82_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_37_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_80_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_38_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_81_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_39_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_83_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_40_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_85_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_41_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_87_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_42_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_89_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_43_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_91_nl;
  wire[7:0] weight_mem_run_1_for_5_mux_44_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_93_nl;
  wire[7:0] data_in_tmp_operator_for_mux_34_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_95_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_46_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_44_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_42_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_40_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_38_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_36_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_34_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_32_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_33_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_35_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_37_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_39_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_41_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_43_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_45_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_47_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_30_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_28_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_26_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_24_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_22_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_20_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_18_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_16_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_17_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_19_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_21_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_23_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_25_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_27_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_29_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_31_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_30_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_28_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_26_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_24_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_22_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_20_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_18_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_16_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_17_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_19_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_21_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_23_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_25_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_27_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_29_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_31_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_1_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_2_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_3_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_4_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_5_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_6_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_7_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_8_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_9_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_10_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_11_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_12_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_13_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_14_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_15_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_14_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_13_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_12_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_11_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_10_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_9_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_8_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_7_nl;
  wire[7:0] PEManager_16U_ClusterLookup_for_mux_1_nl;
  wire mux_22_nl;
  wire nand_198_nl;
  wire nor_475_nl;
  wire pe_config_is_cluster_not_39_nl;
  wire[11:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_40_nl;
  wire[11:0] PECore_RunFSM_switch_lp_mux_28_nl;
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_43_nl;
  wire PECore_RunFSM_switch_lp_mux_29_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3212_nl;
  wire weight_mem_run_1_if_for_if_and_702_nl;
  wire PECore_DecodeAxi_mux_134_nl;
  wire PECore_DecodeAxi_if_mux_122_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_mux_5_nl;
  wire PECore_DecodeAxi_mux_135_nl;
  wire PECore_DecodeAxi_if_mux_123_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_or_nl;
  wire PECore_RunFSM_case_0_if_mux_1_nl;
  wire or_1624_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_465_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_466_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_468_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_469_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_470_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_471_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_472_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_473_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_474_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_475_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_476_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_477_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_478_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_479_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_1_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_2995_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_2994_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_2992_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_2988_nl;
  wire[15:0] operator_16_false_1_acc_12_nl;
  wire[16:0] nl_operator_16_false_1_acc_12_nl;
  wire[14:0] operator_16_false_1_acc_nl;
  wire[15:0] nl_operator_16_false_1_acc_nl;
  wire[15:0] operator_16_false_1_acc_11_nl;
  wire[16:0] nl_operator_16_false_1_acc_11_nl;
  wire[13:0] operator_16_false_1_acc_8_nl;
  wire[14:0] nl_operator_16_false_1_acc_8_nl;
  wire[13:0] operator_16_false_1_mux_20_nl;
  wire[15:0] operator_16_false_1_acc_10_nl;
  wire[16:0] nl_operator_16_false_1_acc_10_nl;
  wire[14:0] operator_16_false_1_acc_7_nl;
  wire[15:0] nl_operator_16_false_1_acc_7_nl;
  wire[15:0] operator_16_false_1_acc_9_nl;
  wire[16:0] nl_operator_16_false_1_acc_9_nl;
  wire[12:0] operator_16_false_1_acc_3_nl;
  wire[13:0] nl_operator_16_false_1_acc_3_nl;
  wire[15:0] PECore_RunFSM_case_2_else_for_10_operator_16_false_1_acc_nl;
  wire[16:0] nl_PECore_RunFSM_case_2_else_for_10_operator_16_false_1_acc_nl;
  wire[14:0] operator_16_false_1_acc_4_nl;
  wire[15:0] nl_operator_16_false_1_acc_4_nl;
  wire[15:0] PECore_RunFSM_case_2_else_for_12_operator_16_false_1_acc_nl;
  wire[16:0] nl_PECore_RunFSM_case_2_else_for_12_operator_16_false_1_acc_nl;
  wire[13:0] operator_16_false_1_acc_5_nl;
  wire[14:0] nl_operator_16_false_1_acc_5_nl;
  wire[15:0] PECore_RunFSM_case_2_else_for_14_operator_16_false_1_acc_nl;
  wire[16:0] nl_PECore_RunFSM_case_2_else_for_14_operator_16_false_1_acc_nl;
  wire[14:0] operator_16_false_1_acc_6_nl;
  wire[15:0] nl_operator_16_false_1_acc_6_nl;
  wire[15:0] PECore_RunFSM_case_2_else_for_16_operator_16_false_1_acc_nl;
  wire[16:0] nl_PECore_RunFSM_case_2_else_for_16_operator_16_false_1_acc_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_1_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_435_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_436_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_438_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_439_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_440_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_441_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_442_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_443_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_444_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_445_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_446_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_447_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_448_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_449_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_2_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3009_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3008_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3006_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3002_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_2_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_405_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_406_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_408_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_409_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_410_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_411_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_412_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_413_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_414_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_415_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_416_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_417_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_418_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_419_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_3_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3023_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3022_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3020_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3016_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_3_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_375_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_376_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_378_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_379_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_380_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_381_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_382_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_383_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_384_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_385_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_386_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_387_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_388_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_389_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_4_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3037_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3036_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3034_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3030_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_4_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_345_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_346_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_348_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_349_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_350_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_351_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_352_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_353_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_354_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_355_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_356_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_357_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_358_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_359_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_5_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3051_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3050_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3048_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3044_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_5_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_315_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_316_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_318_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_319_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_320_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_321_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_322_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_323_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_324_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_325_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_326_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_327_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_328_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_329_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_6_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3065_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3064_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3062_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3058_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_6_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_285_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_286_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_288_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_289_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_290_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_291_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_292_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_293_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_294_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_295_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_296_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_297_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_298_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_299_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_7_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3079_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3078_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3076_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3072_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_7_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_255_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_256_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_258_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_259_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_260_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_261_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_262_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_263_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_264_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_265_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_266_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_267_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_268_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_269_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_8_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3093_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3092_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3090_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3086_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_8_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_225_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_226_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_228_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_229_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_230_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_231_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_232_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_233_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_234_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_235_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_236_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_237_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_238_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_239_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_9_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3107_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3106_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3104_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3100_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_9_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_195_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_196_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_198_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_199_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_200_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_201_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_202_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_203_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_204_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_205_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_206_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_207_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_208_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_209_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_10_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3121_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3120_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3118_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3114_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_10_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_165_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_166_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_168_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_169_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_170_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_171_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_172_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_173_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_174_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_175_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_176_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_177_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_178_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_179_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_11_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3135_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3134_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3132_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3128_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_11_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_135_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_136_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_138_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_139_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_140_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_141_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_142_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_143_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_144_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_145_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_146_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_147_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_148_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_149_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_12_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3149_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3148_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3146_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3142_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_12_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_105_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_106_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_108_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_109_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_110_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_111_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_112_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_113_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_114_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_115_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_116_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_117_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_118_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_119_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_13_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3163_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3162_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3160_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3156_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_13_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_75_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_76_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_78_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_79_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_80_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_81_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_82_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_83_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_84_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_85_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_86_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_87_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_88_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_89_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_14_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3177_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3176_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3174_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3170_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_14_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_45_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_46_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_48_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_49_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_50_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_51_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_52_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_53_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_54_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_55_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_56_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_57_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_58_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_59_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_15_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3191_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3190_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3188_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3184_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_15_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_15_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_16_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_18_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_19_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_20_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_21_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_22_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_23_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_24_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_25_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_26_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_27_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_28_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_and_29_nl;
  wire weight_mem_read_arbxbar_xbar_for_3_16_operator_8_false_operator_8_false_operator_8_false_or_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3216_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3218_nl;
  wire Arbiter_16U_Roundrobin_pick_mux_3219_nl;
  wire weight_mem_run_1_if_for_if_and_697_nl;
  wire weight_mem_run_1_if_for_if_and_693_nl;
  wire weight_mem_run_1_if_for_if_and_689_nl;
  wire weight_mem_run_1_if_for_if_and_690_nl;
  wire weight_mem_run_1_if_for_if_and_694_nl;
  wire weight_mem_run_1_if_for_if_and_698_nl;
  wire weight_mem_run_1_if_for_if_and_703_nl;
  wire weight_mem_run_1_if_for_if_and_701_nl;
  wire weight_mem_run_1_if_for_if_and_699_nl;
  wire weight_mem_run_1_if_for_if_and_695_nl;
  wire weight_mem_run_1_if_for_if_and_688_nl;
  wire weight_mem_run_1_if_for_if_and_692_nl;
  wire weight_mem_run_1_if_for_if_and_696_nl;
  wire weight_mem_run_1_if_for_if_and_700_nl;
  wire PECore_DecodeAxi_mux_149_nl;
  wire PECore_DecodeAxi_if_mux_135_nl;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_56_nl;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_54_nl;
  wire[7:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_mux1h_nl;
  wire PECore_UpdateFSM_switch_lp_or_nl;
  wire PECore_UpdateFSM_switch_lp_and_2_nl;
  wire PECore_UpdateFSM_switch_lp_and_3_nl;
  wire[7:0] PECore_DecodeAxi_if_mux_68_nl;
  wire[3:0] PECore_DecodeAxi_if_mux_69_nl;
  wire weight_mem_run_1_if_for_if_and_691_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_260_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_262_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_264_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_266_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_268_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_270_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_272_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_274_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_276_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_278_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_280_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_282_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_284_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_286_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_256_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_258_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_332_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_347_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_362_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_377_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_392_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_407_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_422_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_437_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_452_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_467_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_482_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_497_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_512_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_527_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_302_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_317_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_331_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_346_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_361_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_376_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_391_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_406_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_421_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_436_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_451_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_466_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_481_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_496_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_511_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_526_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_301_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_316_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_330_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_345_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_360_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_375_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_390_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_405_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_420_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_435_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_450_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_465_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_480_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_495_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_510_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_525_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_300_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_315_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_329_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_344_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_359_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_374_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_389_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_404_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_419_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_434_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_449_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_464_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_479_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_494_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_509_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_524_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_299_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_314_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_328_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_343_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_358_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_373_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_388_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_403_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_418_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_433_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_448_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_463_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_478_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_493_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_508_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_523_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_298_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_313_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_327_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_342_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_357_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_372_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_387_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_402_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_417_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_432_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_447_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_462_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_477_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_492_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_507_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_522_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_297_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_312_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_326_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_341_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_356_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_371_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_386_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_401_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_416_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_431_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_446_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_461_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_476_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_491_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_506_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_521_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_296_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_311_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_325_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_340_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_355_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_370_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_385_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_400_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_415_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_430_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_445_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_460_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_475_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_490_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_505_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_520_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_295_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_310_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_324_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_339_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_354_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_369_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_384_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_399_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_414_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_429_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_444_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_459_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_474_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_489_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_504_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_519_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_294_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_309_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_323_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_338_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_353_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_368_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_383_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_398_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_413_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_428_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_443_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_458_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_473_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_488_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_503_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_518_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_293_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_308_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_322_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_337_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_352_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_367_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_382_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_397_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_412_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_427_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_442_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_457_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_472_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_487_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_502_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_517_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_292_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_307_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_321_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_336_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_351_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_366_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_381_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_396_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_411_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_426_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_441_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_456_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_471_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_486_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_501_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_516_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_291_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_306_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_320_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_335_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_350_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_365_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_380_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_395_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_410_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_425_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_440_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_455_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_470_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_485_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_500_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_515_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_290_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_305_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_319_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_334_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_349_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_364_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_379_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_394_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_409_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_424_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_439_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_454_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_469_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_484_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_499_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_514_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_289_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_304_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_318_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_333_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_348_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_363_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_378_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_393_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_408_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_423_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_438_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_453_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_468_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_483_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_498_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_513_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_288_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_303_nl;
  wire[7:0] while_mux_111_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_36_nl;
  wire[7:0] while_mux_110_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_35_nl;
  wire[7:0] while_mux_109_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_34_nl;
  wire[7:0] while_mux_108_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_33_nl;
  wire[7:0] while_mux_107_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_32_nl;
  wire[7:0] while_mux_106_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_31_nl;
  wire[7:0] while_mux_105_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_30_nl;
  wire[7:0] while_mux_104_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_29_nl;
  wire[7:0] while_mux_103_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_28_nl;
  wire[7:0] while_mux_102_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_27_nl;
  wire[7:0] while_mux_101_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_26_nl;
  wire[7:0] while_mux_100_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_25_nl;
  wire[7:0] while_mux_99_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_24_nl;
  wire[7:0] while_mux_98_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_23_nl;
  wire[7:0] while_mux_97_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_22_nl;
  wire[7:0] while_mux_96_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_21_nl;
  wire[7:0] mux1h_7_nl;
  wire[7:0] PEManager_16U_GetInputAddr_1_acc_nl;
  wire[8:0] nl_PEManager_16U_GetInputAddr_1_acc_nl;
  wire[7:0] PEManager_16U_GetBiasAddr_acc_nl;
  wire[8:0] nl_PEManager_16U_GetBiasAddr_acc_nl;
  wire PECore_DecodeAxi_if_and_nl;
  wire PECore_DecodeAxi_if_and_1_nl;
  wire not_3760_nl;
  wire[7:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_35_nl;
  wire[7:0] PEManager_16U_GetInputAddr_acc_nl;
  wire[8:0] nl_PEManager_16U_GetInputAddr_acc_nl;
  wire or_1589_nl;
  wire mux_601_nl;
  wire and_1488_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_53_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_133_nl;
  wire[3:0] PEManager_16U_ClusterLookup_for_mux_5_nl;
  wire[3:0] PEManager_16U_ClusterLookup_for_mux_138_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_55_nl;
  wire[3:0] PECore_DecodeAxiRead_case_4_switch_lp_and_1_nl;
  wire[3:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_5_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_132_nl;
  wire and_5134_nl;
  wire and_5136_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_and_1_nl;
  wire crossbar_spec_PE_Weight_WordType_16U_16U_source_tmp_and_2_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_57_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_131_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_59_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_130_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_61_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_129_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_63_nl;
  wire[3:0] PEManager_16U_ClusterLookup_1_for_mux_128_nl;
  wire[3:0] PEManager_16U_ClusterLookup_for_mux_78_nl;
  wire[3:0] PEManager_16U_ClusterLookup_for_mux_137_nl;
  wire[3:0] PEManager_16U_ClusterLookup_for_mux_76_nl;
  wire[3:0] PEManager_16U_ClusterLookup_for_mux_136_nl;
  wire[5:0] PEManager_16U_ClusterLookup_for_mux_67_nl;
  wire[1:0] PECore_DecodeAxiRead_case_4_switch_lp_and_9_nl;
  wire[1:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_10_nl;
  wire[1:0] PEManager_16U_ClusterLookup_for_mux_135_nl;
  wire[2:0] PEManager_16U_ClusterLookup_for_mux_69_nl;
  wire[4:0] PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_12_nl;
  wire[4:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_2_nl;
  wire[4:0] PECore_RunBias_if_for_12_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_12_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_12_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_12_operator_33_true_acc_nl;
  wire[4:0] PEManager_16U_ClusterLookup_for_mux_134_nl;
  wire[5:0] PEManager_16U_ClusterLookup_for_mux_71_nl;
  wire[1:0] PECore_DecodeAxiRead_case_4_switch_lp_and_7_nl;
  wire[1:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_4_nl;
  wire[1:0] PEManager_16U_ClusterLookup_for_mux_133_nl;
  wire[2:0] PEManager_16U_ClusterLookup_for_mux_2_nl;
  wire[4:0] PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_10_nl;
  wire[4:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_nl;
  wire[4:0] PEManager_16U_ClusterLookup_for_mux_132_nl;
  wire[5:0] PEManager_16U_ClusterLookup_for_mux_73_nl;
  wire[1:0] PECore_DecodeAxiRead_case_4_switch_lp_and_6_nl;
  wire[1:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_1_nl;
  wire[1:0] PEManager_16U_ClusterLookup_for_mux_131_nl;
  wire[2:0] PEManager_16U_ClusterLookup_for_mux_75_nl;
  wire[4:0] PEManager_16U_ClusterLookup_for_mux_130_nl;
  wire[4:0] PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_11_nl;
  wire[4:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_1_nl;
  wire[4:0] PECore_RunBias_if_for_2_operator_34_true_acc_nl;
  wire[5:0] nl_PECore_RunBias_if_for_2_operator_34_true_acc_nl;
  wire[2:0] PECore_RunBias_if_for_2_operator_33_true_acc_nl;
  wire[3:0] nl_PECore_RunBias_if_for_2_operator_33_true_acc_nl;
  wire PECore_RunMac_if_and_803_nl;
  wire[3:0] PEManager_16U_ClusterLookup_for_mux_77_nl;
  wire[3:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl;
  wire[3:0] PECore_DecodeAxiRead_case_4_switch_lp_mux1h_24_nl;
  wire[3:0] PEManager_16U_ClusterLookup_for_mux_129_nl;
  wire rva_out_reg_data_and_1_nl;
  wire PECore_RunMac_if_and_801_nl;
  wire PEManager_16U_ClusterLookup_for_mux_79_nl;
  wire[6:0] PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_13_nl;
  wire[6:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl;
  wire[6:0] PEManager_16U_ClusterLookup_for_mux_128_nl;
  wire[3:0] operator_4_false_mux_2_nl;
  wire[2:0] PECore_RunBias_if_for_1_operator_33_true_acc_1_nl;
  wire[3:0] nl_PECore_RunBias_if_for_1_operator_33_true_acc_1_nl;
  wire[7:0] operator_8_false_mux_2_nl;
  wire and_5952_nl;
  wire[13:0] operator_32_true_acc_nl;
  wire[14:0] nl_operator_32_true_acc_nl;
  wire[12:0] operator_32_true_mux1h_40_nl;
  wire[13:0] operator_32_true_acc_1_nl;
  wire[14:0] nl_operator_32_true_acc_1_nl;
  wire[12:0] operator_32_true_mux1h_41_nl;
  wire[13:0] operator_32_true_acc_2_nl;
  wire[14:0] nl_operator_32_true_acc_2_nl;
  wire[12:0] operator_32_true_mux1h_42_nl;
  wire[13:0] operator_32_true_acc_3_nl;
  wire[14:0] nl_operator_32_true_acc_3_nl;
  wire[12:0] operator_32_true_mux1h_43_nl;
  wire[19:0] adpfloat_tmp_to_fixed_20U_14U_if_1_adpfloat_tmp_to_fixed_20U_14U_if_1_mux_2_nl;
  wire[19:0] adpfloat_tmp_to_fixed_20U_14U_if_1_mux1h_8_nl;
  wire[19:0] adpfloat_tmp_to_fixed_20U_14U_if_1_adpfloat_tmp_to_fixed_20U_14U_if_1_mux_3_nl;
  wire[19:0] adpfloat_tmp_to_fixed_20U_14U_if_1_mux1h_9_nl;
  wire[32:0] operator_32_true_acc_nl_1;
  wire[33:0] nl_operator_32_true_acc_nl_1;
  wire[31:0] operator_32_true_mux1h_8_nl;
  wire[32:0] operator_32_true_acc_1_nl_1;
  wire[33:0] nl_operator_32_true_acc_1_nl_1;
  wire[31:0] operator_32_true_mux1h_9_nl;
  wire[32:0] operator_32_true_acc_2_nl_1;
  wire[33:0] nl_operator_32_true_acc_2_nl_1;
  wire[31:0] operator_32_true_mux1h_10_nl;
  wire[32:0] operator_32_true_acc_3_nl_1;
  wire[33:0] nl_operator_32_true_acc_3_nl_1;
  wire[31:0] operator_32_true_mux1h_11_nl;
  wire[31:0] PECore_RunMac_if_for_mux1h_4_nl;
  wire[31:0] PECore_RunMac_if_for_mux1h_5_nl;
  wire[31:0] PECore_RunMac_if_for_mux1h_6_nl;
  wire[31:0] PECore_RunMac_if_for_mux1h_7_nl;
  wire[19:0] and_5953_nl;
  wire[19:0] mux1h_16_nl;
  wire[19:0] PECore_RunBias_if_for_if_or_8_nl;
  wire[19:0] PECore_RunBias_if_for_if_mux1h_4_nl;
  wire PECore_RunBias_if_for_if_and_8_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_8_nl;
  wire PECore_RunBias_if_for_if_or_9_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_12_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_13_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_14_nl;
  wire nor_599_nl;
  wire[19:0] and_5961_nl;
  wire[19:0] mux_645_nl;
  wire[19:0] PECore_RunBias_if_for_if_or_10_nl;
  wire[19:0] PECore_RunBias_if_for_if_mux1h_5_nl;
  wire PECore_RunBias_if_for_if_and_9_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_9_nl;
  wire PECore_RunBias_if_for_if_and_10_nl;
  wire or_3882_nl;
  wire nor_603_nl;
  wire[19:0] and_5968_nl;
  wire[19:0] mux_646_nl;
  wire[19:0] PECore_RunBias_if_for_if_or_11_nl;
  wire[19:0] PECore_RunBias_if_for_if_mux1h_6_nl;
  wire PECore_RunBias_if_for_if_and_11_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_10_nl;
  wire PECore_RunBias_if_for_if_and_12_nl;
  wire or_3883_nl;
  wire nor_607_nl;
  wire[19:0] and_5975_nl;
  wire[19:0] mux_647_nl;
  wire[19:0] PECore_RunBias_if_for_if_or_12_nl;
  wire[19:0] PECore_RunBias_if_for_if_mux1h_7_nl;
  wire PECore_RunBias_if_for_if_and_13_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_11_nl;
  wire PECore_RunBias_if_for_if_and_14_nl;
  wire or_3884_nl;
  wire nor_611_nl;
  wire[2:0] operator_3_false_mux_2_nl;
  wire[2:0] PECore_RunBias_if_right_shift_mux_2_nl;
  wire[2:0] operator_3_false_mux_3_nl;
  wire[2:0] PECore_RunBias_if_right_shift_mux_3_nl;
  wire and_5982_nl;
  wire PEManager_16U_GetInputAddr_1_PEManager_16U_GetInputAddr_1_nor_nl;
  wire PEManager_16U_GetInputAddr_1_and_1_nl;
  wire PEManager_16U_GetInputAddr_1_and_2_nl;
  wire PEManager_16U_GetInputAddr_1_and_3_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_adpfloat_tmp_to_fixed_20U_14U_nor_8_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_16_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_17_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_18_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_adpfloat_tmp_to_fixed_20U_14U_nor_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_20_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_21_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_22_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_23_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_24_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_25_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_26_nl;
  wire adpfloat_tmp_to_fixed_20U_14U_and_27_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[7:0] PECore_RunMac_if_mux1h_63_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_127_nl;
  wire[7:0] PECore_RunMac_if_mux1h_62_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_126_nl;
  wire[7:0] PECore_RunMac_if_mux1h_61_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_124_nl;
  wire[7:0] PECore_RunMac_if_mux1h_60_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_122_nl;
  wire[7:0] PECore_RunMac_if_mux1h_59_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_120_nl;
  wire[7:0] PECore_RunMac_if_mux1h_58_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_118_nl;
  wire[7:0] PECore_RunMac_if_mux1h_57_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_116_nl;
  wire[7:0] PECore_RunMac_if_mux1h_56_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_114_nl;
  wire[7:0] PECore_RunMac_if_mux1h_55_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_112_nl;
  wire[7:0] PECore_RunMac_if_mux1h_54_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_113_nl;
  wire[7:0] PECore_RunMac_if_mux1h_53_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_115_nl;
  wire[7:0] PECore_RunMac_if_mux1h_52_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_117_nl;
  wire[7:0] PECore_RunMac_if_mux1h_51_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_119_nl;
  wire[7:0] PECore_RunMac_if_mux1h_50_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_121_nl;
  wire[7:0] PECore_RunMac_if_mux1h_49_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_123_nl;
  wire[7:0] PECore_RunMac_if_mux1h_48_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_125_nl;
  wire [127:0] nl_Datapath_for_1_ProductSum_cmp_in_1_data_rsc_dat;
  
  wire[7:0] PECore_RunMac_if_mux1h_47_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_111_nl;
  wire[7:0] PECore_RunMac_if_mux1h_46_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_109_nl;
  wire[7:0] PECore_RunMac_if_mux1h_45_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_107_nl;
  wire[7:0] PECore_RunMac_if_mux1h_44_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_105_nl;
  wire[7:0] PECore_RunMac_if_mux1h_43_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_103_nl;
  wire[7:0] PECore_RunMac_if_mux1h_42_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_101_nl;
  wire[7:0] PECore_RunMac_if_mux1h_41_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_99_nl;
  wire[7:0] PECore_RunMac_if_mux1h_40_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_97_nl;
  wire[7:0] PECore_RunMac_if_mux1h_39_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_96_nl;
  wire[7:0] PECore_RunMac_if_mux1h_38_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_98_nl;
  wire[7:0] PECore_RunMac_if_mux1h_37_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_100_nl;
  wire[7:0] PECore_RunMac_if_mux1h_36_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_102_nl;
  wire[7:0] PECore_RunMac_if_mux1h_35_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_104_nl;
  wire[7:0] PECore_RunMac_if_mux1h_34_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_106_nl;
  wire[7:0] PECore_RunMac_if_mux1h_33_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_108_nl;
  wire[7:0] PECore_RunMac_if_mux1h_32_nl;
  wire[7:0] PEManager_16U_ClusterLookup_1_for_mux_110_nl;
  wire [127:0] nl_Datapath_for_1_ProductSum_cmp_1_in_1_data_rsc_dat;

  always @(posedge clk) begin 
    if (~rst) begin
      pe_config_input_counter_sva <= 0;
    end
    else begin
      pe_config_input_counter_sva <= 1;
    end
  end
    


endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore
// ------------------------------------------------------------------


module PECore (
  clk, rst, start_val, start_rdy, start_msg, input_port_val, input_port_rdy, input_port_msg,
      rva_in_val, rva_in_rdy, rva_in_msg, rva_out_val, rva_out_rdy, rva_out_msg,
      act_port_val, act_port_rdy, act_port_msg, SC_SRAM_CONFIG
);
  input clk;
  input rst;
  input start_val;
  output start_rdy;
  input start_msg;
  input input_port_val;
  output input_port_rdy;
  input [137:0] input_port_msg;
  input rva_in_val;
  output rva_in_rdy;
  input [168:0] rva_in_msg;
  output rva_out_val;
  input rva_out_rdy;
  output [127:0] rva_out_msg;
  output act_port_val;
  input act_port_rdy;
  output [319:0] act_port_msg;
  input [31:0] SC_SRAM_CONFIG;


  // Interconnect Declarations
  wire weight_mem_banks_bank_array_impl_data0_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data0_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data0_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data0_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data1_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data1_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data1_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data1_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data1_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data2_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data2_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data2_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data2_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data2_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data3_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data3_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data3_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data3_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data3_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data4_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data4_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data4_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data4_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data4_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data5_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data5_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data5_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data5_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data5_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data6_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data6_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data6_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data6_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data6_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data7_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data7_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data7_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data7_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data7_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data8_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data8_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data8_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data8_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data8_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data9_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data9_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data9_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data9_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data9_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data10_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data10_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data10_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data10_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data10_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data11_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data11_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data11_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data11_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data11_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data12_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data12_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data12_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data12_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data12_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data13_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data13_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data13_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data13_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data13_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data14_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data14_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data14_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data14_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data14_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data15_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data15_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_array_impl_data15_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data15_rsci_radr_d;
  wire weight_mem_banks_bank_array_impl_data15_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire input_mem_banks_bank_array_impl_data0_rsci_clken_d;
  wire [127:0] input_mem_banks_bank_array_impl_data0_rsci_d_d;
  wire [127:0] input_mem_banks_bank_array_impl_data0_rsci_q_d;
  wire [7:0] input_mem_banks_bank_array_impl_data0_rsci_radr_d;
  wire [7:0] input_mem_banks_bank_array_impl_data0_rsci_wadr_d;
  wire input_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire weight_mem_banks_bank_array_impl_data0_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data0_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data0_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data0_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data0_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data0_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data1_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data1_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data1_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data1_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data1_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data1_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data2_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data2_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data2_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data2_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data2_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data2_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data3_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data3_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data3_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data3_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data3_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data3_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data4_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data4_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data4_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data4_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data4_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data4_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data5_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data5_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data5_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data5_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data5_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data5_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data6_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data6_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data6_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data6_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data6_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data6_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data7_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data7_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data7_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data7_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data7_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data7_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data8_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data8_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data8_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data8_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data8_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data8_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data9_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data9_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data9_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data9_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data9_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data9_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data10_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data10_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data10_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data10_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data10_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data10_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data11_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data11_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data11_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data11_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data11_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data11_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data12_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data12_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data12_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data12_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data12_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data12_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data13_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data13_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data13_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data13_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data13_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data13_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data14_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data14_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data14_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data14_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data14_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data14_rsc_wadr;
  wire weight_mem_banks_bank_array_impl_data15_rsc_clken;
  wire [127:0] weight_mem_banks_bank_array_impl_data15_rsc_q;
  wire [11:0] weight_mem_banks_bank_array_impl_data15_rsc_radr;
  wire weight_mem_banks_bank_array_impl_data15_rsc_we;
  wire [127:0] weight_mem_banks_bank_array_impl_data15_rsc_d;
  wire [11:0] weight_mem_banks_bank_array_impl_data15_rsc_wadr;
  wire input_mem_banks_bank_array_impl_data0_rsc_clken;
  wire [127:0] input_mem_banks_bank_array_impl_data0_rsc_q;
  wire [7:0] input_mem_banks_bank_array_impl_data0_rsc_radr;
  wire input_mem_banks_bank_array_impl_data0_rsc_we;
  wire [127:0] input_mem_banks_bank_array_impl_data0_rsc_d;
  wire [7:0] input_mem_banks_bank_array_impl_data0_rsc_wadr;
  wire [11:0] weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_iff;
  wire weight_mem_banks_bank_array_impl_data0_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data1_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data2_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data3_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data4_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data5_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data6_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data7_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data8_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data9_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data10_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data11_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data12_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data13_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data14_rsci_we_d_iff;
  wire weight_mem_banks_bank_array_impl_data15_rsci_we_d_iff;
  wire input_mem_banks_bank_array_impl_data0_rsci_we_d_iff;

  // Helper signals
  wire [2:0] state;
  assign state = {PECore_PECoreRun_inst.state_2_0_sva_2, PECore_PECoreRun_inst.state_2_0_sva_1, PECore_PECoreRun_inst.state_2_0_sva_0};

  wire is_start;
  assign is_start = PECore_PECoreRun_inst.is_start_sva;

  // PE_Config signals
  wire pe_config_is_valid = PECore_PECoreRun_inst.pe_config_is_valid_sva;
  wire pe_config_is_zero_first = PECore_PECoreRun_inst.pe_config_is_zero_first_sva;
  wire pe_config_is_cluster = PECore_PECoreRun_inst.pe_config_is_cluster_sva;
  wire pe_config_is_bias = PECore_PECoreRun_inst.pe_config_is_bias_sva;
  wire [3:0] pe_config_num_manager = PECore_PECoreRun_inst.pe_config_num_manager_sva;
  wire [7:0] pe_config_num_output = PECore_PECoreRun_inst.pe_config_num_output_sva;
  wire pe_config_manager_counter = PECore_PECoreRun_inst.pe_config_manager_counter_sva;
  wire [7:0] pe_config_input_counter = PECore_PECoreRun_inst.pe_config_input_counter_sva;
  wire [7:0] pe_config_output_counter = PECore_PECoreRun_inst.pe_config_output_counter_sva;

  // RVA_IN Decode
  wire rva_in_rw = rva_in_msg[168];
  wire [15:0] rva_in_wstrb = rva_in_msg[167:152];
  wire [23:0] rva_in_addr = rva_in_msg[151:128];
  wire [127:0] rva_in_data = rva_in_msg[127:0];

  
  PECore_PECore_PECoreRun PECore_PECoreRun_inst (
      .clk(clk),
      .rst(rst),
      .start_val(start_val),
      .start_rdy(start_rdy),
      .start_msg(start_msg),
      .input_port_val(input_port_val),
      .input_port_rdy(input_port_rdy),
      .input_port_msg(input_port_msg),
      .rva_in_val(rva_in_val),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_msg(rva_in_msg),
      .rva_out_val(rva_out_val),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_msg(rva_out_msg),
      .act_port_val(act_port_val),
      .act_port_rdy(act_port_rdy),
      .act_port_msg(act_port_msg),
      .SC_SRAM_CONFIG(SC_SRAM_CONFIG),
      .weight_mem_banks_bank_array_impl_data0_rsci_clken_d(weight_mem_banks_bank_array_impl_data0_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data0_rsci_d_d(weight_mem_banks_bank_array_impl_data0_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data0_rsci_q_d(weight_mem_banks_bank_array_impl_data0_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data0_rsci_radr_d(weight_mem_banks_bank_array_impl_data0_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data1_rsci_clken_d(weight_mem_banks_bank_array_impl_data1_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data1_rsci_d_d(weight_mem_banks_bank_array_impl_data1_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data1_rsci_q_d(weight_mem_banks_bank_array_impl_data1_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data1_rsci_radr_d(weight_mem_banks_bank_array_impl_data1_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data1_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data1_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data2_rsci_clken_d(weight_mem_banks_bank_array_impl_data2_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data2_rsci_d_d(weight_mem_banks_bank_array_impl_data2_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data2_rsci_q_d(weight_mem_banks_bank_array_impl_data2_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data2_rsci_radr_d(weight_mem_banks_bank_array_impl_data2_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data2_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data2_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data3_rsci_clken_d(weight_mem_banks_bank_array_impl_data3_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data3_rsci_d_d(weight_mem_banks_bank_array_impl_data3_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data3_rsci_q_d(weight_mem_banks_bank_array_impl_data3_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data3_rsci_radr_d(weight_mem_banks_bank_array_impl_data3_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data3_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data3_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data4_rsci_clken_d(weight_mem_banks_bank_array_impl_data4_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data4_rsci_d_d(weight_mem_banks_bank_array_impl_data4_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data4_rsci_q_d(weight_mem_banks_bank_array_impl_data4_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data4_rsci_radr_d(weight_mem_banks_bank_array_impl_data4_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data4_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data4_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data5_rsci_clken_d(weight_mem_banks_bank_array_impl_data5_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data5_rsci_d_d(weight_mem_banks_bank_array_impl_data5_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data5_rsci_q_d(weight_mem_banks_bank_array_impl_data5_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data5_rsci_radr_d(weight_mem_banks_bank_array_impl_data5_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data5_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data5_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data6_rsci_clken_d(weight_mem_banks_bank_array_impl_data6_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data6_rsci_d_d(weight_mem_banks_bank_array_impl_data6_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data6_rsci_q_d(weight_mem_banks_bank_array_impl_data6_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data6_rsci_radr_d(weight_mem_banks_bank_array_impl_data6_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data6_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data6_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data7_rsci_clken_d(weight_mem_banks_bank_array_impl_data7_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data7_rsci_d_d(weight_mem_banks_bank_array_impl_data7_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data7_rsci_q_d(weight_mem_banks_bank_array_impl_data7_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data7_rsci_radr_d(weight_mem_banks_bank_array_impl_data7_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data7_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data7_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data8_rsci_clken_d(weight_mem_banks_bank_array_impl_data8_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data8_rsci_d_d(weight_mem_banks_bank_array_impl_data8_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data8_rsci_q_d(weight_mem_banks_bank_array_impl_data8_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data8_rsci_radr_d(weight_mem_banks_bank_array_impl_data8_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data8_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data8_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data9_rsci_clken_d(weight_mem_banks_bank_array_impl_data9_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data9_rsci_d_d(weight_mem_banks_bank_array_impl_data9_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data9_rsci_q_d(weight_mem_banks_bank_array_impl_data9_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data9_rsci_radr_d(weight_mem_banks_bank_array_impl_data9_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data9_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data9_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data10_rsci_clken_d(weight_mem_banks_bank_array_impl_data10_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data10_rsci_d_d(weight_mem_banks_bank_array_impl_data10_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data10_rsci_q_d(weight_mem_banks_bank_array_impl_data10_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data10_rsci_radr_d(weight_mem_banks_bank_array_impl_data10_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data10_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data10_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data11_rsci_clken_d(weight_mem_banks_bank_array_impl_data11_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data11_rsci_d_d(weight_mem_banks_bank_array_impl_data11_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data11_rsci_q_d(weight_mem_banks_bank_array_impl_data11_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data11_rsci_radr_d(weight_mem_banks_bank_array_impl_data11_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data11_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data11_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data12_rsci_clken_d(weight_mem_banks_bank_array_impl_data12_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data12_rsci_d_d(weight_mem_banks_bank_array_impl_data12_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data12_rsci_q_d(weight_mem_banks_bank_array_impl_data12_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data12_rsci_radr_d(weight_mem_banks_bank_array_impl_data12_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data12_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data12_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data13_rsci_clken_d(weight_mem_banks_bank_array_impl_data13_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data13_rsci_d_d(weight_mem_banks_bank_array_impl_data13_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data13_rsci_q_d(weight_mem_banks_bank_array_impl_data13_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data13_rsci_radr_d(weight_mem_banks_bank_array_impl_data13_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data13_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data13_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data14_rsci_clken_d(weight_mem_banks_bank_array_impl_data14_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data14_rsci_d_d(weight_mem_banks_bank_array_impl_data14_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data14_rsci_q_d(weight_mem_banks_bank_array_impl_data14_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data14_rsci_radr_d(weight_mem_banks_bank_array_impl_data14_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data14_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data14_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data15_rsci_clken_d(weight_mem_banks_bank_array_impl_data15_rsci_clken_d),
      .weight_mem_banks_bank_array_impl_data15_rsci_d_d(weight_mem_banks_bank_array_impl_data15_rsci_d_d),
      .weight_mem_banks_bank_array_impl_data15_rsci_q_d(weight_mem_banks_bank_array_impl_data15_rsci_q_d),
      .weight_mem_banks_bank_array_impl_data15_rsci_radr_d(weight_mem_banks_bank_array_impl_data15_rsci_radr_d),
      .weight_mem_banks_bank_array_impl_data15_rsci_readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_array_impl_data15_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .input_mem_banks_bank_array_impl_data0_rsci_clken_d(input_mem_banks_bank_array_impl_data0_rsci_clken_d),
      .input_mem_banks_bank_array_impl_data0_rsci_d_d(input_mem_banks_bank_array_impl_data0_rsci_d_d),
      .input_mem_banks_bank_array_impl_data0_rsci_q_d(input_mem_banks_bank_array_impl_data0_rsci_q_d),
      .input_mem_banks_bank_array_impl_data0_rsci_radr_d(input_mem_banks_bank_array_impl_data0_rsci_radr_d),
      .input_mem_banks_bank_array_impl_data0_rsci_wadr_d(input_mem_banks_bank_array_impl_data0_rsci_wadr_d),
      .input_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d(input_mem_banks_bank_array_impl_data0_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_pff(weight_mem_banks_bank_array_impl_data0_rsci_wadr_d_iff),
      .weight_mem_banks_bank_array_impl_data0_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data0_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data1_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data1_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data2_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data2_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data3_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data3_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data4_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data4_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data5_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data5_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data6_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data6_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data7_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data7_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data8_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data8_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data9_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data9_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data10_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data10_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data11_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data11_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data12_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data12_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data13_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data13_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data14_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data14_rsci_we_d_iff),
      .weight_mem_banks_bank_array_impl_data15_rsci_we_d_pff(weight_mem_banks_bank_array_impl_data15_rsci_we_d_iff),
      .input_mem_banks_bank_array_impl_data0_rsci_we_d_pff(input_mem_banks_bank_array_impl_data0_rsci_we_d_iff)
    );
endmodule