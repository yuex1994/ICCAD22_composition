// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun (
  clk, rst, start_val, start_rdy, start_msg, act_port_val, act_port_rdy, act_port_msg,
      rva_in_val, rva_in_rdy, rva_in_msg, rva_out_val, rva_out_rdy, rva_out_msg,
      output_port_val, output_port_rdy, output_port_msg, done_val, done_rdy, done_msg
);
  input clk;
  input rst;
  input start_val;
  output start_rdy;
  input start_msg;
  input act_port_val;
  output act_port_rdy;
  input [319:0] act_port_msg;
  input rva_in_val;
  output rva_in_rdy;
  input [168:0] rva_in_msg;
  output rva_out_val;
  input rva_out_rdy;
  output [127:0] rva_out_msg;
  output output_port_val;
  input output_port_rdy;
  output [137:0] output_port_msg;
  output done_val;
  input done_rdy;
  output done_msg;


  // Interconnect Declarations
  wire ActUnitRun_wen;
  wire ActUnitRun_wten;
  wire [127:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  wire [11:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_return_rsc_z_mxwt;
  wire [319:0] act_port_PopNB_mioi_data_data_rsc_z_mxwt;
  wire act_port_PopNB_mioi_return_rsc_z_mxwt;
  wire rva_out_Push_mioi_wen_comp;
  wire start_PopNB_mioi_data_rsc_z_mxwt;
  wire start_PopNB_mioi_return_rsc_z_mxwt;
  wire output_port_Push_mioi_wen_comp;
  wire done_Push_mioi_wen_comp;
  wire [2:0] fsm_output;
  wire act_config_InstIncr_if_if_unequal_tmp;
  wire [8:0] operator_8_false_acc_tmp;
  wire [9:0] nl_operator_8_false_acc_tmp;
  wire act_config_InstIncr_if_equal_1_tmp;
  wire [6:0] operator_6_false_acc_tmp;
  wire [7:0] nl_operator_6_false_acc_tmp;
  wire ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_1_tmp;
  wire [7:0] act_config_in_InstFetch_mux_tmp;
  wire [4:0] while_mux_125_tmp;
  wire mux_tmp_1;
  wire and_dcpl;
  wire and_dcpl_1;
  wire and_dcpl_5;
  wire and_dcpl_8;
  wire and_dcpl_11;
  wire or_dcpl_8;
  wire or_dcpl_9;
  wire and_dcpl_31;
  wire nor_tmp_6;
  wire mux_tmp_16;
  wire or_dcpl_13;
  wire or_dcpl_15;
  wire or_dcpl_22;
  wire not_tmp_34;
  wire or_dcpl_27;
  wire and_dcpl_45;
  wire or_dcpl_33;
  wire or_dcpl_34;
  wire or_dcpl_35;
  wire or_dcpl_38;
  wire or_dcpl_41;
  wire or_dcpl_44;
  wire or_dcpl_47;
  wire or_dcpl_56;
  wire or_dcpl_57;
  wire or_dcpl_66;
  wire or_dcpl_75;
  wire or_dcpl_76;
  wire or_dcpl_85;
  wire or_dcpl_94;
  wire or_dcpl_95;
  wire or_dcpl_104;
  wire or_dcpl_116;
  wire and_dcpl_65;
  wire or_tmp_61;
  wire and_158_cse;
  wire act_config_InstIncr_if_act_config_InstIncr_if_if_act_config_InstIncr_if_if_nor_mdf_sva_1;
  wire act_config_InstIncr_act_config_InstIncr_if_and_svs_1;
  wire act_config_ActConfigRead_else_unequal_tmp_1;
  wire act_config_ActConfigRead_unequal_tmp_1;
  wire ActUnit_RunInst_switch_lp_and_66_tmp_1;
  reg ActUnit_RunInst_switch_lp_equal_tmp_2;
  reg is_start_sva;
  wire ActUnit_RunInst_switch_lp_equal_tmp_20;
  reg ActUnit_RunInst_switch_lp_equal_tmp_1;
  reg ActUnit_RunInst_switch_lp_equal_tmp_3;
  reg ActUnit_RunInst_switch_lp_nor_tmp;
  reg ActUnit_RunInst_switch_lp_equal_tmp_4;
  reg ActUnit_RunInst_switch_lp_equal_tmp_5;
  reg ActUnit_RunInst_switch_lp_equal_tmp_6;
  reg ActUnit_RunInst_switch_lp_equal_tmp_7;
  reg ActUnit_RunInst_switch_lp_equal_tmp_8;
  reg ActUnit_RunInst_switch_lp_equal_tmp_9;
  reg ActUnit_RunInst_switch_lp_equal_tmp_10;
  wire ActUnit_RunInst_switch_lp_and_ssc_sva_1;
  wire ActUnit_RunInst_switch_lp_and_50_tmp_1;
  wire ActUnit_RunInst_switch_lp_and_ssc_1_sva_1;
  wire ActUnit_RunInst_switch_lp_and_34_tmp_1;
  wire ActUnit_RunInst_switch_lp_and_ssc_2_sva_1;
  wire ActUnit_RunInst_switch_lp_and_18_tmp_1;
  wire ActUnit_RunInst_switch_lp_nor_ssc_sva_1;
  wire ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0;
  wire ActUnit_RunInst_switch_lp_equal_tmp_11;
  wire ActUnit_RunInst_switch_lp_equal_tmp_12;
  wire ActUnit_RunInst_switch_lp_equal_tmp_13;
  wire ActUnit_RunInst_switch_lp_equal_tmp_14;
  wire ActUnit_RunInst_switch_lp_equal_tmp_15;
  wire ActUnit_RunInst_switch_lp_equal_tmp_16;
  wire ActUnit_RunInst_switch_lp_equal_tmp_17;
  wire ActUnit_RunInst_switch_lp_equal_tmp_18;
  wire ActUnit_RunInst_switch_lp_equal_tmp_19;
  wire ActUnit_RunInst_switch_lp_nor_tmp_1;
  wire is_incr_lpi_1_dfm_2;
  wire ActUnit_RunLoad_if_else_and_ssc_sva_1;
  wire ActUnit_PushOutput_and_tmp_1;
  wire act_config_is_zero_first_sva_dfm_4_mx0;
  wire ActUnit_RunLoad_if_else_and_ssc_1_sva_1;
  wire ActUnit_RunLoad_if_else_and_ssc_2_sva_1;
  wire ActUnit_RunLoad_if_else_nor_ssc_sva_1;
  reg ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_cse;
  reg [4:0] act_config_inst_counter_sva;
  wire [7:0] ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_mx1_tmp_7_0;
  reg act_config_is_valid_sva;
  wire ActUnit_DecodeAxiRead_unequal_tmp_1;
  wire [1:0] nvhls_get_slc_2U_NVUINT8_return_3_sva_1;
  reg [7:0] act_config_inst_regs_0_sva_dfm_5;
  reg [7:0] act_config_inst_regs_1_sva_dfm_5;
  reg [7:0] act_config_inst_regs_2_sva_dfm_5;
  reg [7:0] act_config_inst_regs_3_sva_dfm_5;
  reg [7:0] act_config_inst_regs_4_sva_dfm_5;
  reg [7:0] act_config_inst_regs_5_sva_dfm_5;
  reg [7:0] act_config_inst_regs_6_sva_dfm_5;
  reg [7:0] act_config_inst_regs_7_sva_dfm_5;
  reg [7:0] act_config_inst_regs_8_sva_dfm_5;
  reg [7:0] act_config_inst_regs_9_sva_dfm_5;
  reg [7:0] act_config_inst_regs_10_sva_dfm_5;
  reg [7:0] act_config_inst_regs_11_sva_dfm_5;
  reg [7:0] act_config_inst_regs_12_sva_dfm_5;
  reg [7:0] act_config_inst_regs_13_sva_dfm_5;
  reg [7:0] act_config_inst_regs_14_sva_dfm_5;
  reg [7:0] act_config_inst_regs_15_sva_dfm_5;
  reg [7:0] act_config_inst_regs_16_sva_dfm_6;
  reg [7:0] act_config_inst_regs_17_sva_dfm_6;
  reg [7:0] act_config_inst_regs_18_sva_dfm_6;
  reg [7:0] act_config_inst_regs_19_sva_dfm_6;
  reg [7:0] act_config_inst_regs_20_sva_dfm_6;
  reg [7:0] act_config_inst_regs_21_sva_dfm_6;
  reg [7:0] act_config_inst_regs_22_sva_dfm_6;
  reg [7:0] act_config_inst_regs_23_sva_dfm_6;
  reg [7:0] act_config_inst_regs_24_sva_dfm_6;
  reg [7:0] act_config_inst_regs_25_sva_dfm_6;
  reg [7:0] act_config_inst_regs_26_sva_dfm_6;
  reg [7:0] act_config_inst_regs_27_sva_dfm_6;
  reg [7:0] act_config_inst_regs_28_sva_dfm_6;
  reg [7:0] act_config_inst_regs_29_sva_dfm_6;
  reg [7:0] act_config_inst_regs_30_sva_dfm_6;
  reg [7:0] act_config_inst_regs_31_sva_dfm_6;
  reg [7:0] reg_ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_ftd_12;
  wire act_mem_banks_write_if_for_if_mux_cse;
  wire act_mem_banks_write_if_for_if_mux_1_cse;
  wire act_mem_banks_read_for_mux_16_cse;
  wire act_mem_banks_read_for_mux_17_cse;
  wire ActUnit_DecodeAxiRead_and_9_cse;
  wire ActUnit_DecodeAxiRead_and_10_cse;
  reg reg_done_Push_mioi_iswt0_cse;
  reg reg_output_port_Push_mioi_iswt0_cse;
  reg reg_start_PopNB_mioi_iswt0_cse;
  reg reg_rva_out_Push_mioi_iswt0_cse;
  reg reg_act_port_PopNB_mioi_iswt0_cse;
  reg reg_rva_in_PopNB_mioi_iswt0_cse;
  wire act_regs_data_and_cse;
  wire act_config_adpfloat_bias_and_cse;
  wire act_config_inst_regs_and_cse;
  wire act_config_inst_regs_and_16_cse;
  wire act_mem_banks_bank_array_impl_data0_and_cse;
  wire act_mem_banks_bank_array_impl_data0_and_1_cse;
  wire act_mem_banks_bank_array_impl_data0_and_2_cse;
  wire act_mem_banks_bank_array_impl_data0_and_3_cse;
  wire act_mem_banks_bank_array_impl_data0_and_4_cse;
  wire act_mem_banks_bank_array_impl_data0_and_5_cse;
  wire act_mem_banks_bank_array_impl_data0_and_6_cse;
  wire act_mem_banks_bank_array_impl_data0_and_7_cse;
  wire act_mem_banks_bank_array_impl_data0_and_8_cse;
  wire act_mem_banks_bank_array_impl_data0_and_9_cse;
  wire act_mem_banks_bank_array_impl_data0_and_10_cse;
  wire act_mem_banks_bank_array_impl_data0_and_11_cse;
  wire act_mem_banks_bank_array_impl_data0_and_12_cse;
  wire act_mem_banks_bank_array_impl_data0_and_13_cse;
  wire act_mem_banks_bank_array_impl_data0_and_14_cse;
  wire act_mem_banks_bank_array_impl_data0_and_15_cse;
  wire act_mem_banks_bank_array_impl_data0_and_16_cse;
  wire act_mem_banks_bank_array_impl_data0_and_17_cse;
  wire act_mem_banks_bank_array_impl_data0_and_18_cse;
  wire act_mem_banks_bank_array_impl_data0_and_19_cse;
  wire act_mem_banks_bank_array_impl_data0_and_20_cse;
  wire act_mem_banks_bank_array_impl_data0_and_21_cse;
  wire act_mem_banks_bank_array_impl_data0_and_22_cse;
  wire act_mem_banks_bank_array_impl_data0_and_23_cse;
  wire act_mem_banks_bank_array_impl_data0_and_24_cse;
  wire act_mem_banks_bank_array_impl_data0_and_25_cse;
  wire act_mem_banks_bank_array_impl_data0_and_26_cse;
  wire act_mem_banks_bank_array_impl_data0_and_27_cse;
  wire act_mem_banks_bank_array_impl_data0_and_28_cse;
  wire act_mem_banks_bank_array_impl_data0_and_29_cse;
  wire act_mem_banks_bank_array_impl_data0_and_30_cse;
  wire act_mem_banks_bank_array_impl_data0_and_31_cse;
  wire act_mem_banks_read_read_data_and_cse;
  wire or_55_cse;
  wire or_58_cse;
  wire ActUnit_CheckStart_if_ActUnit_CheckStart_if_and_1_cse;
  wire ActUnit_RunInst_switch_lp_nor_13_cse;
  wire or_16_cse;
  wire mux_5_cse;
  wire act_port_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct_mx0;
  wire rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct_mx0;
  reg [7:0] act_config_output_counter_sva;
  reg [7:0] act_config_output_addr_base_sva;
  wire output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct_mx0;
  wire done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct_mx0;
  wire [7:0] act_mem_banks_read_for_mux_mx0w0;
  wire act_config_ActConfigRead_else_else_not_22;
  wire [7:0] act_mem_banks_read_for_mux_1_mx0w0;
  wire [7:0] act_mem_banks_read_for_mux_2_mx0w0;
  wire [7:0] act_mem_banks_read_for_mux_3_mx0w0;
  wire [7:0] act_mem_banks_read_for_mux_4_mx0w0;
  wire [7:0] act_mem_banks_read_for_mux_5_mx0w0;
  wire [7:0] act_mem_banks_read_for_mux_6_mx0w0;
  wire [7:0] act_mem_banks_read_for_mux_7_mx0w0;
  wire ActUnit_DecodeAxiRead_and_cse_1;
  wire [7:0] act_mem_banks_read_for_mux_8_mx0w0;
  wire [7:0] act_mem_banks_read_for_mux_9_mx0w0;
  reg [4:0] act_config_buffer_addr_base_sva;
  wire [7:0] act_mem_banks_read_for_mux_10_mx0w0;
  wire [7:0] act_mem_banks_read_for_mux_11_mx0w0;
  reg [7:0] act_config_num_output_sva;
  wire [7:0] act_mem_banks_read_for_mux_12_mx0w0;
  reg [5:0] act_config_num_inst_sva;
  wire [7:0] act_mem_banks_read_for_mux_13_mx0w0;
  reg [2:0] act_config_adpfloat_bias_sva;
  wire [7:0] act_mem_banks_read_for_mux_14_mx0w0;
  reg act_config_is_zero_first_sva;
  reg act_config_inst_regs_1_sva_0;
  reg act_config_inst_regs_17_sva_0;
  wire [7:0] act_mem_banks_read_for_mux_15_mx0w0;
  reg ActUnit_RunInst_switch_lp_nor_7_itm;
  reg act_config_inst_regs_16_sva_0;
  wire or_dcpl;
  wire or_dcpl_122;
  wire or_dcpl_123;
  wire or_dcpl_124;
  wire and_tmp;
  wire and_dcpl_73;
  wire while_asn_1364;
  wire while_asn_1378;
  wire [19:0] act_regs_data_0_15_sva_dfm_3;
  wire while_asn_1374;
  wire [19:0] act_regs_data_1_15_sva_dfm_3;
  wire while_asn_1370;
  wire [19:0] act_regs_data_2_15_sva_dfm_3;
  wire while_asn_1366;
  wire [19:0] act_regs_data_3_15_sva_dfm_3;
  wire [19:0] act_regs_data_0_14_sva_dfm_3;
  wire [19:0] act_regs_data_1_14_sva_dfm_3;
  wire [19:0] act_regs_data_2_14_sva_dfm_3;
  wire [19:0] act_regs_data_3_14_sva_dfm_3;
  wire [19:0] act_regs_data_0_13_sva_dfm_3;
  wire [19:0] act_regs_data_1_13_sva_dfm_3;
  wire [19:0] act_regs_data_2_13_sva_dfm_3;
  wire [19:0] act_regs_data_3_13_sva_dfm_3;
  wire [19:0] act_regs_data_0_12_sva_dfm_3;
  wire [19:0] act_regs_data_1_12_sva_dfm_3;
  wire [19:0] act_regs_data_2_12_sva_dfm_3;
  wire [19:0] act_regs_data_3_12_sva_dfm_3;
  wire [19:0] act_regs_data_0_11_sva_dfm_3;
  wire [19:0] act_regs_data_1_11_sva_dfm_3;
  wire [19:0] act_regs_data_2_11_sva_dfm_3;
  wire [19:0] act_regs_data_3_11_sva_dfm_3;
  wire [19:0] act_regs_data_0_10_sva_dfm_3;
  wire [19:0] act_regs_data_1_10_sva_dfm_3;
  wire [19:0] act_regs_data_2_10_sva_dfm_3;
  wire [19:0] act_regs_data_3_10_sva_dfm_3;
  wire [19:0] act_regs_data_0_9_sva_dfm_3;
  wire [19:0] act_regs_data_1_9_sva_dfm_3;
  wire [19:0] act_regs_data_2_9_sva_dfm_3;
  wire [19:0] act_regs_data_3_9_sva_dfm_3;
  wire [19:0] act_regs_data_0_8_sva_dfm_3;
  wire [19:0] act_regs_data_1_8_sva_dfm_3;
  wire [19:0] act_regs_data_2_8_sva_dfm_3;
  wire [19:0] act_regs_data_3_8_sva_dfm_3;
  wire [19:0] act_regs_data_0_7_sva_dfm_3;
  wire [19:0] act_regs_data_1_7_sva_dfm_3;
  wire [19:0] act_regs_data_2_7_sva_dfm_3;
  wire [19:0] act_regs_data_3_7_sva_dfm_3;
  wire [19:0] act_regs_data_0_6_sva_dfm_3;
  wire [19:0] act_regs_data_1_6_sva_dfm_3;
  wire [19:0] act_regs_data_2_6_sva_dfm_3;
  wire [19:0] act_regs_data_3_6_sva_dfm_3;
  wire [19:0] act_regs_data_0_5_sva_dfm_3;
  wire [19:0] act_regs_data_1_5_sva_dfm_3;
  wire [19:0] act_regs_data_2_5_sva_dfm_3;
  wire [19:0] act_regs_data_3_5_sva_dfm_3;
  wire [19:0] act_regs_data_0_4_sva_dfm_3;
  wire [19:0] act_regs_data_1_4_sva_dfm_3;
  wire [19:0] act_regs_data_2_4_sva_dfm_3;
  wire [19:0] act_regs_data_3_4_sva_dfm_3;
  wire [19:0] act_regs_data_0_3_sva_dfm_3;
  wire [19:0] act_regs_data_1_3_sva_dfm_3;
  wire [19:0] act_regs_data_2_3_sva_dfm_3;
  wire [19:0] act_regs_data_3_3_sva_dfm_3;
  wire [19:0] act_regs_data_0_2_sva_dfm_3;
  wire [19:0] act_regs_data_1_2_sva_dfm_3;
  wire [19:0] act_regs_data_2_2_sva_dfm_3;
  wire [19:0] act_regs_data_3_2_sva_dfm_3;
  wire [19:0] act_regs_data_0_1_sva_dfm_3;
  wire [19:0] act_regs_data_1_1_sva_dfm_3;
  wire [19:0] act_regs_data_2_1_sva_dfm_3;
  wire [19:0] act_regs_data_3_1_sva_dfm_3;
  wire [19:0] act_regs_data_0_0_sva_dfm_3;
  wire [19:0] act_regs_data_1_0_sva_dfm_3;
  wire [19:0] act_regs_data_2_0_sva_dfm_3;
  wire [19:0] act_regs_data_3_0_sva_dfm_3;
  wire act_config_output_counter_sva_mx0c1;
  wire or_887_tmp;
  reg [319:0] ActUnit_RunInst_case_8_EAdd_act_regs_data_sva;
  reg [319:0] ActUnit_RunInst_case_9_EMul_act_regs_data_sva;
  reg [319:0] ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva;
  reg [319:0] ActUnit_RunInst_case_11_Tanh_act_regs_data_sva;
  reg [319:0] ActUnit_RunInst_case_12_Relu_act_regs_data_sva;
  reg [319:0] ActUnit_RunInst_case_13_OneX_act_regs_data_sva;
  wire and_1551_tmp;
  wire nor_18_cse;
  wire nor_19_cse;
  wire nor_20_cse;
  wire nor_21_cse;
  wire or_884_itm;
  wire [127:0] out_data_out;
  wire or_tmp_756;
  reg [19:0] act_regs_data_1_15_sva;
  reg [19:0] act_regs_data_2_0_sva;
  reg [19:0] act_regs_data_1_14_sva;
  reg [19:0] act_regs_data_2_1_sva;
  reg [19:0] act_regs_data_1_13_sva;
  reg [19:0] act_regs_data_2_2_sva;
  reg [19:0] act_regs_data_1_12_sva;
  reg [19:0] act_regs_data_2_3_sva;
  reg [19:0] act_regs_data_1_11_sva;
  reg [19:0] act_regs_data_2_4_sva;
  reg [19:0] act_regs_data_1_10_sva;
  reg [19:0] act_regs_data_2_5_sva;
  reg [19:0] act_regs_data_1_9_sva;
  reg [19:0] act_regs_data_2_6_sva;
  reg [19:0] act_regs_data_1_8_sva;
  reg [19:0] act_regs_data_2_7_sva;
  reg [19:0] act_regs_data_1_7_sva;
  reg [19:0] act_regs_data_2_8_sva;
  reg [19:0] act_regs_data_1_6_sva;
  reg [19:0] act_regs_data_2_9_sva;
  reg [19:0] act_regs_data_1_5_sva;
  reg [19:0] act_regs_data_2_10_sva;
  reg [19:0] act_regs_data_1_4_sva;
  reg [19:0] act_regs_data_2_11_sva;
  reg [19:0] act_regs_data_1_3_sva;
  reg [19:0] act_regs_data_2_12_sva;
  reg [19:0] act_regs_data_1_2_sva;
  reg [19:0] act_regs_data_2_13_sva;
  reg [19:0] act_regs_data_1_1_sva;
  reg [19:0] act_regs_data_2_14_sva;
  reg [19:0] act_regs_data_1_0_sva;
  reg [19:0] act_regs_data_2_15_sva;
  reg [19:0] act_regs_data_0_15_sva;
  reg [19:0] act_regs_data_3_0_sva;
  reg [19:0] act_regs_data_0_14_sva;
  reg [19:0] act_regs_data_3_1_sva;
  reg [19:0] act_regs_data_0_13_sva;
  reg [19:0] act_regs_data_3_2_sva;
  reg [19:0] act_regs_data_0_12_sva;
  reg [19:0] act_regs_data_3_3_sva;
  reg [19:0] act_regs_data_0_11_sva;
  reg [19:0] act_regs_data_3_4_sva;
  reg [19:0] act_regs_data_0_10_sva;
  reg [19:0] act_regs_data_3_5_sva;
  reg [19:0] act_regs_data_0_9_sva;
  reg [19:0] act_regs_data_3_6_sva;
  reg [19:0] act_regs_data_0_8_sva;
  reg [19:0] act_regs_data_3_7_sva;
  reg [19:0] act_regs_data_0_7_sva;
  reg [19:0] act_regs_data_3_8_sva;
  reg [19:0] act_regs_data_0_6_sva;
  reg [19:0] act_regs_data_3_9_sva;
  reg [19:0] act_regs_data_0_5_sva;
  reg [19:0] act_regs_data_3_10_sva;
  reg [19:0] act_regs_data_0_4_sva;
  reg [19:0] act_regs_data_3_11_sva;
  reg [19:0] act_regs_data_0_3_sva;
  reg [19:0] act_regs_data_3_12_sva;
  reg [19:0] act_regs_data_0_2_sva;
  reg [19:0] act_regs_data_3_13_sva;
  reg [19:0] act_regs_data_0_1_sva;
  reg [19:0] act_regs_data_3_14_sva;
  reg [19:0] act_regs_data_0_0_sva;
  reg [19:0] act_regs_data_3_15_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [4:0] act_read_addrs_lpi_1_dfm_5;
  reg [7:0] act_write_data_data_0_0_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_1_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_2_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_3_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_4_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_5_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_6_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_7_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_8_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_9_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_10_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_11_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_12_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_13_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_14_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_15_lpi_1_dfm_4;
  reg [4:0] act_write_addrs_lpi_1_dfm_5;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_7_0_sva_dfm;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_127_120;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_119_112;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_111_104;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_103_96;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_95_88;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_87_80;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_79_72;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_71_64;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_63_56;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_55_48;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_47_40;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_39_32;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_31_24;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_23_16;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_15_8;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_7_0;
  wire act_config_is_valid_sva_mx0c0;
  wire ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0;
  wire is_start_sva_mx0c1;
  wire [4:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_3_mx0w2;
  wire act_write_addrs_lpi_1_dfm_5_mx0c2;
  wire ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_cse_1;
  wire ActUnit_RunInst_switch_lp_nor_7_itm_mx0w0;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [4:0] while_mux_124_ssc_mx0;
  wire [4:0] act_read_addrs_lpi_1_dfm_9;
  wire [7:0] act_write_data_data_0_0_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_1_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_2_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_3_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_4_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_5_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_6_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_7_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_8_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_9_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_10_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_11_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_12_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_13_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_14_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_15_lpi_1_dfm_5_mx0;
  wire while_asn_1290;
  wire while_asn_1292;
  wire while_asn_1294;
  wire while_asn_1296;
  wire while_asn_1298;
  wire while_asn_1300;
  wire while_asn_1302;
  wire while_asn_1304;
  wire while_asn_1306;
  wire while_asn_1308;
  wire while_asn_1310;
  wire while_asn_1312;
  wire while_asn_1314;
  wire while_asn_1316;
  wire while_asn_1318;
  wire while_asn_1320;
  wire while_asn_1322;
  wire while_asn_1324;
  wire while_asn_1326;
  wire while_asn_1328;
  wire while_asn_1330;
  wire while_asn_1332;
  wire while_asn_1334;
  wire while_asn_1336;
  wire while_asn_1338;
  wire while_asn_1340;
  wire while_asn_1342;
  wire while_asn_1344;
  wire while_asn_1346;
  wire while_asn_1348;
  wire while_asn_1350;
  wire while_asn_1352;
  wire while_asn_1354;
  wire while_asn_1356;
  wire while_asn_1358;
  wire while_asn_1360;
  wire [319:0] libraries_EAdd_0d1aed8b807329bc366abb192bb53bb66056_1;
  wire [319:0] libraries_EMul_50466378fb684d7351699b7bf1bdec8c6525_1;
  wire [319:0] libraries_Sigmoid_6ea22cc51ee279163d827d3cc5db43491cd81_1;
  wire [319:0] libraries_Tanh_0c47cc570305d1d8c1a9dd465101e61217b26_1;
  wire [319:0] libraries_Relu_29d7978308309996bcf6431af85e65007d30_1;
  wire [319:0] libraries_OneX_6a9c88d8c3af0ca712acdf3bbda5530a55e7_1;
  wire [319:0] libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1;
  reg [2:0] act_config_in_InstFetch_return_sva_4_2;
  wire mux_10_cse;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_cse;
  wire act_write_data_data_and_cse;
  wire ActUnit_PushAxiRsp_if_and_cse;
  wire ActUnit_PushAxiRsp_if_and_1_cse;
  wire mux_tmp_118;
  wire not_tmp_67;
  wire or_tmp_791;
  wire or_958_cse;
  wire or_957_cse;
  wire or_956_cse;
  wire or_955_cse;
  wire or_954_cse;
  wire or_953_cse;
  wire or_952_cse;
  wire or_951_cse;
  wire or_950_cse;
  wire or_949_cse;
  wire or_948_cse;
  wire or_947_cse;
  wire or_946_cse;
  wire or_945_cse;
  wire or_944_cse;
  wire or_943_cse;
  wire or_942_cse;
  wire or_941_cse;
  wire or_940_cse;
  wire or_939_cse;
  wire or_938_cse;
  wire or_937_cse;
  wire or_936_cse;
  wire or_935_cse;
  wire or_934_cse;
  wire or_933_cse;
  wire or_932_cse;
  wire or_931_cse;
  wire or_930_cse;
  wire or_929_cse;
  wire or_928_cse;
  wire or_925_cse;
  reg reg_act_regs_data_3_15_enexo;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo;
  reg reg_act_config_inst_counter_enexo;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_1;
  reg reg_act_regs_data_1_14_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_1;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_2;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_2;
  reg reg_act_regs_data_1_13_enexo;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_3;
  reg reg_act_regs_data_0_12_enexo;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_4;
  reg reg_act_regs_data_0_11_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_4;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_5;
  reg reg_act_regs_data_0_10_enexo;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_6;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_6;
  reg reg_act_regs_data_3_9_enexo;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_7;
  reg reg_act_regs_data_2_8_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_7;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_8;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_8;
  reg reg_act_regs_data_0_7_enexo;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_9;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_9;
  reg reg_act_regs_data_1_6_enexo;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_10;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_10;
  reg reg_act_regs_data_3_5_enexo;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_11;
  reg reg_act_regs_data_2_4_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_11;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_12;
  reg reg_act_regs_data_3_3_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_12;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_13;
  reg reg_act_regs_data_1_2_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_13;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_14;
  reg reg_act_regs_data_0_1_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_14;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_15;
  reg reg_act_regs_data_1_0_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_15;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_18_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_19_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_20_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_21_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_22_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_23_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_24_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_25_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_26_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_27_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_28_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_29_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_30_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_31_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_32_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_33_enex5;
  wire [19:0] nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [7:0] z_out_7_0;
  wire [8:0] nl_z_out_7_0;

  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_prb;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_prb;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb;
  wire[0:0] pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb;
  wire[0:0] pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb;
  wire[0:0] nor_12_nl;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1;
  wire[0:0] act_config_InstIncr_if_act_config_InstIncr_if_and_1_nl;
  wire[0:0] ActUnit_DecodeAxi_mux_88_nl;
  wire[0:0] ActUnit_DecodeAxi_if_mux_82_nl;
  wire[0:0] ActUnit_DecodeAxiWrite_mux_36_nl;
  wire[0:0] act_config_ActConfigWrite_mux_33_nl;
  wire[7:0] mux_91_nl;
  wire[0:0] and_1557_nl;
  wire[0:0] not_235_nl;
  wire[4:0] and_1554_nl;
  wire[4:0] while_while_while_or_nl;
  wire[0:0] while_while_not_nl;
  wire[0:0] mux_19_nl;
  wire[0:0] nand_6_nl;
  wire[0:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_2_nl;
  wire[0:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_33_nl;
  wire[0:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_5_nl;
  wire[0:0] mux_158_nl;
  wire[0:0] or_960_nl;
  wire[0:0] mux_157_nl;
  wire[0:0] mux_156_nl;
  wire[0:0] mux_155_nl;
  wire[0:0] mux_154_nl;
  wire[0:0] mux_153_nl;
  wire[0:0] mux_152_nl;
  wire[0:0] mux_151_nl;
  wire[0:0] mux_150_nl;
  wire[0:0] mux_149_nl;
  wire[0:0] and_1734_nl;
  wire[0:0] and_1733_nl;
  wire[0:0] mux_148_nl;
  wire[0:0] and_1732_nl;
  wire[0:0] and_1731_nl;
  wire[0:0] mux_147_nl;
  wire[0:0] mux_146_nl;
  wire[0:0] and_1730_nl;
  wire[0:0] and_1729_nl;
  wire[0:0] mux_145_nl;
  wire[0:0] and_1728_nl;
  wire[0:0] and_1727_nl;
  wire[0:0] mux_144_nl;
  wire[0:0] mux_143_nl;
  wire[0:0] mux_142_nl;
  wire[0:0] and_1726_nl;
  wire[0:0] and_1725_nl;
  wire[0:0] mux_141_nl;
  wire[0:0] and_1724_nl;
  wire[0:0] and_1723_nl;
  wire[0:0] mux_140_nl;
  wire[0:0] mux_139_nl;
  wire[0:0] and_1722_nl;
  wire[0:0] and_1721_nl;
  wire[0:0] mux_138_nl;
  wire[0:0] and_1720_nl;
  wire[0:0] and_1719_nl;
  wire[0:0] mux_137_nl;
  wire[0:0] mux_136_nl;
  wire[0:0] mux_135_nl;
  wire[0:0] mux_134_nl;
  wire[0:0] and_1718_nl;
  wire[0:0] and_1717_nl;
  wire[0:0] mux_133_nl;
  wire[0:0] and_1716_nl;
  wire[0:0] and_1715_nl;
  wire[0:0] mux_132_nl;
  wire[0:0] mux_131_nl;
  wire[0:0] and_1714_nl;
  wire[0:0] and_1713_nl;
  wire[0:0] mux_130_nl;
  wire[0:0] and_1712_nl;
  wire[0:0] and_1711_nl;
  wire[0:0] mux_129_nl;
  wire[0:0] mux_128_nl;
  wire[0:0] mux_127_nl;
  wire[0:0] and_1710_nl;
  wire[0:0] and_1709_nl;
  wire[0:0] mux_126_nl;
  wire[0:0] and_1708_nl;
  wire[0:0] and_1707_nl;
  wire[0:0] mux_125_nl;
  wire[0:0] mux_124_nl;
  wire[0:0] and_1706_nl;
  wire[0:0] and_1705_nl;
  wire[0:0] mux_123_nl;
  wire[0:0] and_1704_nl;
  wire[0:0] and_1703_nl;
  wire[0:0] nand_nl;
  wire[0:0] while_else_1_while_else_1_nand_nl;
  wire[0:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_31_nl;
  wire[0:0] mux_4_nl;
  wire[0:0] nor_16_nl;
  wire[0:0] or_1_nl;
  wire[4:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_21_nl;
  wire[0:0] ActUnit_DecodeAxiWrite_else_not_17_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_1_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_4_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_7_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_9_nl;
  wire[1:0] act_config_ActConfigWrite_if_mux_3_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_11_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_13_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_15_nl;
  wire[1:0] act_config_ActConfigWrite_if_mux_5_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_17_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_19_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_21_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_23_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_25_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_27_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_29_nl;
  wire[0:0] ActUnit_DecodeAxi_mux_89_nl;
  wire[0:0] ActUnit_DecodeAxi_if_mux_83_nl;
  wire[0:0] ActUnit_DecodeAxiWrite_mux_37_nl;
  wire[0:0] act_config_ActConfigWrite_mux_34_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_22_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_23_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_24_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_25_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_26_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_27_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_28_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_29_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_30_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_31_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_32_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_33_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_34_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_35_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_36_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_37_nl;
  wire[4:0] ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_and_1_nl;
  wire[0:0] mux_nl;
  wire[0:0] nor_14_nl;
  wire[0:0] mux_15_nl;
  wire[0:0] or_64_nl;
  wire[0:0] mux_121_nl;
  wire[0:0] mux_120_nl;
  wire[0:0] mux_119_nl;
  wire[0:0] mux_118_nl;
  wire[0:0] mux_117_nl;
  wire[0:0] mux_116_nl;
  wire[0:0] mux_115_nl;
  wire[0:0] mux_114_nl;
  wire[0:0] mux_113_nl;
  wire[0:0] mux_112_nl;
  wire[0:0] mux_111_nl;
  wire[0:0] mux_110_nl;
  wire[0:0] mux_109_nl;
  wire[0:0] mux_108_nl;
  wire[0:0] mux_107_nl;
  wire[0:0] mux_106_nl;
  wire[0:0] mux_105_nl;
  wire[0:0] mux_104_nl;
  wire[0:0] mux_103_nl;
  wire[0:0] mux_102_nl;
  wire[0:0] mux_101_nl;
  wire[0:0] mux_100_nl;
  wire[0:0] mux_99_nl;
  wire[0:0] mux_98_nl;
  wire[0:0] mux_97_nl;
  wire[0:0] mux_96_nl;
  wire[0:0] mux_95_nl;
  wire[0:0] mux_94_nl;
  wire[0:0] mux_93_nl;
  wire[0:0] mux_92_nl;
  wire[2:0] operator_8_false_operator_8_false_and_1_nl;
  wire[0:0] operator_8_false_nor_1_nl;
  wire[4:0] operator_8_false_operator_8_false_mux_2_nl;
  wire[4:0] operator_8_false_operator_8_false_mux_3_nl;

  // Interconnect Declarations for Component Instantiations 
  
  wire[7:0] ActUnit_PushAxiRsp_if_mux_10_nl;
  wire[7:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_47_nl;
  wire[7:0] act_config_ActConfigRead_else_else_mux_18_nl;
  wire[7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_40_nl;
  wire[7:0] ActUnit_PushAxiRsp_if_mux_9_nl;
  wire[7:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_45_nl;
  wire[7:0] act_config_ActConfigRead_else_else_mux_17_nl;
  wire[7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_39_nl;
  wire[7:0] ActUnit_PushAxiRsp_if_mux_8_nl;
  wire[7:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_43_nl;
  wire[7:0] act_config_ActConfigRead_else_else_mux_16_nl;
  wire[7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_38_nl;
  wire[7:0] ActUnit_PushAxiRsp_if_mux_7_nl;
  wire[7:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_41_nl;
  wire[7:0] act_config_ActConfigRead_else_else_mux_15_nl;
  wire[7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_37_nl;
  wire[7:0] ActUnit_PushAxiRsp_if_mux_6_nl;
  wire[7:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_39_nl;
  wire[7:0] act_config_ActConfigRead_else_else_mux_14_nl;
  wire[7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_36_nl;
  wire[7:0] ActUnit_PushAxiRsp_if_mux_5_nl;
  wire[7:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_37_nl;
  wire[7:0] act_config_ActConfigRead_else_else_mux_13_nl;
  wire[7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_35_nl;
  wire[7:0] ActUnit_PushAxiRsp_if_mux_4_nl;
  wire[7:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_35_nl;
  wire[7:0] act_config_ActConfigRead_else_else_mux_12_nl;
  wire[7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_34_nl;
  wire[7:0] and_1686_nl;
  wire[7:0] mux1h_65_nl;
  wire[0:0] not_366_nl;
  wire[7:0] ActUnit_PushAxiRsp_if_mux_2_nl;
  wire[7:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_33_nl;
  wire[7:0] act_config_ActConfigRead_else_else_mux_11_nl;
  wire[7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_33_nl;
  wire[2:0] act_mem_banks_read_read_data_mux_9_nl;
  wire[2:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_31_nl;
  wire[2:0] act_config_ActConfigRead_else_else_mux_10_nl;
  wire[2:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_32_nl;
  wire[4:0] and_1687_nl;
  wire[4:0] mux1h_66_nl;
  wire[0:0] not_370_nl;
  wire[7:0] ActUnit_PushAxiRsp_if_mux_1_nl;
  wire[7:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_29_nl;
  wire[7:0] act_config_ActConfigRead_else_else_mux_9_nl;
  wire[7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_31_nl;
  wire[7:0] and_1688_nl;
  wire[7:0] mux1h_67_nl;
  wire[0:0] not_374_nl;
  wire[1:0] act_mem_banks_read_read_data_mux_7_nl;
  wire[1:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_27_nl;
  wire[1:0] act_config_ActConfigRead_else_else_mux_8_nl;
  wire[1:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_30_nl;
  wire[5:0] and_1689_nl;
  wire[5:0] mux1h_68_nl;
  wire[0:0] act_mem_banks_read_read_data_and_19_nl;
  wire[0:0] act_mem_banks_read_read_data_and_20_nl;
  wire[0:0] act_mem_banks_read_read_data_and_21_nl;
  wire[0:0] not_378_nl;
  wire[4:0] act_mem_banks_read_read_data_mux_5_nl;
  wire[4:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_25_nl;
  wire[4:0] act_config_ActConfigRead_else_else_mux_7_nl;
  wire[4:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_29_nl;
  wire[2:0] and_1690_nl;
  wire[2:0] mux1h_69_nl;
  wire[0:0] not_382_nl;
  wire[6:0] act_mem_banks_read_read_data_mux_3_nl;
  wire[6:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_23_nl;
  wire[6:0] act_config_ActConfigRead_else_else_mux_6_nl;
  wire[6:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_28_nl;
  wire[0:0] act_mem_banks_read_read_data_mux_2_nl;
  wire[0:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_50_nl;
  wire[0:0] ActUnit_DecodeAxiRead_mux_27_nl;
  wire[0:0] act_config_ActConfigRead_else_mux_18_nl;
  wire[0:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_19_nl;
  wire[6:0] act_mem_banks_read_read_data_mux_1_nl;
  wire[6:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_21_nl;
  wire[6:0] act_config_ActConfigRead_else_else_mux_5_nl;
  wire[6:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_27_nl;
  wire[0:0] act_mem_banks_read_read_data_mux_nl;
  wire[0:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_49_nl;
  wire[0:0] ActUnit_DecodeAxiRead_mux_28_nl;
  wire[0:0] act_config_ActConfigRead_else_mux_20_nl;
  wire[0:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_21_nl;
  wire [127:0] nl_ActUnit_ActUnitRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun;

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit
// ------------------------------------------------------------------


module ActUnit (
  clk, rst, start_val, start_rdy, start_msg, act_port_val, act_port_rdy, act_port_msg,
      rva_in_val, rva_in_rdy, rva_in_msg, rva_out_val, rva_out_rdy, rva_out_msg,
      output_port_val, output_port_rdy, output_port_msg, done_val, done_rdy, done_msg
);
  input clk;
  input rst;
  input start_val;
  output start_rdy;
  input start_msg;
  input act_port_val;
  output act_port_rdy;
  input [319:0] act_port_msg;
  input rva_in_val;
  output rva_in_rdy;
  input [168:0] rva_in_msg;
  output rva_out_val;
  input rva_out_rdy;
  output [127:0] rva_out_msg;
  output output_port_val;
  input output_port_rdy;
  output [137:0] output_port_msg;
  output done_val;
  input done_rdy;
  output done_msg;

    // helpful signals for verification

    wire is_start = run.is_start_sva;
    wire state = is_start ? (run.fsm_output[1]? 3'b001:3'b010) : 3'b000;

    // Act_config
    wire act_config_is_valid = run.act_config_is_valid_sva;
    wire act_config_is_zero_first = run.act_config_is_zero_first_sva;
    wire [2:0] act_config_adpfloat_bias = run.act_config_adpfloat_bias_sva;
    wire [5:0] act_config_num_inst = run.act_config_num_inst_sva;
    wire [7:0] act_config_num_ouput = run.act_config_num_output_sva;
    wire [4:0] act_config_buffer_addr_base = run.act_config_buffer_addr_base_sva;
    wire [7:0] act_config_output_addr_base = run.act_config_output_addr_base_sva;
    wire [4:0] act_config_inst_counter = act_config_inst_counter_sva;
    wire [7:0] act_config_output_counter = act_config_output_counter_sva;



  // Interconnect Declarations for Component Instantiations 
  ActUnit_ActUnit_ActUnitRun run (
      .clk(clk),
      .rst(rst),
      .start_val(start_val),
      .start_rdy(start_rdy),
      .start_msg(start_msg),
      .act_port_val(act_port_val),
      .act_port_rdy(act_port_rdy),
      .act_port_msg(act_port_msg),
      .rva_in_val(rva_in_val),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_msg(rva_in_msg),
      .rva_out_val(rva_out_val),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_msg(rva_out_msg),
      .output_port_val(output_port_val),
      .output_port_rdy(output_port_rdy),
      .output_port_msg(output_port_msg),
      .done_val(done_val),
      .done_rdy(done_rdy),
      .done_msg(done_msg)
    );
endmodule



