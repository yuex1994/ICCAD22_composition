// ================================================================
// NVDLA Open Source Project
//
// Copyright(c) 2016 - 2017 NVIDIA Corporation. Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with
// this distribution for more information.
// ================================================================
// File Name: NV_NVDLA_SDP_CORE_x.v
module SDP_X_mgc_in_wire_wait_v1 (ld, vd, d, lz, vz, z);
  parameter integer rscid = 1;
  parameter integer width = 8;
  input ld;
  output vd;
  output [width-1:0] d;
  output lz;
  input vz;
  input [width-1:0] z;
  wire vd;
  wire [width-1:0] d;
  wire lz;
  assign d = z;
  assign lz = ld;
  assign vd = vz;
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/SDP_X_mgc_out_stdreg_wait_v1.v
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
// All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------
module SDP_X_mgc_out_stdreg_wait_v1 (ld, vd, d, lz, vz, z);
  parameter integer rscid = 1;
  parameter integer width = 8;
  input ld;
  output vd;
  input [width-1:0] d;
  output lz;
  input vz;
  output [width-1:0] z;
  wire vd;
  wire lz;
  wire [width-1:0] z;
  assign z = d;
  assign lz = ld;
  assign vd = vz;
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/SDP_X_mgc_io_sync_v1.v
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
// All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------
module SDP_X_mgc_io_sync_v1 (ld, lz);
    parameter valid = 0;
    input ld;
    output lz;
    wire lz;
    assign lz = ld;
endmodule
module SDP_X_mgc_in_sync_v1 (vd, vz);
    parameter valid = 1;
    output vd;
    input vz;
    wire vd;
    assign vd = vz;
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/SDP_X_mgc_in_wire_v1.v
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
// All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------
module SDP_X_mgc_in_wire_v1 (d, z);
  parameter integer rscid = 1;
  parameter integer width = 8;
  output [width-1:0] d;
  input [width-1:0] z;
  wire [width-1:0] d;
  assign d = z;
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/SDP_X_mgc_chan_in_v2.v
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
// All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------
module SDP_X_mgc_chan_in_v2 (ld, vd, d, lz, vz, z, sd, sld, sz, slz);
  parameter integer rscid = 1;
  parameter integer width = 8;
  parameter integer sz_width = 8;
  input ld;
  output vd;
  output [width-1:0] d;
  output lz;
  input vz;
  input [width-1:0] z;
  output [sz_width-1:0] sd;
  input sld;
  input [sz_width-1:0] sz;
  output slz;
  wire vd;
  wire [width-1:0] d;
  wire lz;
  assign d = z;
  assign lz = ld;
  assign vd = vz;
  assign sd = sz;
  assign slz = sld;
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_r_beh_v4.v
module SDP_X_mgc_shift_r_v4(a,s,z);
   parameter width_a = 4;
   parameter signd_a = 1;
   parameter width_s = 2;
   parameter width_z = 8;
   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;
   generate
     if (signd_a)
     begin: SIGNED
       assign z = fshr_u(a,s,a[width_a-1]);
     end
     else
     begin: UNSIGNED
       assign z = fshr_u(a,s,1'b0);
     end
   endgenerate
//Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u = result[olen-1:0];
      end
   endfunction // fshl_u
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v4.v
module SDP_X_mgc_shift_l_v4(a,s,z);
   parameter width_a = 4;
   parameter signd_a = 1;
   parameter width_s = 2;
   parameter width_z = 8;
   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;
   generate
   if (signd_a)
   begin: SIGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSIGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate
//Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 = result[olen-1:0];
      end
   endfunction // fshl_u
//Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u
endmodule
//------> ../td_ccore_solutions/leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_0/rtl.v
// ----------------------------------------------------------------------
// HLS HDL: Verilog Netlister
// HLS Version: 10.0/264918 Production Release
// HLS Date: Mon Aug 8 13:35:54 PDT 2016
//
// Generated by: ezhang@hk-sim-11-144
// Generated date: Sun Dec 11 15:25:45 2016
// ----------------------------------------------------------------------
//
// ------------------------------------------------------------------
// Design Unit: SDP_X_leading_sign_23_0
// ------------------------------------------------------------------
module SDP_X_leading_sign_23_0 (
  mantissa, rtn
);
  input [22:0] mantissa;
  output [4:0] rtn;
// Interconnect Declarations
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_10;
  wire[0:0] IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl;
  wire[0:0] IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl;
  wire[0:0] IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl;
  wire[0:0] IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl;
// Interconnect Declarations for Component Instantiations
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2 = ~((mantissa[20:19]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1 = ~((mantissa[22:21]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1 = ~((mantissa[18:17]!=2'b00));
  assign c_h_1_2 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1 & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3 = (mantissa[16:15]==2'b00)
      & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2 = ~((mantissa[12:11]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 = ~((mantissa[14:13]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1 = ~((mantissa[10:9]!=2'b00));
  assign c_h_1_5 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4 = (mantissa[8:7]==2'b00)
      & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1 & c_h_1_5;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2 = ~((mantissa[4:3]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 = ~((mantissa[6:5]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1 = ~((mantissa[2:1]!=2'b00));
  assign c_h_1_9 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2;
  assign c_h_1_10 = c_h_1_6 & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl = c_h_1_6 & (~ IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4);
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl = c_h_1_2 & (c_h_1_5 | (~
      IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3)) & (c_h_1_9 | (~ c_h_1_10));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1
      & (IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1 | (~ IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2))
      & (~((~(IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 & (IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1
      | (~ IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2)))) & c_h_1_6))
      & (~((~(IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 & (IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1
      | (~ IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2)))) & c_h_1_10));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl
      = ((~((mantissa[22]) | (~((mantissa[21:20]!=2'b01))))) & (~(((mantissa[18])
      | (~((mantissa[17:16]!=2'b01)))) & c_h_1_2)) & (~((~((~((mantissa[14]) | (~((mantissa[13:12]!=2'b01)))))
      & (~(((mantissa[10]) | (~((mantissa[9:8]!=2'b01)))) & c_h_1_5)))) & c_h_1_6))
      & (~((~((~((mantissa[6]) | (~((mantissa[5:4]!=2'b01))))) & (~((~((mantissa[2:1]==2'b01)))
      & c_h_1_9)))) & c_h_1_10))) | ((~ (mantissa[0])) & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1
      & c_h_1_9 & c_h_1_10);
  assign rtn = {c_h_1_10 , (IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl) , (IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl)
      , (IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl) , (IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl)};
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_bl_beh_v4.v
module SDP_X_mgc_shift_bl_v4(a,s,z);
   parameter width_a = 4;
   parameter signd_a = 1;
   parameter width_s = 2;
   parameter width_z = 8;
   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;
   generate if ( signd_a )
   begin: SIGNED
     assign z = fshl_s(a,s,a[width_a-1]);
   end
   else
   begin: UNSIGNED
     assign z = fshl_s(a,s,1'b0);
   end
   endgenerate
//Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 = result[olen-1:0];
      end
   endfunction // fshl_u
//Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u
//Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u = result[olen-1:0];
      end
   endfunction // fshl_u
//Shift left - signed shift argument
   function [width_z-1:0] fshl_s;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      reg [width_a:0] sbit_arg1;
      begin
// Ignoring the possibility that arg2[width_s-1] could be X
// because of customer complaints regarding X'es in simulation results
        if ( arg2[width_s-1] == 1'b0 )
        begin
          sbit_arg1[width_a:0] = {(width_a+1){1'b0}};
          fshl_s = fshl_u(arg1, arg2, sbit);
        end
        else
        begin
          sbit_arg1[width_a] = sbit;
          sbit_arg1[width_a-1:0] = arg1;
          fshl_s = fshr_u(sbit_arg1[width_a:1], ~arg2, sbit);
        end
      end
   endfunction
endmodule
//------> ../td_ccore_solutions/leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_0/rtl.v
// ----------------------------------------------------------------------
// HLS HDL: Verilog Netlister
// HLS Version: 10.0/264918 Production Release
// HLS Date: Mon Aug 8 13:35:54 PDT 2016
//
// Generated by: ezhang@hk-sim-10-065
// Generated date: Mon Jul 3 13:20:08 2017
// ----------------------------------------------------------------------
//
// ------------------------------------------------------------------
// Design Unit: SDP_X_leading_sign_49_0
// ------------------------------------------------------------------
module SDP_X_leading_sign_49_0 (
  mantissa, rtn
);
  input [48:0] mantissa;
  output [5:0] rtn;
// Interconnect Declarations
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_12;
  wire c_h_1_13;
  wire c_h_1_14;
  wire c_h_1_17;
  wire c_h_1_20;
  wire c_h_1_21;
  wire c_h_1_22;
  wire c_h_1_23;
  wire[0:0] IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl;
  wire[0:0] IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl;
  wire[0:0] IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl;
  wire[0:0] IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl;
  wire[0:0] IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl;
// Interconnect Declarations for Component Instantiations
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2 = ~((mantissa[46:45]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1 = ~((mantissa[48:47]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1 = ~((mantissa[44:43]!=2'b00));
  assign c_h_1_2 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3 = (mantissa[42:41]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2 = ~((mantissa[38:37]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 = ~((mantissa[40:39]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1 = ~((mantissa[36:35]!=2'b00));
  assign c_h_1_5 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4 = (mantissa[34:33]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1 & c_h_1_5;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2 = ~((mantissa[30:29]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 = ~((mantissa[32:31]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1 = ~((mantissa[28:27]!=2'b00));
  assign c_h_1_9 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3 = (mantissa[26:25]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2 = ~((mantissa[22:21]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1 = ~((mantissa[24:23]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1 = ~((mantissa[20:19]!=2'b00));
  assign c_h_1_12 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5 = (mantissa[18:17]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1 & c_h_1_12 & c_h_1_13;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2 = ~((mantissa[14:13]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1 = ~((mantissa[16:15]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1 = ~((mantissa[12:11]!=2'b00));
  assign c_h_1_17 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3 = (mantissa[10:9]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2 = ~((mantissa[6:5]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 = ~((mantissa[8:7]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1 = ~((mantissa[4:3]!=2'b00));
  assign c_h_1_20 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2;
  assign c_h_1_21 = c_h_1_17 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4 = (mantissa[2:1]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1 & c_h_1_20;
  assign c_h_1_22 = c_h_1_21 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4;
  assign c_h_1_23 = c_h_1_14 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl = c_h_1_14 & (c_h_1_22
      | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl = c_h_1_6 & (c_h_1_13 |
      (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4)) & (~((~(c_h_1_21
      & (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4))) & c_h_1_23));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl = c_h_1_2 & (c_h_1_5 |
      (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3)) & (~((~(c_h_1_9
      & (c_h_1_12 | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3))))
      & c_h_1_14)) & (~(((~(c_h_1_17 & (c_h_1_20 | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3))))
      | c_h_1_22) & c_h_1_23));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1
      & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1 | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2))
      & (~((~(IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1
      | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2)))) & c_h_1_6))
      & (~((~(IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1
      | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2)) & (~((~(IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1
      & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1 | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2))))
      & c_h_1_13)))) & c_h_1_14)) & (~(((~(IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1
      & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1 | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2))
      & (~((~(IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1
      | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2)))) & c_h_1_21))))
      | c_h_1_22) & c_h_1_23));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl
      = ((~((mantissa[48]) | (~((mantissa[47:46]!=2'b01))))) & (~(((mantissa[44])
      | (~((mantissa[43:42]!=2'b01)))) & c_h_1_2)) & (~((~((~((mantissa[40]) | (~((mantissa[39:38]!=2'b01)))))
      & (~(((mantissa[36]) | (~((mantissa[35:34]!=2'b01)))) & c_h_1_5)))) & c_h_1_6))
      & (~((~((~((mantissa[32]) | (~((mantissa[31:30]!=2'b01))))) & (~(((mantissa[28])
      | (~((mantissa[27:26]!=2'b01)))) & c_h_1_9)) & (~((~((~((mantissa[24]) | (~((mantissa[23:22]!=2'b01)))))
      & (~(((mantissa[20]) | (~((mantissa[19:18]!=2'b01)))) & c_h_1_12)))) & c_h_1_13))))
      & c_h_1_14)) & (~(((~((~((mantissa[16]) | (~((mantissa[15:14]!=2'b01))))) &
      (~(((mantissa[12]) | (~((mantissa[11:10]!=2'b01)))) & c_h_1_17)) & (~((~((~((mantissa[8])
      | (~((mantissa[7:6]!=2'b01))))) & (~(((mantissa[4]) | (~((mantissa[3:2]!=2'b01))))
      & c_h_1_20)))) & c_h_1_21)))) | c_h_1_22) & c_h_1_23))) | ((~ (mantissa[0]))
      & c_h_1_22 & c_h_1_23);
  assign rtn = {c_h_1_23 , (IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl) , (IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl)
      , (IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl) , (IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl)
      , (IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl)};
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_out_fifo_wait_core_v2001_v9.v
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
// All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------
module SDP_X_mgc_out_fifo_wait_core_v9 (clk, en, arst, srst, ld, vd, d, lz, vz, z, sd);
    parameter integer rscid = 0; // resource ID
    parameter integer width = 8; // fifo width
    parameter integer sz_width = 8; // size of port for elements in fifo
    parameter integer fifo_sz = 8; // fifo depth
    parameter integer ph_clk = 1; // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en = 1; // clock enable polarity
    parameter integer ph_arst = 1; // async reset polarity
    parameter integer ph_srst = 1; // sync reset polarity
    parameter integer ph_log2 = 3; // log2(fifo_sz)
   localparam integer fifo_b = width * fifo_sz;
    input clk;
    input en;
    input arst;
    input srst;
    input ld; // load data
    output vd; // fifo full active low
    input [width-1:0] d;
    output lz; // fifo ready to send
    input vz; // dest ready for data
    output [width-1:0] z;
    output [sz_width-1:0] sd;
    localparam integer fifo_mx = (fifo_sz > 0) ? (fifo_sz-1) : 0 ;
    localparam integer fifo_mx_over_8 = fifo_mx / 8 ;
    reg [fifo_mx:0] stat_pre;
    reg [fifo_mx:0] stat;
    reg [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff_pre;
    reg [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff;
    wire [fifo_mx:0] en_l;
    wire [fifo_mx_over_8:0] en_l_s;
    reg [width-1:0] buff_nxt;
    reg stat_nxt;
    reg stat_before;
    reg stat_after;
    reg [fifo_mx:0] en_l_var;
    integer i;
    genvar eni;
    wire [32:0] size_t;
    reg [31:0] count;
    reg [31:0] count_t;
    reg [32:0] n_elem;
// synopsys translate_off
    reg [31:0] peak = 32'b0;
// synopsys translate_on
    wire active;
    assign active = ld | vz; // (ld & ~vd) | (vz & ~lz);
    genvar igen;
    generate
    if ( fifo_sz > 0 )
    begin: FIFO_REG
      wire [31:0] delta;
// 0 : 32'b0 if ld==0 and (vz & stat[fifo_sz-1])==0
// or if ld==1 and (vz & stat[fifo_sz-1])==1
// +1 : 32'b1 if ld==1 and (vz & stat[fifo_sz-1])==0
// -1 : {32{1'b1}} if ld==0 and (vz & stat[fifo_sz-1])==1
      assign delta = {{31{(~ld & (vz & stat[fifo_sz-1]))}} , (vz & stat[fifo_sz-1]) ^ ld};
      assign vd = vz | ~stat[0];
      assign lz = ld | stat[fifo_sz-1];
      assign size_t = count + delta;
      assign sd = size_t[sz_width-1:0];
      assign z = (stat[fifo_sz-1]) ? buff[fifo_b-1:width*(fifo_sz-1)] : d;
      always @(*)
      begin: FIFOPROC
        n_elem = 33'b0;
        for (i = fifo_sz-1; i >= 0; i = i - 1)
        begin
          stat_before = (i != 0) ? stat[i-1] : 1'b0;
          stat_after = (i != (fifo_sz-1)) ? stat[i+1] : 1'b1;
          stat_nxt = stat_after &
                    (stat_before | (stat[i] & (~vz)) | (stat[i] & ld) | (ld & (~vz)));
          stat_pre[i] = stat_nxt;
          if (vz & stat_before )
            begin
              buff_nxt[0+:width] = buff[width*(i-1)+:width];
              en_l_var[i] = 1'b1;
            end
          else if (ld & ~((~vz) & stat[i]))
            begin
              buff_nxt = d;
              en_l_var[i] = 1'b1;
            end
          else
            begin
              buff_nxt = d; // Don't care input to disabled flop
              en_l_var[i] = 1'b0;
            end
          buff_pre[width*i+:width] = buff_nxt[0+:width];
          if ((stat_after == 1'b1) & (stat[i] == 1'b0))
            n_elem = ($unsigned(fifo_sz) - 1) - $unsigned(i);
        end
        if ( stat[fifo_sz-1] == 1'b0 )
          count_t = 32'b0;
        else if ( stat[0] == 1'b1 )
          count_t = fifo_sz;
        else
          count_t = n_elem[31:0];
        count = count_t;
// synopsys translate_off
        if ( peak < count )
          peak = count;
// synopsys translate_on
      end
      if (ph_en) begin: PH_EN_HI
        assign en_l_s[fifo_mx_over_8] = en & active;
        for (igen = 0 ; igen < fifo_sz ; igen = igen + 1) begin: NEED_A_LABEL
          assign en_l[igen] = en & en_l_var[igen];
        end
        for (igen = 1 ; igen <= fifo_mx_over_8 ; igen = igen + 1) begin: NEED_A_LABEL2
          assign en_l_s[igen-1] = en & (stat[igen*8]) & (active);
        end
      end
      else begin: PH_EN_LO
        assign en_l_s[fifo_mx_over_8] = en | ~active;
        for (igen = 0 ; igen < fifo_sz ; igen = igen + 1) begin: NEED_A_LABEL3
          assign en_l[igen] = en | ~en_l_var[igen];
        end
        for (igen = 1 ; igen <= fifo_mx_over_8 ; igen = igen + 1) begin: NEED_A_LABEL2
          assign en_l_s[igen-1] = en | (~stat[igen*8]) | (~active);
        end
      end
// Output registers:
      for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
      begin: BUF_GEN
        if (ph_clk==1) begin: POS_BUF
          if (ph_arst==0) begin: LABEL1
            always @(posedge clk or negedge arst)
            if (arst == 1'b0) begin
              stat[eni] <= 1'b0;
            end
            else if (srst == ph_srst) begin
              stat[eni] <= 1'b0;
            end
            else if (en_l_s[eni/8] == ph_en) begin
              stat[eni] <= stat_pre[eni];
            end
          end
          else begin: LABEL2 // ph_arst==1
            always @(posedge clk or posedge arst)
            if (arst == 1'b1) begin
              stat[eni] <= 1'b0;
            end
            else if (srst == ph_srst) begin
              stat[eni] <= 1'b0;
            end
            else if (en_l_s[eni/8] == ph_en) begin
              stat[eni] <= stat_pre[eni];
            end
          end
        end
        else begin: NEG_BUF
          if (ph_arst==0) begin: LABEL3
            always @(negedge clk or negedge arst)
            if (arst == 1'b0) begin
              stat[eni] <= 1'b0;
            end
            else if (srst == ph_srst) begin
              stat[eni] <= 1'b0;
            end
            else if (en_l_s[eni/8] == ph_en) begin
              stat[eni] <= stat_pre[eni];
            end
          end
          else begin: LABEL4 // ph_arst==1
            always @(negedge clk or posedge arst)
            if (arst == 1'b1) begin
              stat[eni] <= 1'b0;
            end
            else if (srst == ph_srst) begin
              stat[eni] <= 1'b0;
            end
            else if (en_l_s[eni/8] == ph_en) begin
              stat[eni] <= stat_pre[eni];
            end
          end
        end
      end
      for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
      begin: STATGEN2
        if (ph_clk==1) begin: POS_STAT
          if (ph_arst==0) begin: LABEL5
            always @(posedge clk or negedge arst)
            if (arst == 1'b0) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (srst == ph_srst) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (en_l[eni] == ph_en) begin
              buff[width*eni+:width] <= buff_pre[width*eni+:width];
            end
          end
          else begin: LABEL6 // ph_arst==1
            always @(posedge clk or posedge arst)
            if (arst == 1'b1) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (srst == ph_srst) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (en_l[eni] == ph_en) begin
              buff[width*eni+:width] <= buff_pre[width*eni+:width];
            end
          end
        end
        else begin: NEG_STAT // ph_clk==0
          if (ph_arst==0) begin: LABEL7
            always @(negedge clk or negedge arst)
            if (arst == 1'b0) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (srst == ph_srst) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (en_l[eni] == ph_en) begin
              buff[width*eni+:width] <= buff_pre[width*eni+:width];
            end
          end
          else begin: LABEL8 // ph_arst==1
            always @(negedge clk or posedge arst)
            if (arst == 1'b1) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (srst == ph_srst) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (en_l[eni] == ph_en) begin
              buff[width*eni+:width] <= buff_pre[width*eni+:width];
            end
          end
        end
      end
    end
    else
    begin: FEED_THRU
      assign vd = vz;
      assign lz = ld;
      assign z = d;
      assign sd = ld & ~vz;
    end
    endgenerate
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_pipe_v2001_v10.v
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
// All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------
/*
 *
 *             _______________________________________________
 * WRITER    |                                               |          READER
 *           |           MGC_PIPE                            |
 *           |           __________________________          |
 *        --<| vdout  --<| vd ---------------  vz<|-----ldin<|---
 *           |           |      FIFO              |          |
 *        ---|>ldout  ---|>ld ---------------- lz |> ---vdin |>--
 *        ---|>dout -----|>d  ---------------- dz |> ----din |>--
 *           |           |________________________|          |
 *           |_______________________________________________|
 *
 *    vdout - can be considered as a notFULL signal
 *    vdin  - can be considered as a notEMPTY signal
 *    write_stall - an internal debug signal formed from ldout & !vdout
 *    read_stall  - an internal debug signal formed from ldin & !vdin
 *
 */
// two clock pipe
module SDP_X_mgc_pipe_v10 (clk, en, arst, srst, ldin, vdin, din, ldout, vdout, dout, sd);
    parameter integer rscid = 0; // resource ID
    parameter integer width = 8; // fifo width
    parameter integer sz_width = 8; // width of size of elements in fifo
    parameter integer fifo_sz = 8; // fifo depth
    parameter integer log2_sz = 3; // log2(fifo_sz)
    parameter integer ph_clk = 1; // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en = 1; // clock enable polarity
    parameter integer ph_arst = 1; // async reset polarity
    parameter integer ph_srst = 1; // sync reset polarity
    input clk;
    input en;
    input arst;
    input srst;
    input ldin;
    output vdin;
    output [width-1:0] din;
    input ldout;
    output vdout;
    input [width-1:0] dout;
    output [sz_width-1:0] sd;
// synopsys translate_off
    wire write_stall;
    wire read_stall;
    assign write_stall = ldout & !vdout;
    assign read_stall = ldin & !vdin;
// synopsys translate_on
    SDP_X_mgc_out_fifo_wait_core_v9
    #(
        .rscid (rscid),
        .width (width),
        .sz_width (sz_width),
        .fifo_sz (fifo_sz),
        .ph_clk (ph_clk),
        .ph_en (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst),
        .ph_log2 (log2_sz)
    )
    FIFO
    (
        .clk (clk),
        .en (en),
        .arst (arst),
        .srst (srst),
        .ld (ldout),
        .vd (vdout),
        .d (dout),
        .lz (vdin),
        .vz (ldin),
        .z (din),
        .sd (sd)
    );
endmodule
//------> ./rtl.v
// ----------------------------------------------------------------------
// HLS HDL: Verilog Netlister
// HLS Version: 10.0/264918 Production Release
// HLS Date: Mon Aug 8 13:35:54 PDT 2016
//
// Generated by: ezhang@hk-sim-11-191
// Generated date: Thu Jul 6 11:21:49 2017
// ----------------------------------------------------------------------
//
// ------------------------------------------------------------------
// Design Unit: SDP_X_cfg_alu_shift_value_rsc_triosy_obj_unreg
// ------------------------------------------------------------------
module SDP_X_cfg_alu_shift_value_rsc_triosy_obj_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_cfg_alu_src_rsc_triosy_obj_unreg
// ------------------------------------------------------------------
module SDP_X_cfg_alu_src_rsc_triosy_obj_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_cfg_alu_algo_rsc_triosy_obj_unreg
// ------------------------------------------------------------------
module SDP_X_cfg_alu_algo_rsc_triosy_obj_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_cfg_alu_bypass_rsc_triosy_obj_unreg
// ------------------------------------------------------------------
module SDP_X_cfg_alu_bypass_rsc_triosy_obj_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_cfg_alu_op_rsc_triosy_obj_unreg
// ------------------------------------------------------------------
module SDP_X_cfg_alu_op_rsc_triosy_obj_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_chn_alu_out_rsci_unreg
// ------------------------------------------------------------------
module SDP_X_chn_alu_out_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_chn_alu_op_rsci_unreg
// ------------------------------------------------------------------
module SDP_X_chn_alu_op_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_chn_alu_in_rsci_unreg
// ------------------------------------------------------------------
module SDP_X_chn_alu_in_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_core_fsm
// FSM Module
// ------------------------------------------------------------------
module SDP_X_X_alu_core_core_fsm (
  nvdla_core_clk, nvdla_core_rstn, core_wen, fsm_output
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;
// FSM State Type Declaration for X_alu_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;
  reg [0:0] state_var;
  reg [0:0] state_var_NS;
// Interconnect Declarations for Component Instantiations
  always @(*)
  begin : X_alu_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
// core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_staller
// ------------------------------------------------------------------
module SDP_X_X_alu_core_staller (
  nvdla_core_clk, nvdla_core_rstn, core_wen, chn_alu_in_rsci_wen_comp, core_wten,
      chn_alu_op_rsci_wen_comp, chn_alu_out_rsci_wen_comp
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output core_wen;
  input chn_alu_in_rsci_wen_comp;
  output core_wten;
  reg core_wten;
  input chn_alu_op_rsci_wen_comp;
  input chn_alu_out_rsci_wen_comp;
// Interconnect Declarations for Component Instantiations
  assign core_wen = chn_alu_in_rsci_wen_comp & chn_alu_op_rsci_wen_comp & chn_alu_out_rsci_wen_comp;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_cfg_alu_shift_value_rsc_triosy_obj_cfg_alu_shift_value_rsc_triosy_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_alu_core_cfg_alu_shift_value_rsc_triosy_obj_cfg_alu_shift_value_rsc_triosy_wait_dp
    (
  nvdla_core_clk, nvdla_core_rstn, cfg_alu_shift_value_rsc_triosy_obj_bawt, cfg_alu_shift_value_rsc_triosy_obj_biwt,
      cfg_alu_shift_value_rsc_triosy_obj_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_alu_shift_value_rsc_triosy_obj_bawt;
  input cfg_alu_shift_value_rsc_triosy_obj_biwt;
  input cfg_alu_shift_value_rsc_triosy_obj_bdwt;
// Interconnect Declarations
  reg cfg_alu_shift_value_rsc_triosy_obj_bcwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_alu_shift_value_rsc_triosy_obj_bawt = cfg_alu_shift_value_rsc_triosy_obj_biwt
      | cfg_alu_shift_value_rsc_triosy_obj_bcwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_shift_value_rsc_triosy_obj_bcwt <= 1'b0;
    end
    else begin
      cfg_alu_shift_value_rsc_triosy_obj_bcwt <= ~((~(cfg_alu_shift_value_rsc_triosy_obj_bcwt
          | cfg_alu_shift_value_rsc_triosy_obj_biwt)) | cfg_alu_shift_value_rsc_triosy_obj_bdwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_cfg_alu_shift_value_rsc_triosy_obj_cfg_alu_shift_value_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_alu_core_cfg_alu_shift_value_rsc_triosy_obj_cfg_alu_shift_value_rsc_triosy_wait_ctrl
    (
  cfg_alu_shift_value_rsc_triosy_obj_oswt, core_wen, core_wten, cfg_alu_shift_value_rsc_triosy_obj_iswt0,
      cfg_alu_shift_value_rsc_triosy_obj_biwt, cfg_alu_shift_value_rsc_triosy_obj_bdwt
);
  input cfg_alu_shift_value_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_alu_shift_value_rsc_triosy_obj_iswt0;
  output cfg_alu_shift_value_rsc_triosy_obj_biwt;
  output cfg_alu_shift_value_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_alu_shift_value_rsc_triosy_obj_biwt = (~ core_wten) & cfg_alu_shift_value_rsc_triosy_obj_iswt0;
  assign cfg_alu_shift_value_rsc_triosy_obj_bdwt = cfg_alu_shift_value_rsc_triosy_obj_oswt
      & core_wen;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_cfg_alu_src_rsc_triosy_obj_cfg_alu_src_rsc_triosy_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_alu_core_cfg_alu_src_rsc_triosy_obj_cfg_alu_src_rsc_triosy_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, cfg_alu_src_rsc_triosy_obj_bawt, cfg_alu_src_rsc_triosy_obj_biwt,
      cfg_alu_src_rsc_triosy_obj_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_alu_src_rsc_triosy_obj_bawt;
  input cfg_alu_src_rsc_triosy_obj_biwt;
  input cfg_alu_src_rsc_triosy_obj_bdwt;
// Interconnect Declarations
  reg cfg_alu_src_rsc_triosy_obj_bcwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_alu_src_rsc_triosy_obj_bawt = cfg_alu_src_rsc_triosy_obj_biwt | cfg_alu_src_rsc_triosy_obj_bcwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_src_rsc_triosy_obj_bcwt <= 1'b0;
    end
    else begin
      cfg_alu_src_rsc_triosy_obj_bcwt <= ~((~(cfg_alu_src_rsc_triosy_obj_bcwt | cfg_alu_src_rsc_triosy_obj_biwt))
          | cfg_alu_src_rsc_triosy_obj_bdwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_cfg_alu_src_rsc_triosy_obj_cfg_alu_src_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_alu_core_cfg_alu_src_rsc_triosy_obj_cfg_alu_src_rsc_triosy_wait_ctrl (
  cfg_alu_src_rsc_triosy_obj_oswt, core_wen, core_wten, cfg_alu_src_rsc_triosy_obj_iswt0,
      cfg_alu_src_rsc_triosy_obj_biwt, cfg_alu_src_rsc_triosy_obj_bdwt
);
  input cfg_alu_src_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_alu_src_rsc_triosy_obj_iswt0;
  output cfg_alu_src_rsc_triosy_obj_biwt;
  output cfg_alu_src_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_alu_src_rsc_triosy_obj_biwt = (~ core_wten) & cfg_alu_src_rsc_triosy_obj_iswt0;
  assign cfg_alu_src_rsc_triosy_obj_bdwt = cfg_alu_src_rsc_triosy_obj_oswt & core_wen;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_cfg_alu_algo_rsc_triosy_obj_cfg_alu_algo_rsc_triosy_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_alu_core_cfg_alu_algo_rsc_triosy_obj_cfg_alu_algo_rsc_triosy_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, cfg_alu_algo_rsc_triosy_obj_bawt, cfg_alu_algo_rsc_triosy_obj_biwt,
      cfg_alu_algo_rsc_triosy_obj_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_alu_algo_rsc_triosy_obj_bawt;
  input cfg_alu_algo_rsc_triosy_obj_biwt;
  input cfg_alu_algo_rsc_triosy_obj_bdwt;
// Interconnect Declarations
  reg cfg_alu_algo_rsc_triosy_obj_bcwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_alu_algo_rsc_triosy_obj_bawt = cfg_alu_algo_rsc_triosy_obj_biwt | cfg_alu_algo_rsc_triosy_obj_bcwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_algo_rsc_triosy_obj_bcwt <= 1'b0;
    end
    else begin
      cfg_alu_algo_rsc_triosy_obj_bcwt <= ~((~(cfg_alu_algo_rsc_triosy_obj_bcwt |
          cfg_alu_algo_rsc_triosy_obj_biwt)) | cfg_alu_algo_rsc_triosy_obj_bdwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_cfg_alu_algo_rsc_triosy_obj_cfg_alu_algo_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_alu_core_cfg_alu_algo_rsc_triosy_obj_cfg_alu_algo_rsc_triosy_wait_ctrl (
  cfg_alu_algo_rsc_triosy_obj_oswt, core_wen, core_wten, cfg_alu_algo_rsc_triosy_obj_iswt0,
      cfg_alu_algo_rsc_triosy_obj_biwt, cfg_alu_algo_rsc_triosy_obj_bdwt
);
  input cfg_alu_algo_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_alu_algo_rsc_triosy_obj_iswt0;
  output cfg_alu_algo_rsc_triosy_obj_biwt;
  output cfg_alu_algo_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_alu_algo_rsc_triosy_obj_biwt = (~ core_wten) & cfg_alu_algo_rsc_triosy_obj_iswt0;
  assign cfg_alu_algo_rsc_triosy_obj_bdwt = cfg_alu_algo_rsc_triosy_obj_oswt & core_wen;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_cfg_alu_bypass_rsc_triosy_obj_cfg_alu_bypass_rsc_triosy_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_alu_core_cfg_alu_bypass_rsc_triosy_obj_cfg_alu_bypass_rsc_triosy_wait_dp
    (
  nvdla_core_clk, nvdla_core_rstn, cfg_alu_bypass_rsc_triosy_obj_bawt, cfg_alu_bypass_rsc_triosy_obj_biwt,
      cfg_alu_bypass_rsc_triosy_obj_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_alu_bypass_rsc_triosy_obj_bawt;
  input cfg_alu_bypass_rsc_triosy_obj_biwt;
  input cfg_alu_bypass_rsc_triosy_obj_bdwt;
// Interconnect Declarations
  reg cfg_alu_bypass_rsc_triosy_obj_bcwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_alu_bypass_rsc_triosy_obj_bawt = cfg_alu_bypass_rsc_triosy_obj_biwt
      | cfg_alu_bypass_rsc_triosy_obj_bcwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_bypass_rsc_triosy_obj_bcwt <= 1'b0;
    end
    else begin
      cfg_alu_bypass_rsc_triosy_obj_bcwt <= ~((~(cfg_alu_bypass_rsc_triosy_obj_bcwt
          | cfg_alu_bypass_rsc_triosy_obj_biwt)) | cfg_alu_bypass_rsc_triosy_obj_bdwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_cfg_alu_bypass_rsc_triosy_obj_cfg_alu_bypass_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_alu_core_cfg_alu_bypass_rsc_triosy_obj_cfg_alu_bypass_rsc_triosy_wait_ctrl
    (
  cfg_alu_bypass_rsc_triosy_obj_oswt, core_wen, core_wten, cfg_alu_bypass_rsc_triosy_obj_iswt0,
      cfg_alu_bypass_rsc_triosy_obj_biwt, cfg_alu_bypass_rsc_triosy_obj_bdwt
);
  input cfg_alu_bypass_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_alu_bypass_rsc_triosy_obj_iswt0;
  output cfg_alu_bypass_rsc_triosy_obj_biwt;
  output cfg_alu_bypass_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_alu_bypass_rsc_triosy_obj_biwt = (~ core_wten) & cfg_alu_bypass_rsc_triosy_obj_iswt0;
  assign cfg_alu_bypass_rsc_triosy_obj_bdwt = cfg_alu_bypass_rsc_triosy_obj_oswt
      & core_wen;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_cfg_alu_op_rsc_triosy_obj_cfg_alu_op_rsc_triosy_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_alu_core_cfg_alu_op_rsc_triosy_obj_cfg_alu_op_rsc_triosy_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, cfg_alu_op_rsc_triosy_obj_bawt, cfg_alu_op_rsc_triosy_obj_biwt,
      cfg_alu_op_rsc_triosy_obj_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_alu_op_rsc_triosy_obj_bawt;
  input cfg_alu_op_rsc_triosy_obj_biwt;
  input cfg_alu_op_rsc_triosy_obj_bdwt;
// Interconnect Declarations
  reg cfg_alu_op_rsc_triosy_obj_bcwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_alu_op_rsc_triosy_obj_bawt = cfg_alu_op_rsc_triosy_obj_biwt | cfg_alu_op_rsc_triosy_obj_bcwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_op_rsc_triosy_obj_bcwt <= 1'b0;
    end
    else begin
      cfg_alu_op_rsc_triosy_obj_bcwt <= ~((~(cfg_alu_op_rsc_triosy_obj_bcwt | cfg_alu_op_rsc_triosy_obj_biwt))
          | cfg_alu_op_rsc_triosy_obj_bdwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_cfg_alu_op_rsc_triosy_obj_cfg_alu_op_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_alu_core_cfg_alu_op_rsc_triosy_obj_cfg_alu_op_rsc_triosy_wait_ctrl (
  cfg_alu_op_rsc_triosy_obj_oswt, core_wen, core_wten, cfg_alu_op_rsc_triosy_obj_iswt0,
      cfg_alu_op_rsc_triosy_obj_biwt, cfg_alu_op_rsc_triosy_obj_bdwt
);
  input cfg_alu_op_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_alu_op_rsc_triosy_obj_iswt0;
  output cfg_alu_op_rsc_triosy_obj_biwt;
  output cfg_alu_op_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_alu_op_rsc_triosy_obj_biwt = (~ core_wten) & cfg_alu_op_rsc_triosy_obj_iswt0;
  assign cfg_alu_op_rsc_triosy_obj_bdwt = cfg_alu_op_rsc_triosy_obj_oswt & core_wen;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_chn_alu_out_rsci_chn_alu_out_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_alu_core_chn_alu_out_rsci_chn_alu_out_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_out_rsci_oswt, chn_alu_out_rsci_bawt,
      chn_alu_out_rsci_wen_comp, chn_alu_out_rsci_biwt, chn_alu_out_rsci_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_alu_out_rsci_oswt;
  output chn_alu_out_rsci_bawt;
  output chn_alu_out_rsci_wen_comp;
  input chn_alu_out_rsci_biwt;
  input chn_alu_out_rsci_bdwt;
// Interconnect Declarations
  reg chn_alu_out_rsci_bcwt;
// Interconnect Declarations for Component Instantiations
  assign chn_alu_out_rsci_bawt = chn_alu_out_rsci_biwt | chn_alu_out_rsci_bcwt;
  assign chn_alu_out_rsci_wen_comp = (~ chn_alu_out_rsci_oswt) | chn_alu_out_rsci_bawt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_bcwt <= 1'b0;
    end
    else begin
      chn_alu_out_rsci_bcwt <= ~((~(chn_alu_out_rsci_bcwt | chn_alu_out_rsci_biwt))
          | chn_alu_out_rsci_bdwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_chn_alu_out_rsci_chn_alu_out_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_alu_core_chn_alu_out_rsci_chn_alu_out_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_out_rsci_oswt, core_wen, core_wten, chn_alu_out_rsci_iswt0,
      chn_alu_out_rsci_ld_core_psct, chn_alu_out_rsci_biwt, chn_alu_out_rsci_bdwt,
      chn_alu_out_rsci_ld_core_sct, chn_alu_out_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_alu_out_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_alu_out_rsci_iswt0;
  input chn_alu_out_rsci_ld_core_psct;
  output chn_alu_out_rsci_biwt;
  output chn_alu_out_rsci_bdwt;
  output chn_alu_out_rsci_ld_core_sct;
  input chn_alu_out_rsci_vd;
// Interconnect Declarations
  wire chn_alu_out_rsci_ogwt;
  wire chn_alu_out_rsci_pdswt0;
  reg chn_alu_out_rsci_icwt;
// Interconnect Declarations for Component Instantiations
  assign chn_alu_out_rsci_pdswt0 = (~ core_wten) & chn_alu_out_rsci_iswt0;
  assign chn_alu_out_rsci_biwt = chn_alu_out_rsci_ogwt & chn_alu_out_rsci_vd;
  assign chn_alu_out_rsci_ogwt = chn_alu_out_rsci_pdswt0 | chn_alu_out_rsci_icwt;
  assign chn_alu_out_rsci_bdwt = chn_alu_out_rsci_oswt & core_wen;
  assign chn_alu_out_rsci_ld_core_sct = chn_alu_out_rsci_ld_core_psct & chn_alu_out_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_icwt <= 1'b0;
    end
    else begin
      chn_alu_out_rsci_icwt <= ~((~(chn_alu_out_rsci_icwt | chn_alu_out_rsci_pdswt0))
          | chn_alu_out_rsci_biwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_chn_alu_op_rsci_chn_alu_op_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_alu_core_chn_alu_op_rsci_chn_alu_op_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_op_rsci_oswt, chn_alu_op_rsci_bawt, chn_alu_op_rsci_wen_comp,
      chn_alu_op_rsci_d_mxwt, chn_alu_op_rsci_biwt, chn_alu_op_rsci_bdwt, chn_alu_op_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_alu_op_rsci_oswt;
  output chn_alu_op_rsci_bawt;
  output chn_alu_op_rsci_wen_comp;
  output [255:0] chn_alu_op_rsci_d_mxwt;
  input chn_alu_op_rsci_biwt;
  input chn_alu_op_rsci_bdwt;
  input [255:0] chn_alu_op_rsci_d;
// Interconnect Declarations
  reg chn_alu_op_rsci_bcwt;
  reg [255:0] chn_alu_op_rsci_d_bfwt;
// Interconnect Declarations for Component Instantiations
  assign chn_alu_op_rsci_bawt = chn_alu_op_rsci_biwt | chn_alu_op_rsci_bcwt;
  assign chn_alu_op_rsci_wen_comp = (~ chn_alu_op_rsci_oswt) | chn_alu_op_rsci_bawt;
  assign chn_alu_op_rsci_d_mxwt = MUX_v_256_2_2(chn_alu_op_rsci_d, chn_alu_op_rsci_d_bfwt,
      chn_alu_op_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_op_rsci_bcwt <= 1'b0;
      chn_alu_op_rsci_d_bfwt <= 256'b0;
    end
    else begin
      chn_alu_op_rsci_bcwt <= ~((~(chn_alu_op_rsci_bcwt | chn_alu_op_rsci_biwt))
          | chn_alu_op_rsci_bdwt);
      chn_alu_op_rsci_d_bfwt <= chn_alu_op_rsci_d_mxwt;
    end
  end
  function [255:0] MUX_v_256_2_2;
    input [255:0] input_0;
    input [255:0] input_1;
    input [0:0] sel;
    reg [255:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_256_2_2 = result;
  end
  endfunction
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_chn_alu_op_rsci_chn_alu_op_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_alu_core_chn_alu_op_rsci_chn_alu_op_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_op_rsci_oswt, core_wen, core_wten, chn_alu_op_rsci_iswt0,
      chn_alu_op_rsci_ld_core_psct, chn_alu_op_rsci_biwt, chn_alu_op_rsci_bdwt, chn_alu_op_rsci_ld_core_sct,
      chn_alu_op_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_alu_op_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_alu_op_rsci_iswt0;
  input chn_alu_op_rsci_ld_core_psct;
  output chn_alu_op_rsci_biwt;
  output chn_alu_op_rsci_bdwt;
  output chn_alu_op_rsci_ld_core_sct;
  input chn_alu_op_rsci_vd;
// Interconnect Declarations
  wire chn_alu_op_rsci_ogwt;
  wire chn_alu_op_rsci_pdswt0;
  reg chn_alu_op_rsci_icwt;
// Interconnect Declarations for Component Instantiations
  assign chn_alu_op_rsci_pdswt0 = (~ core_wten) & chn_alu_op_rsci_iswt0;
  assign chn_alu_op_rsci_biwt = chn_alu_op_rsci_ogwt & chn_alu_op_rsci_vd;
  assign chn_alu_op_rsci_ogwt = chn_alu_op_rsci_pdswt0 | chn_alu_op_rsci_icwt;
  assign chn_alu_op_rsci_bdwt = chn_alu_op_rsci_oswt & core_wen;
  assign chn_alu_op_rsci_ld_core_sct = chn_alu_op_rsci_ld_core_psct & chn_alu_op_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_op_rsci_icwt <= 1'b0;
    end
    else begin
      chn_alu_op_rsci_icwt <= ~((~(chn_alu_op_rsci_icwt | chn_alu_op_rsci_pdswt0))
          | chn_alu_op_rsci_biwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_chn_alu_in_rsci_chn_alu_in_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_alu_core_chn_alu_in_rsci_chn_alu_in_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_in_rsci_oswt, chn_alu_in_rsci_bawt, chn_alu_in_rsci_wen_comp,
      chn_alu_in_rsci_d_mxwt, chn_alu_in_rsci_biwt, chn_alu_in_rsci_bdwt, chn_alu_in_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_alu_in_rsci_oswt;
  output chn_alu_in_rsci_bawt;
  output chn_alu_in_rsci_wen_comp;
  output [511:0] chn_alu_in_rsci_d_mxwt;
  input chn_alu_in_rsci_biwt;
  input chn_alu_in_rsci_bdwt;
  input [511:0] chn_alu_in_rsci_d;
// Interconnect Declarations
  reg chn_alu_in_rsci_bcwt;
  reg [511:0] chn_alu_in_rsci_d_bfwt;
// Interconnect Declarations for Component Instantiations
  assign chn_alu_in_rsci_bawt = chn_alu_in_rsci_biwt | chn_alu_in_rsci_bcwt;
  assign chn_alu_in_rsci_wen_comp = (~ chn_alu_in_rsci_oswt) | chn_alu_in_rsci_bawt;
  assign chn_alu_in_rsci_d_mxwt = MUX_v_512_2_2(chn_alu_in_rsci_d, chn_alu_in_rsci_d_bfwt,
      chn_alu_in_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_in_rsci_bcwt <= 1'b0;
      chn_alu_in_rsci_d_bfwt <= 512'b0;
    end
    else begin
      chn_alu_in_rsci_bcwt <= ~((~(chn_alu_in_rsci_bcwt | chn_alu_in_rsci_biwt))
          | chn_alu_in_rsci_bdwt);
      chn_alu_in_rsci_d_bfwt <= chn_alu_in_rsci_d_mxwt;
    end
  end
  function [511:0] MUX_v_512_2_2;
    input [511:0] input_0;
    input [511:0] input_1;
    input [0:0] sel;
    reg [511:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_512_2_2 = result;
  end
  endfunction
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_chn_alu_in_rsci_chn_alu_in_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_alu_core_chn_alu_in_rsci_chn_alu_in_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_in_rsci_oswt, core_wen, chn_alu_in_rsci_iswt0,
      chn_alu_in_rsci_ld_core_psct, core_wten, chn_alu_in_rsci_biwt, chn_alu_in_rsci_bdwt,
      chn_alu_in_rsci_ld_core_sct, chn_alu_in_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_alu_in_rsci_oswt;
  input core_wen;
  input chn_alu_in_rsci_iswt0;
  input chn_alu_in_rsci_ld_core_psct;
  input core_wten;
  output chn_alu_in_rsci_biwt;
  output chn_alu_in_rsci_bdwt;
  output chn_alu_in_rsci_ld_core_sct;
  input chn_alu_in_rsci_vd;
// Interconnect Declarations
  wire chn_alu_in_rsci_ogwt;
  wire chn_alu_in_rsci_pdswt0;
  reg chn_alu_in_rsci_icwt;
// Interconnect Declarations for Component Instantiations
  assign chn_alu_in_rsci_pdswt0 = (~ core_wten) & chn_alu_in_rsci_iswt0;
  assign chn_alu_in_rsci_biwt = chn_alu_in_rsci_ogwt & chn_alu_in_rsci_vd;
  assign chn_alu_in_rsci_ogwt = chn_alu_in_rsci_pdswt0 | chn_alu_in_rsci_icwt;
  assign chn_alu_in_rsci_bdwt = chn_alu_in_rsci_oswt & core_wen;
  assign chn_alu_in_rsci_ld_core_sct = chn_alu_in_rsci_ld_core_psct & chn_alu_in_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_in_rsci_icwt <= 1'b0;
    end
    else begin
      chn_alu_in_rsci_icwt <= ~((~(chn_alu_in_rsci_icwt | chn_alu_in_rsci_pdswt0))
          | chn_alu_in_rsci_biwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_cfg_mul_src_rsc_triosy_obj_unreg
// ------------------------------------------------------------------
module SDP_X_cfg_mul_src_rsc_triosy_obj_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_cfg_mul_prelu_rsc_triosy_obj_unreg
// ------------------------------------------------------------------
module SDP_X_cfg_mul_prelu_rsc_triosy_obj_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_cfg_mul_bypass_rsc_triosy_obj_unreg
// ------------------------------------------------------------------
module SDP_X_cfg_mul_bypass_rsc_triosy_obj_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_cfg_mul_op_rsc_triosy_obj_unreg
// ------------------------------------------------------------------
module SDP_X_cfg_mul_op_rsc_triosy_obj_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_chn_mul_out_rsci_unreg
// ------------------------------------------------------------------
module SDP_X_chn_mul_out_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_chn_mul_op_rsci_unreg
// ------------------------------------------------------------------
module SDP_X_chn_mul_op_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_chn_mul_in_rsci_unreg
// ------------------------------------------------------------------
module SDP_X_chn_mul_in_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_core_fsm
// FSM Module
// ------------------------------------------------------------------
module SDP_X_X_mul_core_core_fsm (
  nvdla_core_clk, nvdla_core_rstn, core_wen, fsm_output
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;
// FSM State Type Declaration for X_mul_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;
  reg [0:0] state_var;
  reg [0:0] state_var_NS;
// Interconnect Declarations for Component Instantiations
  always @(*)
  begin : X_mul_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
// core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_staller
// ------------------------------------------------------------------
module SDP_X_X_mul_core_staller (
  nvdla_core_clk, nvdla_core_rstn, core_wen, chn_mul_in_rsci_wen_comp, core_wten,
      chn_mul_op_rsci_wen_comp, chn_mul_out_rsci_wen_comp
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output core_wen;
  input chn_mul_in_rsci_wen_comp;
  output core_wten;
  reg core_wten;
  input chn_mul_op_rsci_wen_comp;
  input chn_mul_out_rsci_wen_comp;
// Interconnect Declarations for Component Instantiations
  assign core_wen = chn_mul_in_rsci_wen_comp & chn_mul_op_rsci_wen_comp & chn_mul_out_rsci_wen_comp;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_cfg_mul_src_rsc_triosy_obj_cfg_mul_src_rsc_triosy_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_mul_core_cfg_mul_src_rsc_triosy_obj_cfg_mul_src_rsc_triosy_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, cfg_mul_src_rsc_triosy_obj_bawt, cfg_mul_src_rsc_triosy_obj_biwt,
      cfg_mul_src_rsc_triosy_obj_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_mul_src_rsc_triosy_obj_bawt;
  input cfg_mul_src_rsc_triosy_obj_biwt;
  input cfg_mul_src_rsc_triosy_obj_bdwt;
// Interconnect Declarations
  reg cfg_mul_src_rsc_triosy_obj_bcwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_mul_src_rsc_triosy_obj_bawt = cfg_mul_src_rsc_triosy_obj_biwt | cfg_mul_src_rsc_triosy_obj_bcwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_mul_src_rsc_triosy_obj_bcwt <= 1'b0;
    end
    else begin
      cfg_mul_src_rsc_triosy_obj_bcwt <= ~((~(cfg_mul_src_rsc_triosy_obj_bcwt | cfg_mul_src_rsc_triosy_obj_biwt))
          | cfg_mul_src_rsc_triosy_obj_bdwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_cfg_mul_src_rsc_triosy_obj_cfg_mul_src_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_mul_core_cfg_mul_src_rsc_triosy_obj_cfg_mul_src_rsc_triosy_wait_ctrl (
  cfg_mul_src_rsc_triosy_obj_oswt, core_wen, core_wten, cfg_mul_src_rsc_triosy_obj_iswt0,
      cfg_mul_src_rsc_triosy_obj_biwt, cfg_mul_src_rsc_triosy_obj_bdwt
);
  input cfg_mul_src_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_mul_src_rsc_triosy_obj_iswt0;
  output cfg_mul_src_rsc_triosy_obj_biwt;
  output cfg_mul_src_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_mul_src_rsc_triosy_obj_biwt = (~ core_wten) & cfg_mul_src_rsc_triosy_obj_iswt0;
  assign cfg_mul_src_rsc_triosy_obj_bdwt = cfg_mul_src_rsc_triosy_obj_oswt & core_wen;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_cfg_mul_prelu_rsc_triosy_obj_cfg_mul_prelu_rsc_triosy_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_mul_core_cfg_mul_prelu_rsc_triosy_obj_cfg_mul_prelu_rsc_triosy_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, cfg_mul_prelu_rsc_triosy_obj_bawt, cfg_mul_prelu_rsc_triosy_obj_biwt,
      cfg_mul_prelu_rsc_triosy_obj_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_mul_prelu_rsc_triosy_obj_bawt;
  input cfg_mul_prelu_rsc_triosy_obj_biwt;
  input cfg_mul_prelu_rsc_triosy_obj_bdwt;
// Interconnect Declarations
  reg cfg_mul_prelu_rsc_triosy_obj_bcwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_mul_prelu_rsc_triosy_obj_bawt = cfg_mul_prelu_rsc_triosy_obj_biwt |
      cfg_mul_prelu_rsc_triosy_obj_bcwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_mul_prelu_rsc_triosy_obj_bcwt <= 1'b0;
    end
    else begin
      cfg_mul_prelu_rsc_triosy_obj_bcwt <= ~((~(cfg_mul_prelu_rsc_triosy_obj_bcwt
          | cfg_mul_prelu_rsc_triosy_obj_biwt)) | cfg_mul_prelu_rsc_triosy_obj_bdwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_cfg_mul_prelu_rsc_triosy_obj_cfg_mul_prelu_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_mul_core_cfg_mul_prelu_rsc_triosy_obj_cfg_mul_prelu_rsc_triosy_wait_ctrl
    (
  cfg_mul_prelu_rsc_triosy_obj_oswt, core_wen, core_wten, cfg_mul_prelu_rsc_triosy_obj_iswt0,
      cfg_mul_prelu_rsc_triosy_obj_biwt, cfg_mul_prelu_rsc_triosy_obj_bdwt
);
  input cfg_mul_prelu_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_mul_prelu_rsc_triosy_obj_iswt0;
  output cfg_mul_prelu_rsc_triosy_obj_biwt;
  output cfg_mul_prelu_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_mul_prelu_rsc_triosy_obj_biwt = (~ core_wten) & cfg_mul_prelu_rsc_triosy_obj_iswt0;
  assign cfg_mul_prelu_rsc_triosy_obj_bdwt = cfg_mul_prelu_rsc_triosy_obj_oswt &
      core_wen;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_cfg_mul_bypass_rsc_triosy_obj_cfg_mul_bypass_rsc_triosy_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_mul_core_cfg_mul_bypass_rsc_triosy_obj_cfg_mul_bypass_rsc_triosy_wait_dp
    (
  nvdla_core_clk, nvdla_core_rstn, cfg_mul_bypass_rsc_triosy_obj_bawt, cfg_mul_bypass_rsc_triosy_obj_biwt,
      cfg_mul_bypass_rsc_triosy_obj_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_mul_bypass_rsc_triosy_obj_bawt;
  input cfg_mul_bypass_rsc_triosy_obj_biwt;
  input cfg_mul_bypass_rsc_triosy_obj_bdwt;
// Interconnect Declarations
  reg cfg_mul_bypass_rsc_triosy_obj_bcwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_mul_bypass_rsc_triosy_obj_bawt = cfg_mul_bypass_rsc_triosy_obj_biwt
      | cfg_mul_bypass_rsc_triosy_obj_bcwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_mul_bypass_rsc_triosy_obj_bcwt <= 1'b0;
    end
    else begin
      cfg_mul_bypass_rsc_triosy_obj_bcwt <= ~((~(cfg_mul_bypass_rsc_triosy_obj_bcwt
          | cfg_mul_bypass_rsc_triosy_obj_biwt)) | cfg_mul_bypass_rsc_triosy_obj_bdwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_cfg_mul_bypass_rsc_triosy_obj_cfg_mul_bypass_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_mul_core_cfg_mul_bypass_rsc_triosy_obj_cfg_mul_bypass_rsc_triosy_wait_ctrl
    (
  cfg_mul_bypass_rsc_triosy_obj_oswt, core_wen, core_wten, cfg_mul_bypass_rsc_triosy_obj_iswt0,
      cfg_mul_bypass_rsc_triosy_obj_biwt, cfg_mul_bypass_rsc_triosy_obj_bdwt
);
  input cfg_mul_bypass_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_mul_bypass_rsc_triosy_obj_iswt0;
  output cfg_mul_bypass_rsc_triosy_obj_biwt;
  output cfg_mul_bypass_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_mul_bypass_rsc_triosy_obj_biwt = (~ core_wten) & cfg_mul_bypass_rsc_triosy_obj_iswt0;
  assign cfg_mul_bypass_rsc_triosy_obj_bdwt = cfg_mul_bypass_rsc_triosy_obj_oswt
      & core_wen;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_cfg_mul_op_rsc_triosy_obj_cfg_mul_op_rsc_triosy_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_mul_core_cfg_mul_op_rsc_triosy_obj_cfg_mul_op_rsc_triosy_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, cfg_mul_op_rsc_triosy_obj_bawt, cfg_mul_op_rsc_triosy_obj_biwt,
      cfg_mul_op_rsc_triosy_obj_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_mul_op_rsc_triosy_obj_bawt;
  input cfg_mul_op_rsc_triosy_obj_biwt;
  input cfg_mul_op_rsc_triosy_obj_bdwt;
// Interconnect Declarations
  reg cfg_mul_op_rsc_triosy_obj_bcwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_mul_op_rsc_triosy_obj_bawt = cfg_mul_op_rsc_triosy_obj_biwt | cfg_mul_op_rsc_triosy_obj_bcwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_mul_op_rsc_triosy_obj_bcwt <= 1'b0;
    end
    else begin
      cfg_mul_op_rsc_triosy_obj_bcwt <= ~((~(cfg_mul_op_rsc_triosy_obj_bcwt | cfg_mul_op_rsc_triosy_obj_biwt))
          | cfg_mul_op_rsc_triosy_obj_bdwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_cfg_mul_op_rsc_triosy_obj_cfg_mul_op_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_mul_core_cfg_mul_op_rsc_triosy_obj_cfg_mul_op_rsc_triosy_wait_ctrl (
  cfg_mul_op_rsc_triosy_obj_oswt, core_wen, core_wten, cfg_mul_op_rsc_triosy_obj_iswt0,
      cfg_mul_op_rsc_triosy_obj_biwt, cfg_mul_op_rsc_triosy_obj_bdwt
);
  input cfg_mul_op_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_mul_op_rsc_triosy_obj_iswt0;
  output cfg_mul_op_rsc_triosy_obj_biwt;
  output cfg_mul_op_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_mul_op_rsc_triosy_obj_biwt = (~ core_wten) & cfg_mul_op_rsc_triosy_obj_iswt0;
  assign cfg_mul_op_rsc_triosy_obj_bdwt = cfg_mul_op_rsc_triosy_obj_oswt & core_wen;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_chn_mul_out_rsci_chn_mul_out_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_mul_core_chn_mul_out_rsci_chn_mul_out_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_out_rsci_oswt, chn_mul_out_rsci_bawt,
      chn_mul_out_rsci_wen_comp, chn_mul_out_rsci_biwt, chn_mul_out_rsci_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_mul_out_rsci_oswt;
  output chn_mul_out_rsci_bawt;
  output chn_mul_out_rsci_wen_comp;
  input chn_mul_out_rsci_biwt;
  input chn_mul_out_rsci_bdwt;
// Interconnect Declarations
  reg chn_mul_out_rsci_bcwt;
// Interconnect Declarations for Component Instantiations
  assign chn_mul_out_rsci_bawt = chn_mul_out_rsci_biwt | chn_mul_out_rsci_bcwt;
  assign chn_mul_out_rsci_wen_comp = (~ chn_mul_out_rsci_oswt) | chn_mul_out_rsci_bawt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_out_rsci_bcwt <= 1'b0;
    end
    else begin
      chn_mul_out_rsci_bcwt <= ~((~(chn_mul_out_rsci_bcwt | chn_mul_out_rsci_biwt))
          | chn_mul_out_rsci_bdwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_chn_mul_out_rsci_chn_mul_out_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_mul_core_chn_mul_out_rsci_chn_mul_out_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_out_rsci_oswt, core_wen, core_wten, chn_mul_out_rsci_iswt0,
      chn_mul_out_rsci_ld_core_psct, chn_mul_out_rsci_biwt, chn_mul_out_rsci_bdwt,
      chn_mul_out_rsci_ld_core_sct, chn_mul_out_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_mul_out_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_mul_out_rsci_iswt0;
  input chn_mul_out_rsci_ld_core_psct;
  output chn_mul_out_rsci_biwt;
  output chn_mul_out_rsci_bdwt;
  output chn_mul_out_rsci_ld_core_sct;
  input chn_mul_out_rsci_vd;
// Interconnect Declarations
  wire chn_mul_out_rsci_ogwt;
  wire chn_mul_out_rsci_pdswt0;
  reg chn_mul_out_rsci_icwt;
// Interconnect Declarations for Component Instantiations
  assign chn_mul_out_rsci_pdswt0 = (~ core_wten) & chn_mul_out_rsci_iswt0;
  assign chn_mul_out_rsci_biwt = chn_mul_out_rsci_ogwt & chn_mul_out_rsci_vd;
  assign chn_mul_out_rsci_ogwt = chn_mul_out_rsci_pdswt0 | chn_mul_out_rsci_icwt;
  assign chn_mul_out_rsci_bdwt = chn_mul_out_rsci_oswt & core_wen;
  assign chn_mul_out_rsci_ld_core_sct = chn_mul_out_rsci_ld_core_psct & chn_mul_out_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_out_rsci_icwt <= 1'b0;
    end
    else begin
      chn_mul_out_rsci_icwt <= ~((~(chn_mul_out_rsci_icwt | chn_mul_out_rsci_pdswt0))
          | chn_mul_out_rsci_biwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_chn_mul_op_rsci_chn_mul_op_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_mul_core_chn_mul_op_rsci_chn_mul_op_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_op_rsci_oswt, chn_mul_op_rsci_bawt, chn_mul_op_rsci_wen_comp,
      chn_mul_op_rsci_d_mxwt, chn_mul_op_rsci_biwt, chn_mul_op_rsci_bdwt, chn_mul_op_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_mul_op_rsci_oswt;
  output chn_mul_op_rsci_bawt;
  output chn_mul_op_rsci_wen_comp;
  output [255:0] chn_mul_op_rsci_d_mxwt;
  input chn_mul_op_rsci_biwt;
  input chn_mul_op_rsci_bdwt;
  input [255:0] chn_mul_op_rsci_d;
// Interconnect Declarations
  reg chn_mul_op_rsci_bcwt;
  reg [255:0] chn_mul_op_rsci_d_bfwt;
// Interconnect Declarations for Component Instantiations
  assign chn_mul_op_rsci_bawt = chn_mul_op_rsci_biwt | chn_mul_op_rsci_bcwt;
  assign chn_mul_op_rsci_wen_comp = (~ chn_mul_op_rsci_oswt) | chn_mul_op_rsci_bawt;
  assign chn_mul_op_rsci_d_mxwt = MUX_v_256_2_2(chn_mul_op_rsci_d, chn_mul_op_rsci_d_bfwt,
      chn_mul_op_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_op_rsci_bcwt <= 1'b0;
      chn_mul_op_rsci_d_bfwt <= 256'b0;
    end
    else begin
      chn_mul_op_rsci_bcwt <= ~((~(chn_mul_op_rsci_bcwt | chn_mul_op_rsci_biwt))
          | chn_mul_op_rsci_bdwt);
      chn_mul_op_rsci_d_bfwt <= chn_mul_op_rsci_d_mxwt;
    end
  end
  function [255:0] MUX_v_256_2_2;
    input [255:0] input_0;
    input [255:0] input_1;
    input [0:0] sel;
    reg [255:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_256_2_2 = result;
  end
  endfunction
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_chn_mul_op_rsci_chn_mul_op_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_mul_core_chn_mul_op_rsci_chn_mul_op_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_op_rsci_oswt, core_wen, core_wten, chn_mul_op_rsci_iswt0,
      chn_mul_op_rsci_ld_core_psct, chn_mul_op_rsci_biwt, chn_mul_op_rsci_bdwt, chn_mul_op_rsci_ld_core_sct,
      chn_mul_op_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_mul_op_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_mul_op_rsci_iswt0;
  input chn_mul_op_rsci_ld_core_psct;
  output chn_mul_op_rsci_biwt;
  output chn_mul_op_rsci_bdwt;
  output chn_mul_op_rsci_ld_core_sct;
  input chn_mul_op_rsci_vd;
// Interconnect Declarations
  wire chn_mul_op_rsci_ogwt;
  wire chn_mul_op_rsci_pdswt0;
  reg chn_mul_op_rsci_icwt;
// Interconnect Declarations for Component Instantiations
  assign chn_mul_op_rsci_pdswt0 = (~ core_wten) & chn_mul_op_rsci_iswt0;
  assign chn_mul_op_rsci_biwt = chn_mul_op_rsci_ogwt & chn_mul_op_rsci_vd;
  assign chn_mul_op_rsci_ogwt = chn_mul_op_rsci_pdswt0 | chn_mul_op_rsci_icwt;
  assign chn_mul_op_rsci_bdwt = chn_mul_op_rsci_oswt & core_wen;
  assign chn_mul_op_rsci_ld_core_sct = chn_mul_op_rsci_ld_core_psct & chn_mul_op_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_op_rsci_icwt <= 1'b0;
    end
    else begin
      chn_mul_op_rsci_icwt <= ~((~(chn_mul_op_rsci_icwt | chn_mul_op_rsci_pdswt0))
          | chn_mul_op_rsci_biwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_chn_mul_in_rsci_chn_mul_in_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_mul_core_chn_mul_in_rsci_chn_mul_in_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_in_rsci_oswt, chn_mul_in_rsci_bawt, chn_mul_in_rsci_wen_comp,
      chn_mul_in_rsci_d_mxwt, chn_mul_in_rsci_biwt, chn_mul_in_rsci_bdwt, chn_mul_in_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_mul_in_rsci_oswt;
  output chn_mul_in_rsci_bawt;
  output chn_mul_in_rsci_wen_comp;
  output [527:0] chn_mul_in_rsci_d_mxwt;
  input chn_mul_in_rsci_biwt;
  input chn_mul_in_rsci_bdwt;
  input [527:0] chn_mul_in_rsci_d;
// Interconnect Declarations
  reg chn_mul_in_rsci_bcwt;
  reg [527:0] chn_mul_in_rsci_d_bfwt;
// Interconnect Declarations for Component Instantiations
  assign chn_mul_in_rsci_bawt = chn_mul_in_rsci_biwt | chn_mul_in_rsci_bcwt;
  assign chn_mul_in_rsci_wen_comp = (~ chn_mul_in_rsci_oswt) | chn_mul_in_rsci_bawt;
  assign chn_mul_in_rsci_d_mxwt = MUX_v_528_2_2(chn_mul_in_rsci_d, chn_mul_in_rsci_d_bfwt,
      chn_mul_in_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_in_rsci_bcwt <= 1'b0;
      chn_mul_in_rsci_d_bfwt <= 528'b0;
    end
    else begin
      chn_mul_in_rsci_bcwt <= ~((~(chn_mul_in_rsci_bcwt | chn_mul_in_rsci_biwt))
          | chn_mul_in_rsci_bdwt);
      chn_mul_in_rsci_d_bfwt <= chn_mul_in_rsci_d_mxwt;
    end
  end
  function [527:0] MUX_v_528_2_2;
    input [527:0] input_0;
    input [527:0] input_1;
    input [0:0] sel;
    reg [527:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_528_2_2 = result;
  end
  endfunction
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_chn_mul_in_rsci_chn_mul_in_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_mul_core_chn_mul_in_rsci_chn_mul_in_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_in_rsci_oswt, core_wen, chn_mul_in_rsci_iswt0,
      chn_mul_in_rsci_ld_core_psct, core_wten, chn_mul_in_rsci_biwt, chn_mul_in_rsci_bdwt,
      chn_mul_in_rsci_ld_core_sct, chn_mul_in_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_mul_in_rsci_oswt;
  input core_wen;
  input chn_mul_in_rsci_iswt0;
  input chn_mul_in_rsci_ld_core_psct;
  input core_wten;
  output chn_mul_in_rsci_biwt;
  output chn_mul_in_rsci_bdwt;
  output chn_mul_in_rsci_ld_core_sct;
  input chn_mul_in_rsci_vd;
// Interconnect Declarations
  wire chn_mul_in_rsci_ogwt;
  wire chn_mul_in_rsci_pdswt0;
  reg chn_mul_in_rsci_icwt;
// Interconnect Declarations for Component Instantiations
  assign chn_mul_in_rsci_pdswt0 = (~ core_wten) & chn_mul_in_rsci_iswt0;
  assign chn_mul_in_rsci_biwt = chn_mul_in_rsci_ogwt & chn_mul_in_rsci_vd;
  assign chn_mul_in_rsci_ogwt = chn_mul_in_rsci_pdswt0 | chn_mul_in_rsci_icwt;
  assign chn_mul_in_rsci_bdwt = chn_mul_in_rsci_oswt & core_wen;
  assign chn_mul_in_rsci_ld_core_sct = chn_mul_in_rsci_ld_core_psct & chn_mul_in_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_in_rsci_icwt <= 1'b0;
    end
    else begin
      chn_mul_in_rsci_icwt <= ~((~(chn_mul_in_rsci_icwt | chn_mul_in_rsci_pdswt0))
          | chn_mul_in_rsci_biwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_cfg_mul_shift_value_rsc_triosy_obj_unreg
// ------------------------------------------------------------------
module SDP_X_cfg_mul_shift_value_rsc_triosy_obj_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_chn_trt_out_rsci_unreg
// ------------------------------------------------------------------
module SDP_X_chn_trt_out_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_chn_trt_in_rsci_unreg
// ------------------------------------------------------------------
module SDP_X_chn_trt_in_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_trt_core_core_fsm
// FSM Module
// ------------------------------------------------------------------
module SDP_X_X_trt_core_core_fsm (
  nvdla_core_clk, nvdla_core_rstn, core_wen, fsm_output
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;
// FSM State Type Declaration for X_trt_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;
  reg [0:0] state_var;
  reg [0:0] state_var_NS;
// Interconnect Declarations for Component Instantiations
  always @(*)
  begin : X_trt_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
// core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_trt_core_staller
// ------------------------------------------------------------------
module SDP_X_X_trt_core_staller (
  nvdla_core_clk, nvdla_core_rstn, core_wen, chn_trt_in_rsci_wen_comp, core_wten,
      chn_trt_out_rsci_wen_comp
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output core_wen;
  input chn_trt_in_rsci_wen_comp;
  output core_wten;
  reg core_wten;
  input chn_trt_out_rsci_wen_comp;
// Interconnect Declarations for Component Instantiations
  assign core_wen = chn_trt_in_rsci_wen_comp & chn_trt_out_rsci_wen_comp;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_trt_core_cfg_mul_shift_value_rsc_triosy_obj_cfg_mul_shift_value_rsc_triosy_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_trt_core_cfg_mul_shift_value_rsc_triosy_obj_cfg_mul_shift_value_rsc_triosy_wait_dp
    (
  nvdla_core_clk, nvdla_core_rstn, cfg_mul_shift_value_rsc_triosy_obj_bawt, cfg_mul_shift_value_rsc_triosy_obj_biwt,
      cfg_mul_shift_value_rsc_triosy_obj_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_mul_shift_value_rsc_triosy_obj_bawt;
  input cfg_mul_shift_value_rsc_triosy_obj_biwt;
  input cfg_mul_shift_value_rsc_triosy_obj_bdwt;
// Interconnect Declarations
  reg cfg_mul_shift_value_rsc_triosy_obj_bcwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_mul_shift_value_rsc_triosy_obj_bawt = cfg_mul_shift_value_rsc_triosy_obj_biwt
      | cfg_mul_shift_value_rsc_triosy_obj_bcwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_mul_shift_value_rsc_triosy_obj_bcwt <= 1'b0;
    end
    else begin
      cfg_mul_shift_value_rsc_triosy_obj_bcwt <= ~((~(cfg_mul_shift_value_rsc_triosy_obj_bcwt
          | cfg_mul_shift_value_rsc_triosy_obj_biwt)) | cfg_mul_shift_value_rsc_triosy_obj_bdwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_trt_core_cfg_mul_shift_value_rsc_triosy_obj_cfg_mul_shift_value_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_trt_core_cfg_mul_shift_value_rsc_triosy_obj_cfg_mul_shift_value_rsc_triosy_wait_ctrl
    (
  cfg_mul_shift_value_rsc_triosy_obj_oswt, core_wen, core_wten, cfg_mul_shift_value_rsc_triosy_obj_iswt0,
      cfg_mul_shift_value_rsc_triosy_obj_biwt, cfg_mul_shift_value_rsc_triosy_obj_bdwt
);
  input cfg_mul_shift_value_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_mul_shift_value_rsc_triosy_obj_iswt0;
  output cfg_mul_shift_value_rsc_triosy_obj_biwt;
  output cfg_mul_shift_value_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_mul_shift_value_rsc_triosy_obj_biwt = (~ core_wten) & cfg_mul_shift_value_rsc_triosy_obj_iswt0;
  assign cfg_mul_shift_value_rsc_triosy_obj_bdwt = cfg_mul_shift_value_rsc_triosy_obj_oswt
      & core_wen;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_trt_core_chn_trt_out_rsci_chn_trt_out_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_trt_core_chn_trt_out_rsci_chn_trt_out_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_trt_out_rsci_oswt, chn_trt_out_rsci_bawt,
      chn_trt_out_rsci_wen_comp, chn_trt_out_rsci_biwt, chn_trt_out_rsci_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_trt_out_rsci_oswt;
  output chn_trt_out_rsci_bawt;
  output chn_trt_out_rsci_wen_comp;
  input chn_trt_out_rsci_biwt;
  input chn_trt_out_rsci_bdwt;
// Interconnect Declarations
  reg chn_trt_out_rsci_bcwt;
// Interconnect Declarations for Component Instantiations
  assign chn_trt_out_rsci_bawt = chn_trt_out_rsci_biwt | chn_trt_out_rsci_bcwt;
  assign chn_trt_out_rsci_wen_comp = (~ chn_trt_out_rsci_oswt) | chn_trt_out_rsci_bawt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_out_rsci_bcwt <= 1'b0;
    end
    else begin
      chn_trt_out_rsci_bcwt <= ~((~(chn_trt_out_rsci_bcwt | chn_trt_out_rsci_biwt))
          | chn_trt_out_rsci_bdwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_trt_core_chn_trt_out_rsci_chn_trt_out_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_trt_core_chn_trt_out_rsci_chn_trt_out_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_trt_out_rsci_oswt, core_wen, core_wten, chn_trt_out_rsci_iswt0,
      chn_trt_out_rsci_ld_core_psct, chn_trt_out_rsci_biwt, chn_trt_out_rsci_bdwt,
      chn_trt_out_rsci_ld_core_sct, chn_trt_out_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_trt_out_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_trt_out_rsci_iswt0;
  input chn_trt_out_rsci_ld_core_psct;
  output chn_trt_out_rsci_biwt;
  output chn_trt_out_rsci_bdwt;
  output chn_trt_out_rsci_ld_core_sct;
  input chn_trt_out_rsci_vd;
// Interconnect Declarations
  wire chn_trt_out_rsci_ogwt;
  wire chn_trt_out_rsci_pdswt0;
  reg chn_trt_out_rsci_icwt;
// Interconnect Declarations for Component Instantiations
  assign chn_trt_out_rsci_pdswt0 = (~ core_wten) & chn_trt_out_rsci_iswt0;
  assign chn_trt_out_rsci_biwt = chn_trt_out_rsci_ogwt & chn_trt_out_rsci_vd;
  assign chn_trt_out_rsci_ogwt = chn_trt_out_rsci_pdswt0 | chn_trt_out_rsci_icwt;
  assign chn_trt_out_rsci_bdwt = chn_trt_out_rsci_oswt & core_wen;
  assign chn_trt_out_rsci_ld_core_sct = chn_trt_out_rsci_ld_core_psct & chn_trt_out_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_out_rsci_icwt <= 1'b0;
    end
    else begin
      chn_trt_out_rsci_icwt <= ~((~(chn_trt_out_rsci_icwt | chn_trt_out_rsci_pdswt0))
          | chn_trt_out_rsci_biwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_trt_core_chn_trt_in_rsci_chn_trt_in_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_trt_core_chn_trt_in_rsci_chn_trt_in_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_trt_in_rsci_oswt, chn_trt_in_rsci_bawt, chn_trt_in_rsci_wen_comp,
      chn_trt_in_rsci_d_mxwt, chn_trt_in_rsci_biwt, chn_trt_in_rsci_bdwt, chn_trt_in_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_trt_in_rsci_oswt;
  output chn_trt_in_rsci_bawt;
  output chn_trt_in_rsci_wen_comp;
  output [799:0] chn_trt_in_rsci_d_mxwt;
  input chn_trt_in_rsci_biwt;
  input chn_trt_in_rsci_bdwt;
  input [799:0] chn_trt_in_rsci_d;
// Interconnect Declarations
  reg chn_trt_in_rsci_bcwt;
  reg [799:0] chn_trt_in_rsci_d_bfwt;
// Interconnect Declarations for Component Instantiations
  assign chn_trt_in_rsci_bawt = chn_trt_in_rsci_biwt | chn_trt_in_rsci_bcwt;
  assign chn_trt_in_rsci_wen_comp = (~ chn_trt_in_rsci_oswt) | chn_trt_in_rsci_bawt;
  assign chn_trt_in_rsci_d_mxwt = MUX_v_800_2_2(chn_trt_in_rsci_d, chn_trt_in_rsci_d_bfwt,
      chn_trt_in_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_in_rsci_bcwt <= 1'b0;
      chn_trt_in_rsci_d_bfwt <= 800'b0;
    end
    else begin
      chn_trt_in_rsci_bcwt <= ~((~(chn_trt_in_rsci_bcwt | chn_trt_in_rsci_biwt))
          | chn_trt_in_rsci_bdwt);
      chn_trt_in_rsci_d_bfwt <= chn_trt_in_rsci_d_mxwt;
    end
  end
  function [799:0] MUX_v_800_2_2;
    input [799:0] input_0;
    input [799:0] input_1;
    input [0:0] sel;
    reg [799:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_800_2_2 = result;
  end
  endfunction
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_trt_core_chn_trt_in_rsci_chn_trt_in_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_trt_core_chn_trt_in_rsci_chn_trt_in_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_trt_in_rsci_oswt, core_wen, chn_trt_in_rsci_iswt0,
      chn_trt_in_rsci_ld_core_psct, core_wten, chn_trt_in_rsci_biwt, chn_trt_in_rsci_bdwt,
      chn_trt_in_rsci_ld_core_sct, chn_trt_in_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_trt_in_rsci_oswt;
  input core_wen;
  input chn_trt_in_rsci_iswt0;
  input chn_trt_in_rsci_ld_core_psct;
  input core_wten;
  output chn_trt_in_rsci_biwt;
  output chn_trt_in_rsci_bdwt;
  output chn_trt_in_rsci_ld_core_sct;
  input chn_trt_in_rsci_vd;
// Interconnect Declarations
  wire chn_trt_in_rsci_ogwt;
  wire chn_trt_in_rsci_pdswt0;
  reg chn_trt_in_rsci_icwt;
// Interconnect Declarations for Component Instantiations
  assign chn_trt_in_rsci_pdswt0 = (~ core_wten) & chn_trt_in_rsci_iswt0;
  assign chn_trt_in_rsci_biwt = chn_trt_in_rsci_ogwt & chn_trt_in_rsci_vd;
  assign chn_trt_in_rsci_ogwt = chn_trt_in_rsci_pdswt0 | chn_trt_in_rsci_icwt;
  assign chn_trt_in_rsci_bdwt = chn_trt_in_rsci_oswt & core_wen;
  assign chn_trt_in_rsci_ld_core_sct = chn_trt_in_rsci_ld_core_psct & chn_trt_in_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_in_rsci_icwt <= 1'b0;
    end
    else begin
      chn_trt_in_rsci_icwt <= ~((~(chn_trt_in_rsci_icwt | chn_trt_in_rsci_pdswt0))
          | chn_trt_in_rsci_biwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_cfg_relu_bypass_rsc_triosy_obj_unreg
// ------------------------------------------------------------------
module SDP_X_cfg_relu_bypass_rsc_triosy_obj_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_chn_relu_out_rsci_unreg
// ------------------------------------------------------------------
module SDP_X_chn_relu_out_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_chn_relu_in_rsci_unreg
// ------------------------------------------------------------------
module SDP_X_chn_relu_in_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_relu_core_core_fsm
// FSM Module
// ------------------------------------------------------------------
module SDP_X_X_relu_core_core_fsm (
  nvdla_core_clk, nvdla_core_rstn, core_wen, fsm_output
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;
// FSM State Type Declaration for X_relu_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;
  reg [0:0] state_var;
  reg [0:0] state_var_NS;
// Interconnect Declarations for Component Instantiations
  always @(*)
  begin : X_relu_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
// core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_relu_core_staller
// ------------------------------------------------------------------
module SDP_X_X_relu_core_staller (
  nvdla_core_clk, nvdla_core_rstn, core_wen, chn_relu_in_rsci_wen_comp, core_wten,
      chn_relu_out_rsci_wen_comp
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output core_wen;
  input chn_relu_in_rsci_wen_comp;
  output core_wten;
  reg core_wten;
  input chn_relu_out_rsci_wen_comp;
// Interconnect Declarations for Component Instantiations
  assign core_wen = chn_relu_in_rsci_wen_comp & chn_relu_out_rsci_wen_comp;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_relu_core_cfg_relu_bypass_rsc_triosy_obj_cfg_relu_bypass_rsc_triosy_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_relu_core_cfg_relu_bypass_rsc_triosy_obj_cfg_relu_bypass_rsc_triosy_wait_dp
    (
  nvdla_core_clk, nvdla_core_rstn, cfg_relu_bypass_rsc_triosy_obj_bawt, cfg_relu_bypass_rsc_triosy_obj_biwt,
      cfg_relu_bypass_rsc_triosy_obj_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_relu_bypass_rsc_triosy_obj_bawt;
  input cfg_relu_bypass_rsc_triosy_obj_biwt;
  input cfg_relu_bypass_rsc_triosy_obj_bdwt;
// Interconnect Declarations
  reg cfg_relu_bypass_rsc_triosy_obj_bcwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_relu_bypass_rsc_triosy_obj_bawt = cfg_relu_bypass_rsc_triosy_obj_biwt
      | cfg_relu_bypass_rsc_triosy_obj_bcwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_relu_bypass_rsc_triosy_obj_bcwt <= 1'b0;
    end
    else begin
      cfg_relu_bypass_rsc_triosy_obj_bcwt <= ~((~(cfg_relu_bypass_rsc_triosy_obj_bcwt
          | cfg_relu_bypass_rsc_triosy_obj_biwt)) | cfg_relu_bypass_rsc_triosy_obj_bdwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_relu_core_cfg_relu_bypass_rsc_triosy_obj_cfg_relu_bypass_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_relu_core_cfg_relu_bypass_rsc_triosy_obj_cfg_relu_bypass_rsc_triosy_wait_ctrl
    (
  cfg_relu_bypass_rsc_triosy_obj_oswt, core_wen, core_wten, cfg_relu_bypass_rsc_triosy_obj_iswt0,
      cfg_relu_bypass_rsc_triosy_obj_biwt, cfg_relu_bypass_rsc_triosy_obj_bdwt
);
  input cfg_relu_bypass_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_relu_bypass_rsc_triosy_obj_iswt0;
  output cfg_relu_bypass_rsc_triosy_obj_biwt;
  output cfg_relu_bypass_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  assign cfg_relu_bypass_rsc_triosy_obj_biwt = (~ core_wten) & cfg_relu_bypass_rsc_triosy_obj_iswt0;
  assign cfg_relu_bypass_rsc_triosy_obj_bdwt = cfg_relu_bypass_rsc_triosy_obj_oswt
      & core_wen;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_relu_core_chn_relu_out_rsci_chn_relu_out_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_relu_core_chn_relu_out_rsci_chn_relu_out_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_relu_out_rsci_oswt, chn_relu_out_rsci_bawt,
      chn_relu_out_rsci_wen_comp, chn_relu_out_rsci_biwt, chn_relu_out_rsci_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_relu_out_rsci_oswt;
  output chn_relu_out_rsci_bawt;
  output chn_relu_out_rsci_wen_comp;
  input chn_relu_out_rsci_biwt;
  input chn_relu_out_rsci_bdwt;
// Interconnect Declarations
  reg chn_relu_out_rsci_bcwt;
// Interconnect Declarations for Component Instantiations
  assign chn_relu_out_rsci_bawt = chn_relu_out_rsci_biwt | chn_relu_out_rsci_bcwt;
  assign chn_relu_out_rsci_wen_comp = (~ chn_relu_out_rsci_oswt) | chn_relu_out_rsci_bawt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_relu_out_rsci_bcwt <= 1'b0;
    end
    else begin
      chn_relu_out_rsci_bcwt <= ~((~(chn_relu_out_rsci_bcwt | chn_relu_out_rsci_biwt))
          | chn_relu_out_rsci_bdwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_relu_core_chn_relu_out_rsci_chn_relu_out_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_relu_core_chn_relu_out_rsci_chn_relu_out_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_relu_out_rsci_oswt, core_wen, core_wten, chn_relu_out_rsci_iswt0,
      chn_relu_out_rsci_ld_core_psct, chn_relu_out_rsci_biwt, chn_relu_out_rsci_bdwt,
      chn_relu_out_rsci_ld_core_sct, chn_relu_out_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_relu_out_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_relu_out_rsci_iswt0;
  input chn_relu_out_rsci_ld_core_psct;
  output chn_relu_out_rsci_biwt;
  output chn_relu_out_rsci_bdwt;
  output chn_relu_out_rsci_ld_core_sct;
  input chn_relu_out_rsci_vd;
// Interconnect Declarations
  wire chn_relu_out_rsci_ogwt;
  wire chn_relu_out_rsci_pdswt0;
  reg chn_relu_out_rsci_icwt;
// Interconnect Declarations for Component Instantiations
  assign chn_relu_out_rsci_pdswt0 = (~ core_wten) & chn_relu_out_rsci_iswt0;
  assign chn_relu_out_rsci_biwt = chn_relu_out_rsci_ogwt & chn_relu_out_rsci_vd;
  assign chn_relu_out_rsci_ogwt = chn_relu_out_rsci_pdswt0 | chn_relu_out_rsci_icwt;
  assign chn_relu_out_rsci_bdwt = chn_relu_out_rsci_oswt & core_wen;
  assign chn_relu_out_rsci_ld_core_sct = chn_relu_out_rsci_ld_core_psct & chn_relu_out_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_relu_out_rsci_icwt <= 1'b0;
    end
    else begin
      chn_relu_out_rsci_icwt <= ~((~(chn_relu_out_rsci_icwt | chn_relu_out_rsci_pdswt0))
          | chn_relu_out_rsci_biwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_relu_core_chn_relu_in_rsci_chn_relu_in_wait_dp
// ------------------------------------------------------------------
module SDP_X_X_relu_core_chn_relu_in_rsci_chn_relu_in_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_relu_in_rsci_oswt, chn_relu_in_rsci_bawt,
      chn_relu_in_rsci_wen_comp, chn_relu_in_rsci_d_mxwt, chn_relu_in_rsci_biwt,
      chn_relu_in_rsci_bdwt, chn_relu_in_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_relu_in_rsci_oswt;
  output chn_relu_in_rsci_bawt;
  output chn_relu_in_rsci_wen_comp;
  output [511:0] chn_relu_in_rsci_d_mxwt;
  input chn_relu_in_rsci_biwt;
  input chn_relu_in_rsci_bdwt;
  input [511:0] chn_relu_in_rsci_d;
// Interconnect Declarations
  reg chn_relu_in_rsci_bcwt;
  reg [511:0] chn_relu_in_rsci_d_bfwt;
// Interconnect Declarations for Component Instantiations
  assign chn_relu_in_rsci_bawt = chn_relu_in_rsci_biwt | chn_relu_in_rsci_bcwt;
  assign chn_relu_in_rsci_wen_comp = (~ chn_relu_in_rsci_oswt) | chn_relu_in_rsci_bawt;
  assign chn_relu_in_rsci_d_mxwt = MUX_v_512_2_2(chn_relu_in_rsci_d, chn_relu_in_rsci_d_bfwt,
      chn_relu_in_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_relu_in_rsci_bcwt <= 1'b0;
      chn_relu_in_rsci_d_bfwt <= 512'b0;
    end
    else begin
      chn_relu_in_rsci_bcwt <= ~((~(chn_relu_in_rsci_bcwt | chn_relu_in_rsci_biwt))
          | chn_relu_in_rsci_bdwt);
      chn_relu_in_rsci_d_bfwt <= chn_relu_in_rsci_d_mxwt;
    end
  end
  function [511:0] MUX_v_512_2_2;
    input [511:0] input_0;
    input [511:0] input_1;
    input [0:0] sel;
    reg [511:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_512_2_2 = result;
  end
  endfunction
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_relu_core_chn_relu_in_rsci_chn_relu_in_wait_ctrl
// ------------------------------------------------------------------
module SDP_X_X_relu_core_chn_relu_in_rsci_chn_relu_in_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_relu_in_rsci_oswt, core_wen, chn_relu_in_rsci_iswt0,
      chn_relu_in_rsci_ld_core_psct, core_wten, chn_relu_in_rsci_biwt, chn_relu_in_rsci_bdwt,
      chn_relu_in_rsci_ld_core_sct, chn_relu_in_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_relu_in_rsci_oswt;
  input core_wen;
  input chn_relu_in_rsci_iswt0;
  input chn_relu_in_rsci_ld_core_psct;
  input core_wten;
  output chn_relu_in_rsci_biwt;
  output chn_relu_in_rsci_bdwt;
  output chn_relu_in_rsci_ld_core_sct;
  input chn_relu_in_rsci_vd;
// Interconnect Declarations
  wire chn_relu_in_rsci_ogwt;
  wire chn_relu_in_rsci_pdswt0;
  reg chn_relu_in_rsci_icwt;
// Interconnect Declarations for Component Instantiations
  assign chn_relu_in_rsci_pdswt0 = (~ core_wten) & chn_relu_in_rsci_iswt0;
  assign chn_relu_in_rsci_biwt = chn_relu_in_rsci_ogwt & chn_relu_in_rsci_vd;
  assign chn_relu_in_rsci_ogwt = chn_relu_in_rsci_pdswt0 | chn_relu_in_rsci_icwt;
  assign chn_relu_in_rsci_bdwt = chn_relu_in_rsci_oswt & core_wen;
  assign chn_relu_in_rsci_ld_core_sct = chn_relu_in_rsci_ld_core_psct & chn_relu_in_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_relu_in_rsci_icwt <= 1'b0;
    end
    else begin
      chn_relu_in_rsci_icwt <= ~((~(chn_relu_in_rsci_icwt | chn_relu_in_rsci_pdswt0))
          | chn_relu_in_rsci_biwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_cfg_alu_shift_value_rsc_triosy_obj
// ------------------------------------------------------------------
module SDP_X_X_alu_core_cfg_alu_shift_value_rsc_triosy_obj (
  nvdla_core_clk, nvdla_core_rstn, cfg_alu_shift_value_rsc_triosy_lz, cfg_alu_shift_value_rsc_triosy_obj_oswt,
      core_wen, core_wten, cfg_alu_shift_value_rsc_triosy_obj_iswt0, cfg_alu_shift_value_rsc_triosy_obj_bawt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_alu_shift_value_rsc_triosy_lz;
  input cfg_alu_shift_value_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_alu_shift_value_rsc_triosy_obj_iswt0;
  output cfg_alu_shift_value_rsc_triosy_obj_bawt;
// Interconnect Declarations
  wire cfg_alu_shift_value_rsc_triosy_obj_biwt;
  wire cfg_alu_shift_value_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_io_sync_v1 #(.valid(32'sd0)) cfg_alu_shift_value_rsc_triosy_obj (
      .ld(cfg_alu_shift_value_rsc_triosy_obj_biwt),
      .lz(cfg_alu_shift_value_rsc_triosy_lz)
    );
  SDP_X_X_alu_core_cfg_alu_shift_value_rsc_triosy_obj_cfg_alu_shift_value_rsc_triosy_wait_ctrl
      X_alu_core_cfg_alu_shift_value_rsc_triosy_obj_cfg_alu_shift_value_rsc_triosy_wait_ctrl_inst
      (
      .cfg_alu_shift_value_rsc_triosy_obj_oswt(cfg_alu_shift_value_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_alu_shift_value_rsc_triosy_obj_iswt0(cfg_alu_shift_value_rsc_triosy_obj_iswt0),
      .cfg_alu_shift_value_rsc_triosy_obj_biwt(cfg_alu_shift_value_rsc_triosy_obj_biwt),
      .cfg_alu_shift_value_rsc_triosy_obj_bdwt(cfg_alu_shift_value_rsc_triosy_obj_bdwt)
    );
  SDP_X_X_alu_core_cfg_alu_shift_value_rsc_triosy_obj_cfg_alu_shift_value_rsc_triosy_wait_dp
      X_alu_core_cfg_alu_shift_value_rsc_triosy_obj_cfg_alu_shift_value_rsc_triosy_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_alu_shift_value_rsc_triosy_obj_bawt(cfg_alu_shift_value_rsc_triosy_obj_bawt),
      .cfg_alu_shift_value_rsc_triosy_obj_biwt(cfg_alu_shift_value_rsc_triosy_obj_biwt),
      .cfg_alu_shift_value_rsc_triosy_obj_bdwt(cfg_alu_shift_value_rsc_triosy_obj_bdwt)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_cfg_alu_src_rsc_triosy_obj
// ------------------------------------------------------------------
module SDP_X_X_alu_core_cfg_alu_src_rsc_triosy_obj (
  nvdla_core_clk, nvdla_core_rstn, cfg_alu_src_rsc_triosy_lz, cfg_alu_src_rsc_triosy_obj_oswt,
      core_wen, core_wten, cfg_alu_src_rsc_triosy_obj_iswt0, cfg_alu_src_rsc_triosy_obj_bawt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_alu_src_rsc_triosy_lz;
  input cfg_alu_src_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_alu_src_rsc_triosy_obj_iswt0;
  output cfg_alu_src_rsc_triosy_obj_bawt;
// Interconnect Declarations
  wire cfg_alu_src_rsc_triosy_obj_biwt;
  wire cfg_alu_src_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_io_sync_v1 #(.valid(32'sd0)) cfg_alu_src_rsc_triosy_obj (
      .ld(cfg_alu_src_rsc_triosy_obj_biwt),
      .lz(cfg_alu_src_rsc_triosy_lz)
    );
  SDP_X_X_alu_core_cfg_alu_src_rsc_triosy_obj_cfg_alu_src_rsc_triosy_wait_ctrl X_alu_core_cfg_alu_src_rsc_triosy_obj_cfg_alu_src_rsc_triosy_wait_ctrl_inst
      (
      .cfg_alu_src_rsc_triosy_obj_oswt(cfg_alu_src_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_alu_src_rsc_triosy_obj_iswt0(cfg_alu_src_rsc_triosy_obj_iswt0),
      .cfg_alu_src_rsc_triosy_obj_biwt(cfg_alu_src_rsc_triosy_obj_biwt),
      .cfg_alu_src_rsc_triosy_obj_bdwt(cfg_alu_src_rsc_triosy_obj_bdwt)
    );
  SDP_X_X_alu_core_cfg_alu_src_rsc_triosy_obj_cfg_alu_src_rsc_triosy_wait_dp X_alu_core_cfg_alu_src_rsc_triosy_obj_cfg_alu_src_rsc_triosy_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_alu_src_rsc_triosy_obj_bawt(cfg_alu_src_rsc_triosy_obj_bawt),
      .cfg_alu_src_rsc_triosy_obj_biwt(cfg_alu_src_rsc_triosy_obj_biwt),
      .cfg_alu_src_rsc_triosy_obj_bdwt(cfg_alu_src_rsc_triosy_obj_bdwt)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_cfg_alu_algo_rsc_triosy_obj
// ------------------------------------------------------------------
module SDP_X_X_alu_core_cfg_alu_algo_rsc_triosy_obj (
  nvdla_core_clk, nvdla_core_rstn, cfg_alu_algo_rsc_triosy_lz, cfg_alu_algo_rsc_triosy_obj_oswt,
      core_wen, core_wten, cfg_alu_algo_rsc_triosy_obj_iswt0, cfg_alu_algo_rsc_triosy_obj_bawt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_alu_algo_rsc_triosy_lz;
  input cfg_alu_algo_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_alu_algo_rsc_triosy_obj_iswt0;
  output cfg_alu_algo_rsc_triosy_obj_bawt;
// Interconnect Declarations
  wire cfg_alu_algo_rsc_triosy_obj_biwt;
  wire cfg_alu_algo_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_io_sync_v1 #(.valid(32'sd0)) cfg_alu_algo_rsc_triosy_obj (
      .ld(cfg_alu_algo_rsc_triosy_obj_biwt),
      .lz(cfg_alu_algo_rsc_triosy_lz)
    );
  SDP_X_X_alu_core_cfg_alu_algo_rsc_triosy_obj_cfg_alu_algo_rsc_triosy_wait_ctrl X_alu_core_cfg_alu_algo_rsc_triosy_obj_cfg_alu_algo_rsc_triosy_wait_ctrl_inst
      (
      .cfg_alu_algo_rsc_triosy_obj_oswt(cfg_alu_algo_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_alu_algo_rsc_triosy_obj_iswt0(cfg_alu_algo_rsc_triosy_obj_iswt0),
      .cfg_alu_algo_rsc_triosy_obj_biwt(cfg_alu_algo_rsc_triosy_obj_biwt),
      .cfg_alu_algo_rsc_triosy_obj_bdwt(cfg_alu_algo_rsc_triosy_obj_bdwt)
    );
  SDP_X_X_alu_core_cfg_alu_algo_rsc_triosy_obj_cfg_alu_algo_rsc_triosy_wait_dp X_alu_core_cfg_alu_algo_rsc_triosy_obj_cfg_alu_algo_rsc_triosy_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_alu_algo_rsc_triosy_obj_bawt(cfg_alu_algo_rsc_triosy_obj_bawt),
      .cfg_alu_algo_rsc_triosy_obj_biwt(cfg_alu_algo_rsc_triosy_obj_biwt),
      .cfg_alu_algo_rsc_triosy_obj_bdwt(cfg_alu_algo_rsc_triosy_obj_bdwt)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_cfg_alu_bypass_rsc_triosy_obj
// ------------------------------------------------------------------
module SDP_X_X_alu_core_cfg_alu_bypass_rsc_triosy_obj (
  nvdla_core_clk, nvdla_core_rstn, cfg_alu_bypass_rsc_triosy_lz, cfg_alu_bypass_rsc_triosy_obj_oswt,
      core_wen, core_wten, cfg_alu_bypass_rsc_triosy_obj_iswt0, cfg_alu_bypass_rsc_triosy_obj_bawt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_alu_bypass_rsc_triosy_lz;
  input cfg_alu_bypass_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_alu_bypass_rsc_triosy_obj_iswt0;
  output cfg_alu_bypass_rsc_triosy_obj_bawt;
// Interconnect Declarations
  wire cfg_alu_bypass_rsc_triosy_obj_biwt;
  wire cfg_alu_bypass_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_io_sync_v1 #(.valid(32'sd0)) cfg_alu_bypass_rsc_triosy_obj (
      .ld(cfg_alu_bypass_rsc_triosy_obj_biwt),
      .lz(cfg_alu_bypass_rsc_triosy_lz)
    );
  SDP_X_X_alu_core_cfg_alu_bypass_rsc_triosy_obj_cfg_alu_bypass_rsc_triosy_wait_ctrl X_alu_core_cfg_alu_bypass_rsc_triosy_obj_cfg_alu_bypass_rsc_triosy_wait_ctrl_inst
      (
      .cfg_alu_bypass_rsc_triosy_obj_oswt(cfg_alu_bypass_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_alu_bypass_rsc_triosy_obj_iswt0(cfg_alu_bypass_rsc_triosy_obj_iswt0),
      .cfg_alu_bypass_rsc_triosy_obj_biwt(cfg_alu_bypass_rsc_triosy_obj_biwt),
      .cfg_alu_bypass_rsc_triosy_obj_bdwt(cfg_alu_bypass_rsc_triosy_obj_bdwt)
    );
  SDP_X_X_alu_core_cfg_alu_bypass_rsc_triosy_obj_cfg_alu_bypass_rsc_triosy_wait_dp X_alu_core_cfg_alu_bypass_rsc_triosy_obj_cfg_alu_bypass_rsc_triosy_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_alu_bypass_rsc_triosy_obj_bawt(cfg_alu_bypass_rsc_triosy_obj_bawt),
      .cfg_alu_bypass_rsc_triosy_obj_biwt(cfg_alu_bypass_rsc_triosy_obj_biwt),
      .cfg_alu_bypass_rsc_triosy_obj_bdwt(cfg_alu_bypass_rsc_triosy_obj_bdwt)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_cfg_alu_op_rsc_triosy_obj
// ------------------------------------------------------------------
module SDP_X_X_alu_core_cfg_alu_op_rsc_triosy_obj (
  nvdla_core_clk, nvdla_core_rstn, cfg_alu_op_rsc_triosy_lz, cfg_alu_op_rsc_triosy_obj_oswt,
      core_wen, core_wten, cfg_alu_op_rsc_triosy_obj_iswt0, cfg_alu_op_rsc_triosy_obj_bawt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_alu_op_rsc_triosy_lz;
  input cfg_alu_op_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_alu_op_rsc_triosy_obj_iswt0;
  output cfg_alu_op_rsc_triosy_obj_bawt;
// Interconnect Declarations
  wire cfg_alu_op_rsc_triosy_obj_biwt;
  wire cfg_alu_op_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_io_sync_v1 #(.valid(32'sd0)) cfg_alu_op_rsc_triosy_obj (
      .ld(cfg_alu_op_rsc_triosy_obj_biwt),
      .lz(cfg_alu_op_rsc_triosy_lz)
    );
  SDP_X_X_alu_core_cfg_alu_op_rsc_triosy_obj_cfg_alu_op_rsc_triosy_wait_ctrl X_alu_core_cfg_alu_op_rsc_triosy_obj_cfg_alu_op_rsc_triosy_wait_ctrl_inst
      (
      .cfg_alu_op_rsc_triosy_obj_oswt(cfg_alu_op_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_alu_op_rsc_triosy_obj_iswt0(cfg_alu_op_rsc_triosy_obj_iswt0),
      .cfg_alu_op_rsc_triosy_obj_biwt(cfg_alu_op_rsc_triosy_obj_biwt),
      .cfg_alu_op_rsc_triosy_obj_bdwt(cfg_alu_op_rsc_triosy_obj_bdwt)
    );
  SDP_X_X_alu_core_cfg_alu_op_rsc_triosy_obj_cfg_alu_op_rsc_triosy_wait_dp X_alu_core_cfg_alu_op_rsc_triosy_obj_cfg_alu_op_rsc_triosy_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_alu_op_rsc_triosy_obj_bawt(cfg_alu_op_rsc_triosy_obj_bawt),
      .cfg_alu_op_rsc_triosy_obj_biwt(cfg_alu_op_rsc_triosy_obj_biwt),
      .cfg_alu_op_rsc_triosy_obj_bdwt(cfg_alu_op_rsc_triosy_obj_bdwt)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_chn_alu_out_rsci
// ------------------------------------------------------------------
module SDP_X_X_alu_core_chn_alu_out_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_out_rsc_z, chn_alu_out_rsc_vz, chn_alu_out_rsc_lz,
      chn_alu_out_rsci_oswt, core_wen, core_wten, chn_alu_out_rsci_iswt0, chn_alu_out_rsci_bawt,
      chn_alu_out_rsci_wen_comp, chn_alu_out_rsci_ld_core_psct, chn_alu_out_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output [527:0] chn_alu_out_rsc_z;
  input chn_alu_out_rsc_vz;
  output chn_alu_out_rsc_lz;
  input chn_alu_out_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_alu_out_rsci_iswt0;
  output chn_alu_out_rsci_bawt;
  output chn_alu_out_rsci_wen_comp;
  input chn_alu_out_rsci_ld_core_psct;
  input [527:0] chn_alu_out_rsci_d;
// Interconnect Declarations
  wire chn_alu_out_rsci_biwt;
  wire chn_alu_out_rsci_bdwt;
  wire chn_alu_out_rsci_ld_core_sct;
  wire chn_alu_out_rsci_vd;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_out_stdreg_wait_v1 #(.rscid(32'sd10),
  .width(32'sd528)) chn_alu_out_rsci (
      .ld(chn_alu_out_rsci_ld_core_sct),
      .vd(chn_alu_out_rsci_vd),
      .d(chn_alu_out_rsci_d),
      .lz(chn_alu_out_rsc_lz),
      .vz(chn_alu_out_rsc_vz),
      .z(chn_alu_out_rsc_z)
    );
  SDP_X_X_alu_core_chn_alu_out_rsci_chn_alu_out_wait_ctrl X_alu_core_chn_alu_out_rsci_chn_alu_out_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_out_rsci_oswt(chn_alu_out_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_alu_out_rsci_iswt0(chn_alu_out_rsci_iswt0),
      .chn_alu_out_rsci_ld_core_psct(chn_alu_out_rsci_ld_core_psct),
      .chn_alu_out_rsci_biwt(chn_alu_out_rsci_biwt),
      .chn_alu_out_rsci_bdwt(chn_alu_out_rsci_bdwt),
      .chn_alu_out_rsci_ld_core_sct(chn_alu_out_rsci_ld_core_sct),
      .chn_alu_out_rsci_vd(chn_alu_out_rsci_vd)
    );
  SDP_X_X_alu_core_chn_alu_out_rsci_chn_alu_out_wait_dp X_alu_core_chn_alu_out_rsci_chn_alu_out_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_out_rsci_oswt(chn_alu_out_rsci_oswt),
      .chn_alu_out_rsci_bawt(chn_alu_out_rsci_bawt),
      .chn_alu_out_rsci_wen_comp(chn_alu_out_rsci_wen_comp),
      .chn_alu_out_rsci_biwt(chn_alu_out_rsci_biwt),
      .chn_alu_out_rsci_bdwt(chn_alu_out_rsci_bdwt)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_chn_alu_op_rsci
// ------------------------------------------------------------------
module SDP_X_X_alu_core_chn_alu_op_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_op_rsc_z, chn_alu_op_rsc_vz, chn_alu_op_rsc_lz,
      chn_alu_op_rsci_oswt, core_wen, core_wten, chn_alu_op_rsci_iswt0, chn_alu_op_rsci_bawt,
      chn_alu_op_rsci_wen_comp, chn_alu_op_rsci_ld_core_psct, chn_alu_op_rsci_d_mxwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [255:0] chn_alu_op_rsc_z;
  input chn_alu_op_rsc_vz;
  output chn_alu_op_rsc_lz;
  input chn_alu_op_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_alu_op_rsci_iswt0;
  output chn_alu_op_rsci_bawt;
  output chn_alu_op_rsci_wen_comp;
  input chn_alu_op_rsci_ld_core_psct;
  output [255:0] chn_alu_op_rsci_d_mxwt;
// Interconnect Declarations
  wire chn_alu_op_rsci_biwt;
  wire chn_alu_op_rsci_bdwt;
  wire chn_alu_op_rsci_ld_core_sct;
  wire chn_alu_op_rsci_vd;
  wire [255:0] chn_alu_op_rsci_d;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_in_wire_wait_v1 #(.rscid(32'sd2),
  .width(32'sd256)) chn_alu_op_rsci (
      .ld(chn_alu_op_rsci_ld_core_sct),
      .vd(chn_alu_op_rsci_vd),
      .d(chn_alu_op_rsci_d),
      .lz(chn_alu_op_rsc_lz),
      .vz(chn_alu_op_rsc_vz),
      .z(chn_alu_op_rsc_z)
    );
  SDP_X_X_alu_core_chn_alu_op_rsci_chn_alu_op_wait_ctrl X_alu_core_chn_alu_op_rsci_chn_alu_op_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_op_rsci_oswt(chn_alu_op_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_alu_op_rsci_iswt0(chn_alu_op_rsci_iswt0),
      .chn_alu_op_rsci_ld_core_psct(chn_alu_op_rsci_ld_core_psct),
      .chn_alu_op_rsci_biwt(chn_alu_op_rsci_biwt),
      .chn_alu_op_rsci_bdwt(chn_alu_op_rsci_bdwt),
      .chn_alu_op_rsci_ld_core_sct(chn_alu_op_rsci_ld_core_sct),
      .chn_alu_op_rsci_vd(chn_alu_op_rsci_vd)
    );
  SDP_X_X_alu_core_chn_alu_op_rsci_chn_alu_op_wait_dp X_alu_core_chn_alu_op_rsci_chn_alu_op_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_op_rsci_oswt(chn_alu_op_rsci_oswt),
      .chn_alu_op_rsci_bawt(chn_alu_op_rsci_bawt),
      .chn_alu_op_rsci_wen_comp(chn_alu_op_rsci_wen_comp),
      .chn_alu_op_rsci_d_mxwt(chn_alu_op_rsci_d_mxwt),
      .chn_alu_op_rsci_biwt(chn_alu_op_rsci_biwt),
      .chn_alu_op_rsci_bdwt(chn_alu_op_rsci_bdwt),
      .chn_alu_op_rsci_d(chn_alu_op_rsci_d)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core_chn_alu_in_rsci
// ------------------------------------------------------------------
module SDP_X_X_alu_core_chn_alu_in_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_in_rsc_z, chn_alu_in_rsc_vz, chn_alu_in_rsc_lz,
      chn_alu_in_rsci_oswt, core_wen, chn_alu_in_rsci_iswt0, chn_alu_in_rsci_bawt,
      chn_alu_in_rsci_wen_comp, chn_alu_in_rsci_ld_core_psct, chn_alu_in_rsci_d_mxwt,
      core_wten
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [511:0] chn_alu_in_rsc_z;
  input chn_alu_in_rsc_vz;
  output chn_alu_in_rsc_lz;
  input chn_alu_in_rsci_oswt;
  input core_wen;
  input chn_alu_in_rsci_iswt0;
  output chn_alu_in_rsci_bawt;
  output chn_alu_in_rsci_wen_comp;
  input chn_alu_in_rsci_ld_core_psct;
  output [511:0] chn_alu_in_rsci_d_mxwt;
  input core_wten;
// Interconnect Declarations
  wire chn_alu_in_rsci_biwt;
  wire chn_alu_in_rsci_bdwt;
  wire chn_alu_in_rsci_ld_core_sct;
  wire chn_alu_in_rsci_vd;
  wire [511:0] chn_alu_in_rsci_d;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_in_wire_wait_v1 #(.rscid(32'sd1),
  .width(32'sd512)) chn_alu_in_rsci (
      .ld(chn_alu_in_rsci_ld_core_sct),
      .vd(chn_alu_in_rsci_vd),
      .d(chn_alu_in_rsci_d),
      .lz(chn_alu_in_rsc_lz),
      .vz(chn_alu_in_rsc_vz),
      .z(chn_alu_in_rsc_z)
    );
  SDP_X_X_alu_core_chn_alu_in_rsci_chn_alu_in_wait_ctrl X_alu_core_chn_alu_in_rsci_chn_alu_in_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_in_rsci_oswt(chn_alu_in_rsci_oswt),
      .core_wen(core_wen),
      .chn_alu_in_rsci_iswt0(chn_alu_in_rsci_iswt0),
      .chn_alu_in_rsci_ld_core_psct(chn_alu_in_rsci_ld_core_psct),
      .core_wten(core_wten),
      .chn_alu_in_rsci_biwt(chn_alu_in_rsci_biwt),
      .chn_alu_in_rsci_bdwt(chn_alu_in_rsci_bdwt),
      .chn_alu_in_rsci_ld_core_sct(chn_alu_in_rsci_ld_core_sct),
      .chn_alu_in_rsci_vd(chn_alu_in_rsci_vd)
    );
  SDP_X_X_alu_core_chn_alu_in_rsci_chn_alu_in_wait_dp X_alu_core_chn_alu_in_rsci_chn_alu_in_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_in_rsci_oswt(chn_alu_in_rsci_oswt),
      .chn_alu_in_rsci_bawt(chn_alu_in_rsci_bawt),
      .chn_alu_in_rsci_wen_comp(chn_alu_in_rsci_wen_comp),
      .chn_alu_in_rsci_d_mxwt(chn_alu_in_rsci_d_mxwt),
      .chn_alu_in_rsci_biwt(chn_alu_in_rsci_biwt),
      .chn_alu_in_rsci_bdwt(chn_alu_in_rsci_bdwt),
      .chn_alu_in_rsci_d(chn_alu_in_rsci_d)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_cfg_mul_src_rsc_triosy_obj
// ------------------------------------------------------------------
module SDP_X_X_mul_core_cfg_mul_src_rsc_triosy_obj (
  nvdla_core_clk, nvdla_core_rstn, cfg_mul_src_rsc_triosy_lz, cfg_mul_src_rsc_triosy_obj_oswt,
      core_wen, core_wten, cfg_mul_src_rsc_triosy_obj_iswt0, cfg_mul_src_rsc_triosy_obj_bawt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_mul_src_rsc_triosy_lz;
  input cfg_mul_src_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_mul_src_rsc_triosy_obj_iswt0;
  output cfg_mul_src_rsc_triosy_obj_bawt;
// Interconnect Declarations
  wire cfg_mul_src_rsc_triosy_obj_biwt;
  wire cfg_mul_src_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_io_sync_v1 #(.valid(32'sd0)) cfg_mul_src_rsc_triosy_obj (
      .ld(cfg_mul_src_rsc_triosy_obj_biwt),
      .lz(cfg_mul_src_rsc_triosy_lz)
    );
  SDP_X_X_mul_core_cfg_mul_src_rsc_triosy_obj_cfg_mul_src_rsc_triosy_wait_ctrl X_mul_core_cfg_mul_src_rsc_triosy_obj_cfg_mul_src_rsc_triosy_wait_ctrl_inst
      (
      .cfg_mul_src_rsc_triosy_obj_oswt(cfg_mul_src_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_mul_src_rsc_triosy_obj_iswt0(cfg_mul_src_rsc_triosy_obj_iswt0),
      .cfg_mul_src_rsc_triosy_obj_biwt(cfg_mul_src_rsc_triosy_obj_biwt),
      .cfg_mul_src_rsc_triosy_obj_bdwt(cfg_mul_src_rsc_triosy_obj_bdwt)
    );
  SDP_X_X_mul_core_cfg_mul_src_rsc_triosy_obj_cfg_mul_src_rsc_triosy_wait_dp X_mul_core_cfg_mul_src_rsc_triosy_obj_cfg_mul_src_rsc_triosy_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_mul_src_rsc_triosy_obj_bawt(cfg_mul_src_rsc_triosy_obj_bawt),
      .cfg_mul_src_rsc_triosy_obj_biwt(cfg_mul_src_rsc_triosy_obj_biwt),
      .cfg_mul_src_rsc_triosy_obj_bdwt(cfg_mul_src_rsc_triosy_obj_bdwt)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_cfg_mul_prelu_rsc_triosy_obj
// ------------------------------------------------------------------
module SDP_X_X_mul_core_cfg_mul_prelu_rsc_triosy_obj (
  nvdla_core_clk, nvdla_core_rstn, cfg_mul_prelu_rsc_triosy_lz, cfg_mul_prelu_rsc_triosy_obj_oswt,
      core_wen, core_wten, cfg_mul_prelu_rsc_triosy_obj_iswt0, cfg_mul_prelu_rsc_triosy_obj_bawt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_mul_prelu_rsc_triosy_lz;
  input cfg_mul_prelu_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_mul_prelu_rsc_triosy_obj_iswt0;
  output cfg_mul_prelu_rsc_triosy_obj_bawt;
// Interconnect Declarations
  wire cfg_mul_prelu_rsc_triosy_obj_biwt;
  wire cfg_mul_prelu_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_io_sync_v1 #(.valid(32'sd0)) cfg_mul_prelu_rsc_triosy_obj (
      .ld(cfg_mul_prelu_rsc_triosy_obj_biwt),
      .lz(cfg_mul_prelu_rsc_triosy_lz)
    );
  SDP_X_X_mul_core_cfg_mul_prelu_rsc_triosy_obj_cfg_mul_prelu_rsc_triosy_wait_ctrl X_mul_core_cfg_mul_prelu_rsc_triosy_obj_cfg_mul_prelu_rsc_triosy_wait_ctrl_inst
      (
      .cfg_mul_prelu_rsc_triosy_obj_oswt(cfg_mul_prelu_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_mul_prelu_rsc_triosy_obj_iswt0(cfg_mul_prelu_rsc_triosy_obj_iswt0),
      .cfg_mul_prelu_rsc_triosy_obj_biwt(cfg_mul_prelu_rsc_triosy_obj_biwt),
      .cfg_mul_prelu_rsc_triosy_obj_bdwt(cfg_mul_prelu_rsc_triosy_obj_bdwt)
    );
  SDP_X_X_mul_core_cfg_mul_prelu_rsc_triosy_obj_cfg_mul_prelu_rsc_triosy_wait_dp X_mul_core_cfg_mul_prelu_rsc_triosy_obj_cfg_mul_prelu_rsc_triosy_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_mul_prelu_rsc_triosy_obj_bawt(cfg_mul_prelu_rsc_triosy_obj_bawt),
      .cfg_mul_prelu_rsc_triosy_obj_biwt(cfg_mul_prelu_rsc_triosy_obj_biwt),
      .cfg_mul_prelu_rsc_triosy_obj_bdwt(cfg_mul_prelu_rsc_triosy_obj_bdwt)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_cfg_mul_bypass_rsc_triosy_obj
// ------------------------------------------------------------------
module SDP_X_X_mul_core_cfg_mul_bypass_rsc_triosy_obj (
  nvdla_core_clk, nvdla_core_rstn, cfg_mul_bypass_rsc_triosy_lz, cfg_mul_bypass_rsc_triosy_obj_oswt,
      core_wen, core_wten, cfg_mul_bypass_rsc_triosy_obj_iswt0, cfg_mul_bypass_rsc_triosy_obj_bawt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_mul_bypass_rsc_triosy_lz;
  input cfg_mul_bypass_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_mul_bypass_rsc_triosy_obj_iswt0;
  output cfg_mul_bypass_rsc_triosy_obj_bawt;
// Interconnect Declarations
  wire cfg_mul_bypass_rsc_triosy_obj_biwt;
  wire cfg_mul_bypass_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_io_sync_v1 #(.valid(32'sd0)) cfg_mul_bypass_rsc_triosy_obj (
      .ld(cfg_mul_bypass_rsc_triosy_obj_biwt),
      .lz(cfg_mul_bypass_rsc_triosy_lz)
    );
  SDP_X_X_mul_core_cfg_mul_bypass_rsc_triosy_obj_cfg_mul_bypass_rsc_triosy_wait_ctrl X_mul_core_cfg_mul_bypass_rsc_triosy_obj_cfg_mul_bypass_rsc_triosy_wait_ctrl_inst
      (
      .cfg_mul_bypass_rsc_triosy_obj_oswt(cfg_mul_bypass_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_mul_bypass_rsc_triosy_obj_iswt0(cfg_mul_bypass_rsc_triosy_obj_iswt0),
      .cfg_mul_bypass_rsc_triosy_obj_biwt(cfg_mul_bypass_rsc_triosy_obj_biwt),
      .cfg_mul_bypass_rsc_triosy_obj_bdwt(cfg_mul_bypass_rsc_triosy_obj_bdwt)
    );
  SDP_X_X_mul_core_cfg_mul_bypass_rsc_triosy_obj_cfg_mul_bypass_rsc_triosy_wait_dp X_mul_core_cfg_mul_bypass_rsc_triosy_obj_cfg_mul_bypass_rsc_triosy_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_mul_bypass_rsc_triosy_obj_bawt(cfg_mul_bypass_rsc_triosy_obj_bawt),
      .cfg_mul_bypass_rsc_triosy_obj_biwt(cfg_mul_bypass_rsc_triosy_obj_biwt),
      .cfg_mul_bypass_rsc_triosy_obj_bdwt(cfg_mul_bypass_rsc_triosy_obj_bdwt)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_cfg_mul_op_rsc_triosy_obj
// ------------------------------------------------------------------
module SDP_X_X_mul_core_cfg_mul_op_rsc_triosy_obj (
  nvdla_core_clk, nvdla_core_rstn, cfg_mul_op_rsc_triosy_lz, cfg_mul_op_rsc_triosy_obj_oswt,
      core_wen, core_wten, cfg_mul_op_rsc_triosy_obj_iswt0, cfg_mul_op_rsc_triosy_obj_bawt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_mul_op_rsc_triosy_lz;
  input cfg_mul_op_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_mul_op_rsc_triosy_obj_iswt0;
  output cfg_mul_op_rsc_triosy_obj_bawt;
// Interconnect Declarations
  wire cfg_mul_op_rsc_triosy_obj_biwt;
  wire cfg_mul_op_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_io_sync_v1 #(.valid(32'sd0)) cfg_mul_op_rsc_triosy_obj (
      .ld(cfg_mul_op_rsc_triosy_obj_biwt),
      .lz(cfg_mul_op_rsc_triosy_lz)
    );
  SDP_X_X_mul_core_cfg_mul_op_rsc_triosy_obj_cfg_mul_op_rsc_triosy_wait_ctrl X_mul_core_cfg_mul_op_rsc_triosy_obj_cfg_mul_op_rsc_triosy_wait_ctrl_inst
      (
      .cfg_mul_op_rsc_triosy_obj_oswt(cfg_mul_op_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_mul_op_rsc_triosy_obj_iswt0(cfg_mul_op_rsc_triosy_obj_iswt0),
      .cfg_mul_op_rsc_triosy_obj_biwt(cfg_mul_op_rsc_triosy_obj_biwt),
      .cfg_mul_op_rsc_triosy_obj_bdwt(cfg_mul_op_rsc_triosy_obj_bdwt)
    );
  SDP_X_X_mul_core_cfg_mul_op_rsc_triosy_obj_cfg_mul_op_rsc_triosy_wait_dp X_mul_core_cfg_mul_op_rsc_triosy_obj_cfg_mul_op_rsc_triosy_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_mul_op_rsc_triosy_obj_bawt(cfg_mul_op_rsc_triosy_obj_bawt),
      .cfg_mul_op_rsc_triosy_obj_biwt(cfg_mul_op_rsc_triosy_obj_biwt),
      .cfg_mul_op_rsc_triosy_obj_bdwt(cfg_mul_op_rsc_triosy_obj_bdwt)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_chn_mul_out_rsci
// ------------------------------------------------------------------
module SDP_X_X_mul_core_chn_mul_out_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_out_rsc_z, chn_mul_out_rsc_vz, chn_mul_out_rsc_lz,
      chn_mul_out_rsci_oswt, core_wen, core_wten, chn_mul_out_rsci_iswt0, chn_mul_out_rsci_bawt,
      chn_mul_out_rsci_wen_comp, chn_mul_out_rsci_ld_core_psct, chn_mul_out_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output [799:0] chn_mul_out_rsc_z;
  input chn_mul_out_rsc_vz;
  output chn_mul_out_rsc_lz;
  input chn_mul_out_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_mul_out_rsci_iswt0;
  output chn_mul_out_rsci_bawt;
  output chn_mul_out_rsci_wen_comp;
  input chn_mul_out_rsci_ld_core_psct;
  input [799:0] chn_mul_out_rsci_d;
// Interconnect Declarations
  wire chn_mul_out_rsci_biwt;
  wire chn_mul_out_rsci_bdwt;
  wire chn_mul_out_rsci_ld_core_sct;
  wire chn_mul_out_rsci_vd;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_out_stdreg_wait_v1 #(.rscid(32'sd22),
  .width(32'sd800)) chn_mul_out_rsci (
      .ld(chn_mul_out_rsci_ld_core_sct),
      .vd(chn_mul_out_rsci_vd),
      .d(chn_mul_out_rsci_d),
      .lz(chn_mul_out_rsc_lz),
      .vz(chn_mul_out_rsc_vz),
      .z(chn_mul_out_rsc_z)
    );
  SDP_X_X_mul_core_chn_mul_out_rsci_chn_mul_out_wait_ctrl X_mul_core_chn_mul_out_rsci_chn_mul_out_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_out_rsci_oswt(chn_mul_out_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_mul_out_rsci_iswt0(chn_mul_out_rsci_iswt0),
      .chn_mul_out_rsci_ld_core_psct(chn_mul_out_rsci_ld_core_psct),
      .chn_mul_out_rsci_biwt(chn_mul_out_rsci_biwt),
      .chn_mul_out_rsci_bdwt(chn_mul_out_rsci_bdwt),
      .chn_mul_out_rsci_ld_core_sct(chn_mul_out_rsci_ld_core_sct),
      .chn_mul_out_rsci_vd(chn_mul_out_rsci_vd)
    );
  SDP_X_X_mul_core_chn_mul_out_rsci_chn_mul_out_wait_dp X_mul_core_chn_mul_out_rsci_chn_mul_out_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_out_rsci_oswt(chn_mul_out_rsci_oswt),
      .chn_mul_out_rsci_bawt(chn_mul_out_rsci_bawt),
      .chn_mul_out_rsci_wen_comp(chn_mul_out_rsci_wen_comp),
      .chn_mul_out_rsci_biwt(chn_mul_out_rsci_biwt),
      .chn_mul_out_rsci_bdwt(chn_mul_out_rsci_bdwt)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_chn_mul_op_rsci
// ------------------------------------------------------------------
module SDP_X_X_mul_core_chn_mul_op_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_op_rsc_z, chn_mul_op_rsc_vz, chn_mul_op_rsc_lz,
      chn_mul_op_rsci_oswt, core_wen, core_wten, chn_mul_op_rsci_iswt0, chn_mul_op_rsci_bawt,
      chn_mul_op_rsci_wen_comp, chn_mul_op_rsci_ld_core_psct, chn_mul_op_rsci_d_mxwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [255:0] chn_mul_op_rsc_z;
  input chn_mul_op_rsc_vz;
  output chn_mul_op_rsc_lz;
  input chn_mul_op_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_mul_op_rsci_iswt0;
  output chn_mul_op_rsci_bawt;
  output chn_mul_op_rsci_wen_comp;
  input chn_mul_op_rsci_ld_core_psct;
  output [255:0] chn_mul_op_rsci_d_mxwt;
// Interconnect Declarations
  wire chn_mul_op_rsci_biwt;
  wire chn_mul_op_rsci_bdwt;
  wire chn_mul_op_rsci_ld_core_sct;
  wire chn_mul_op_rsci_vd;
  wire [255:0] chn_mul_op_rsci_d;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_in_wire_wait_v1 #(.rscid(32'sd15),
  .width(32'sd256)) chn_mul_op_rsci (
      .ld(chn_mul_op_rsci_ld_core_sct),
      .vd(chn_mul_op_rsci_vd),
      .d(chn_mul_op_rsci_d),
      .lz(chn_mul_op_rsc_lz),
      .vz(chn_mul_op_rsc_vz),
      .z(chn_mul_op_rsc_z)
    );
  SDP_X_X_mul_core_chn_mul_op_rsci_chn_mul_op_wait_ctrl X_mul_core_chn_mul_op_rsci_chn_mul_op_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_op_rsci_oswt(chn_mul_op_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_mul_op_rsci_iswt0(chn_mul_op_rsci_iswt0),
      .chn_mul_op_rsci_ld_core_psct(chn_mul_op_rsci_ld_core_psct),
      .chn_mul_op_rsci_biwt(chn_mul_op_rsci_biwt),
      .chn_mul_op_rsci_bdwt(chn_mul_op_rsci_bdwt),
      .chn_mul_op_rsci_ld_core_sct(chn_mul_op_rsci_ld_core_sct),
      .chn_mul_op_rsci_vd(chn_mul_op_rsci_vd)
    );
  SDP_X_X_mul_core_chn_mul_op_rsci_chn_mul_op_wait_dp X_mul_core_chn_mul_op_rsci_chn_mul_op_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_op_rsci_oswt(chn_mul_op_rsci_oswt),
      .chn_mul_op_rsci_bawt(chn_mul_op_rsci_bawt),
      .chn_mul_op_rsci_wen_comp(chn_mul_op_rsci_wen_comp),
      .chn_mul_op_rsci_d_mxwt(chn_mul_op_rsci_d_mxwt),
      .chn_mul_op_rsci_biwt(chn_mul_op_rsci_biwt),
      .chn_mul_op_rsci_bdwt(chn_mul_op_rsci_bdwt),
      .chn_mul_op_rsci_d(chn_mul_op_rsci_d)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core_chn_mul_in_rsci
// ------------------------------------------------------------------
module SDP_X_X_mul_core_chn_mul_in_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_in_rsc_slz, chn_mul_in_rsc_sz, chn_mul_in_rsc_z,
      chn_mul_in_rsc_vz, chn_mul_in_rsc_lz, chn_mul_in_rsci_oswt, core_wen, chn_mul_in_rsci_iswt0,
      chn_mul_in_rsci_bawt, chn_mul_in_rsci_wen_comp, chn_mul_in_rsci_ld_core_psct,
      chn_mul_in_rsci_d_mxwt, core_wten
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output chn_mul_in_rsc_slz;
  input chn_mul_in_rsc_sz;
  input [527:0] chn_mul_in_rsc_z;
  input chn_mul_in_rsc_vz;
  output chn_mul_in_rsc_lz;
  input chn_mul_in_rsci_oswt;
  input core_wen;
  input chn_mul_in_rsci_iswt0;
  output chn_mul_in_rsci_bawt;
  output chn_mul_in_rsci_wen_comp;
  input chn_mul_in_rsci_ld_core_psct;
  output [527:0] chn_mul_in_rsci_d_mxwt;
  input core_wten;
// Interconnect Declarations
  wire chn_mul_in_rsci_biwt;
  wire chn_mul_in_rsci_bdwt;
  wire chn_mul_in_rsci_ld_core_sct;
  wire chn_mul_in_rsci_vd;
  wire [527:0] chn_mul_in_rsci_d;
  wire chn_mul_in_rsci_sd;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_chan_in_v2 #(.rscid(32'sd14),
  .width(32'sd528),
  .sz_width(32'sd1)) chn_mul_in_rsci (
      .ld(chn_mul_in_rsci_ld_core_sct),
      .vd(chn_mul_in_rsci_vd),
      .d(chn_mul_in_rsci_d),
      .lz(chn_mul_in_rsc_lz),
      .vz(chn_mul_in_rsc_vz),
      .z(chn_mul_in_rsc_z),
      .sd(chn_mul_in_rsci_sd),
      .sld(1'b0),
      .sz(chn_mul_in_rsc_sz),
      .slz(chn_mul_in_rsc_slz)
    );
  SDP_X_X_mul_core_chn_mul_in_rsci_chn_mul_in_wait_ctrl X_mul_core_chn_mul_in_rsci_chn_mul_in_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_in_rsci_oswt(chn_mul_in_rsci_oswt),
      .core_wen(core_wen),
      .chn_mul_in_rsci_iswt0(chn_mul_in_rsci_iswt0),
      .chn_mul_in_rsci_ld_core_psct(chn_mul_in_rsci_ld_core_psct),
      .core_wten(core_wten),
      .chn_mul_in_rsci_biwt(chn_mul_in_rsci_biwt),
      .chn_mul_in_rsci_bdwt(chn_mul_in_rsci_bdwt),
      .chn_mul_in_rsci_ld_core_sct(chn_mul_in_rsci_ld_core_sct),
      .chn_mul_in_rsci_vd(chn_mul_in_rsci_vd)
    );
  SDP_X_X_mul_core_chn_mul_in_rsci_chn_mul_in_wait_dp X_mul_core_chn_mul_in_rsci_chn_mul_in_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_in_rsci_oswt(chn_mul_in_rsci_oswt),
      .chn_mul_in_rsci_bawt(chn_mul_in_rsci_bawt),
      .chn_mul_in_rsci_wen_comp(chn_mul_in_rsci_wen_comp),
      .chn_mul_in_rsci_d_mxwt(chn_mul_in_rsci_d_mxwt),
      .chn_mul_in_rsci_biwt(chn_mul_in_rsci_biwt),
      .chn_mul_in_rsci_bdwt(chn_mul_in_rsci_bdwt),
      .chn_mul_in_rsci_d(chn_mul_in_rsci_d)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_trt_core_cfg_mul_shift_value_rsc_triosy_obj
// ------------------------------------------------------------------
module SDP_X_X_trt_core_cfg_mul_shift_value_rsc_triosy_obj (
  nvdla_core_clk, nvdla_core_rstn, cfg_mul_shift_value_rsc_triosy_lz, cfg_mul_shift_value_rsc_triosy_obj_oswt,
      core_wen, core_wten, cfg_mul_shift_value_rsc_triosy_obj_iswt0, cfg_mul_shift_value_rsc_triosy_obj_bawt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_mul_shift_value_rsc_triosy_lz;
  input cfg_mul_shift_value_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_mul_shift_value_rsc_triosy_obj_iswt0;
  output cfg_mul_shift_value_rsc_triosy_obj_bawt;
// Interconnect Declarations
  wire cfg_mul_shift_value_rsc_triosy_obj_biwt;
  wire cfg_mul_shift_value_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_io_sync_v1 #(.valid(32'sd0)) cfg_mul_shift_value_rsc_triosy_obj (
      .ld(cfg_mul_shift_value_rsc_triosy_obj_biwt),
      .lz(cfg_mul_shift_value_rsc_triosy_lz)
    );
  SDP_X_X_trt_core_cfg_mul_shift_value_rsc_triosy_obj_cfg_mul_shift_value_rsc_triosy_wait_ctrl
      X_trt_core_cfg_mul_shift_value_rsc_triosy_obj_cfg_mul_shift_value_rsc_triosy_wait_ctrl_inst
      (
      .cfg_mul_shift_value_rsc_triosy_obj_oswt(cfg_mul_shift_value_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_mul_shift_value_rsc_triosy_obj_iswt0(cfg_mul_shift_value_rsc_triosy_obj_iswt0),
      .cfg_mul_shift_value_rsc_triosy_obj_biwt(cfg_mul_shift_value_rsc_triosy_obj_biwt),
      .cfg_mul_shift_value_rsc_triosy_obj_bdwt(cfg_mul_shift_value_rsc_triosy_obj_bdwt)
    );
  SDP_X_X_trt_core_cfg_mul_shift_value_rsc_triosy_obj_cfg_mul_shift_value_rsc_triosy_wait_dp
      X_trt_core_cfg_mul_shift_value_rsc_triosy_obj_cfg_mul_shift_value_rsc_triosy_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_mul_shift_value_rsc_triosy_obj_bawt(cfg_mul_shift_value_rsc_triosy_obj_bawt),
      .cfg_mul_shift_value_rsc_triosy_obj_biwt(cfg_mul_shift_value_rsc_triosy_obj_biwt),
      .cfg_mul_shift_value_rsc_triosy_obj_bdwt(cfg_mul_shift_value_rsc_triosy_obj_bdwt)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_trt_core_chn_trt_out_rsci
// ------------------------------------------------------------------
module SDP_X_X_trt_core_chn_trt_out_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_trt_out_rsc_z, chn_trt_out_rsc_vz, chn_trt_out_rsc_lz,
      chn_trt_out_rsci_oswt, core_wen, core_wten, chn_trt_out_rsci_iswt0, chn_trt_out_rsci_bawt,
      chn_trt_out_rsci_wen_comp, chn_trt_out_rsci_ld_core_psct, chn_trt_out_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output [511:0] chn_trt_out_rsc_z;
  input chn_trt_out_rsc_vz;
  output chn_trt_out_rsc_lz;
  input chn_trt_out_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_trt_out_rsci_iswt0;
  output chn_trt_out_rsci_bawt;
  output chn_trt_out_rsci_wen_comp;
  input chn_trt_out_rsci_ld_core_psct;
  input [511:0] chn_trt_out_rsci_d;
// Interconnect Declarations
  wire chn_trt_out_rsci_biwt;
  wire chn_trt_out_rsci_bdwt;
  wire chn_trt_out_rsci_ld_core_sct;
  wire chn_trt_out_rsci_vd;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_out_stdreg_wait_v1 #(.rscid(32'sd31),
  .width(32'sd512)) chn_trt_out_rsci (
      .ld(chn_trt_out_rsci_ld_core_sct),
      .vd(chn_trt_out_rsci_vd),
      .d(chn_trt_out_rsci_d),
      .lz(chn_trt_out_rsc_lz),
      .vz(chn_trt_out_rsc_vz),
      .z(chn_trt_out_rsc_z)
    );
  SDP_X_X_trt_core_chn_trt_out_rsci_chn_trt_out_wait_ctrl X_trt_core_chn_trt_out_rsci_chn_trt_out_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_trt_out_rsci_oswt(chn_trt_out_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_trt_out_rsci_iswt0(chn_trt_out_rsci_iswt0),
      .chn_trt_out_rsci_ld_core_psct(chn_trt_out_rsci_ld_core_psct),
      .chn_trt_out_rsci_biwt(chn_trt_out_rsci_biwt),
      .chn_trt_out_rsci_bdwt(chn_trt_out_rsci_bdwt),
      .chn_trt_out_rsci_ld_core_sct(chn_trt_out_rsci_ld_core_sct),
      .chn_trt_out_rsci_vd(chn_trt_out_rsci_vd)
    );
  SDP_X_X_trt_core_chn_trt_out_rsci_chn_trt_out_wait_dp X_trt_core_chn_trt_out_rsci_chn_trt_out_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_trt_out_rsci_oswt(chn_trt_out_rsci_oswt),
      .chn_trt_out_rsci_bawt(chn_trt_out_rsci_bawt),
      .chn_trt_out_rsci_wen_comp(chn_trt_out_rsci_wen_comp),
      .chn_trt_out_rsci_biwt(chn_trt_out_rsci_biwt),
      .chn_trt_out_rsci_bdwt(chn_trt_out_rsci_bdwt)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_trt_core_chn_trt_in_rsci
// ------------------------------------------------------------------
module SDP_X_X_trt_core_chn_trt_in_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_trt_in_rsc_slz, chn_trt_in_rsc_sz, chn_trt_in_rsc_z,
      chn_trt_in_rsc_vz, chn_trt_in_rsc_lz, chn_trt_in_rsci_oswt, core_wen, chn_trt_in_rsci_iswt0,
      chn_trt_in_rsci_bawt, chn_trt_in_rsci_wen_comp, chn_trt_in_rsci_ld_core_psct,
      chn_trt_in_rsci_d_mxwt, core_wten
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output chn_trt_in_rsc_slz;
  input chn_trt_in_rsc_sz;
  input [799:0] chn_trt_in_rsc_z;
  input chn_trt_in_rsc_vz;
  output chn_trt_in_rsc_lz;
  input chn_trt_in_rsci_oswt;
  input core_wen;
  input chn_trt_in_rsci_iswt0;
  output chn_trt_in_rsci_bawt;
  output chn_trt_in_rsci_wen_comp;
  input chn_trt_in_rsci_ld_core_psct;
  output [799:0] chn_trt_in_rsci_d_mxwt;
  input core_wten;
// Interconnect Declarations
  wire chn_trt_in_rsci_biwt;
  wire chn_trt_in_rsci_bdwt;
  wire chn_trt_in_rsci_ld_core_sct;
  wire chn_trt_in_rsci_vd;
  wire [799:0] chn_trt_in_rsci_d;
  wire chn_trt_in_rsci_sd;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_chan_in_v2 #(.rscid(32'sd27),
  .width(32'sd800),
  .sz_width(32'sd1)) chn_trt_in_rsci (
      .ld(chn_trt_in_rsci_ld_core_sct),
      .vd(chn_trt_in_rsci_vd),
      .d(chn_trt_in_rsci_d),
      .lz(chn_trt_in_rsc_lz),
      .vz(chn_trt_in_rsc_vz),
      .z(chn_trt_in_rsc_z),
      .sd(chn_trt_in_rsci_sd),
      .sld(1'b0),
      .sz(chn_trt_in_rsc_sz),
      .slz(chn_trt_in_rsc_slz)
    );
  SDP_X_X_trt_core_chn_trt_in_rsci_chn_trt_in_wait_ctrl X_trt_core_chn_trt_in_rsci_chn_trt_in_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_trt_in_rsci_oswt(chn_trt_in_rsci_oswt),
      .core_wen(core_wen),
      .chn_trt_in_rsci_iswt0(chn_trt_in_rsci_iswt0),
      .chn_trt_in_rsci_ld_core_psct(chn_trt_in_rsci_ld_core_psct),
      .core_wten(core_wten),
      .chn_trt_in_rsci_biwt(chn_trt_in_rsci_biwt),
      .chn_trt_in_rsci_bdwt(chn_trt_in_rsci_bdwt),
      .chn_trt_in_rsci_ld_core_sct(chn_trt_in_rsci_ld_core_sct),
      .chn_trt_in_rsci_vd(chn_trt_in_rsci_vd)
    );
  SDP_X_X_trt_core_chn_trt_in_rsci_chn_trt_in_wait_dp X_trt_core_chn_trt_in_rsci_chn_trt_in_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_trt_in_rsci_oswt(chn_trt_in_rsci_oswt),
      .chn_trt_in_rsci_bawt(chn_trt_in_rsci_bawt),
      .chn_trt_in_rsci_wen_comp(chn_trt_in_rsci_wen_comp),
      .chn_trt_in_rsci_d_mxwt(chn_trt_in_rsci_d_mxwt),
      .chn_trt_in_rsci_biwt(chn_trt_in_rsci_biwt),
      .chn_trt_in_rsci_bdwt(chn_trt_in_rsci_bdwt),
      .chn_trt_in_rsci_d(chn_trt_in_rsci_d)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_relu_core_cfg_relu_bypass_rsc_triosy_obj
// ------------------------------------------------------------------
module SDP_X_X_relu_core_cfg_relu_bypass_rsc_triosy_obj (
  nvdla_core_clk, nvdla_core_rstn, cfg_relu_bypass_rsc_triosy_lz, cfg_relu_bypass_rsc_triosy_obj_oswt,
      core_wen, core_wten, cfg_relu_bypass_rsc_triosy_obj_iswt0, cfg_relu_bypass_rsc_triosy_obj_bawt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_relu_bypass_rsc_triosy_lz;
  input cfg_relu_bypass_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_relu_bypass_rsc_triosy_obj_iswt0;
  output cfg_relu_bypass_rsc_triosy_obj_bawt;
// Interconnect Declarations
  wire cfg_relu_bypass_rsc_triosy_obj_biwt;
  wire cfg_relu_bypass_rsc_triosy_obj_bdwt;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_io_sync_v1 #(.valid(32'sd0)) cfg_relu_bypass_rsc_triosy_obj (
      .ld(cfg_relu_bypass_rsc_triosy_obj_biwt),
      .lz(cfg_relu_bypass_rsc_triosy_lz)
    );
  SDP_X_X_relu_core_cfg_relu_bypass_rsc_triosy_obj_cfg_relu_bypass_rsc_triosy_wait_ctrl
      X_relu_core_cfg_relu_bypass_rsc_triosy_obj_cfg_relu_bypass_rsc_triosy_wait_ctrl_inst
      (
      .cfg_relu_bypass_rsc_triosy_obj_oswt(cfg_relu_bypass_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_relu_bypass_rsc_triosy_obj_iswt0(cfg_relu_bypass_rsc_triosy_obj_iswt0),
      .cfg_relu_bypass_rsc_triosy_obj_biwt(cfg_relu_bypass_rsc_triosy_obj_biwt),
      .cfg_relu_bypass_rsc_triosy_obj_bdwt(cfg_relu_bypass_rsc_triosy_obj_bdwt)
    );
  SDP_X_X_relu_core_cfg_relu_bypass_rsc_triosy_obj_cfg_relu_bypass_rsc_triosy_wait_dp X_relu_core_cfg_relu_bypass_rsc_triosy_obj_cfg_relu_bypass_rsc_triosy_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_relu_bypass_rsc_triosy_obj_bawt(cfg_relu_bypass_rsc_triosy_obj_bawt),
      .cfg_relu_bypass_rsc_triosy_obj_biwt(cfg_relu_bypass_rsc_triosy_obj_biwt),
      .cfg_relu_bypass_rsc_triosy_obj_bdwt(cfg_relu_bypass_rsc_triosy_obj_bdwt)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_relu_core_chn_relu_out_rsci
// ------------------------------------------------------------------
module SDP_X_X_relu_core_chn_relu_out_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_relu_out_rsc_z, chn_relu_out_rsc_vz, chn_relu_out_rsc_lz,
      chn_relu_out_rsci_oswt, core_wen, core_wten, chn_relu_out_rsci_iswt0, chn_relu_out_rsci_bawt,
      chn_relu_out_rsci_wen_comp, chn_relu_out_rsci_ld_core_psct, chn_relu_out_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output [511:0] chn_relu_out_rsc_z;
  input chn_relu_out_rsc_vz;
  output chn_relu_out_rsc_lz;
  input chn_relu_out_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_relu_out_rsci_iswt0;
  output chn_relu_out_rsci_bawt;
  output chn_relu_out_rsci_wen_comp;
  input chn_relu_out_rsci_ld_core_psct;
  input [511:0] chn_relu_out_rsci_d;
// Interconnect Declarations
  wire chn_relu_out_rsci_biwt;
  wire chn_relu_out_rsci_bdwt;
  wire chn_relu_out_rsci_ld_core_sct;
  wire chn_relu_out_rsci_vd;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_out_stdreg_wait_v1 #(.rscid(32'sd36),
  .width(32'sd512)) chn_relu_out_rsci (
      .ld(chn_relu_out_rsci_ld_core_sct),
      .vd(chn_relu_out_rsci_vd),
      .d(chn_relu_out_rsci_d),
      .lz(chn_relu_out_rsc_lz),
      .vz(chn_relu_out_rsc_vz),
      .z(chn_relu_out_rsc_z)
    );
  SDP_X_X_relu_core_chn_relu_out_rsci_chn_relu_out_wait_ctrl X_relu_core_chn_relu_out_rsci_chn_relu_out_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_relu_out_rsci_oswt(chn_relu_out_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_relu_out_rsci_iswt0(chn_relu_out_rsci_iswt0),
      .chn_relu_out_rsci_ld_core_psct(chn_relu_out_rsci_ld_core_psct),
      .chn_relu_out_rsci_biwt(chn_relu_out_rsci_biwt),
      .chn_relu_out_rsci_bdwt(chn_relu_out_rsci_bdwt),
      .chn_relu_out_rsci_ld_core_sct(chn_relu_out_rsci_ld_core_sct),
      .chn_relu_out_rsci_vd(chn_relu_out_rsci_vd)
    );
  SDP_X_X_relu_core_chn_relu_out_rsci_chn_relu_out_wait_dp X_relu_core_chn_relu_out_rsci_chn_relu_out_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_relu_out_rsci_oswt(chn_relu_out_rsci_oswt),
      .chn_relu_out_rsci_bawt(chn_relu_out_rsci_bawt),
      .chn_relu_out_rsci_wen_comp(chn_relu_out_rsci_wen_comp),
      .chn_relu_out_rsci_biwt(chn_relu_out_rsci_biwt),
      .chn_relu_out_rsci_bdwt(chn_relu_out_rsci_bdwt)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_relu_core_chn_relu_in_rsci
// ------------------------------------------------------------------
module SDP_X_X_relu_core_chn_relu_in_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_relu_in_rsc_z, chn_relu_in_rsc_vz, chn_relu_in_rsc_lz,
      chn_relu_in_rsci_oswt, core_wen, chn_relu_in_rsci_iswt0, chn_relu_in_rsci_bawt,
      chn_relu_in_rsci_wen_comp, chn_relu_in_rsci_ld_core_psct, chn_relu_in_rsci_d_mxwt,
      core_wten
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [511:0] chn_relu_in_rsc_z;
  input chn_relu_in_rsc_vz;
  output chn_relu_in_rsc_lz;
  input chn_relu_in_rsci_oswt;
  input core_wen;
  input chn_relu_in_rsci_iswt0;
  output chn_relu_in_rsci_bawt;
  output chn_relu_in_rsci_wen_comp;
  input chn_relu_in_rsci_ld_core_psct;
  output [511:0] chn_relu_in_rsci_d_mxwt;
  input core_wten;
// Interconnect Declarations
  wire chn_relu_in_rsci_biwt;
  wire chn_relu_in_rsci_bdwt;
  wire chn_relu_in_rsci_ld_core_sct;
  wire chn_relu_in_rsci_vd;
  wire [511:0] chn_relu_in_rsci_d;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_in_wire_wait_v1 #(.rscid(32'sd33),
  .width(32'sd512)) chn_relu_in_rsci (
      .ld(chn_relu_in_rsci_ld_core_sct),
      .vd(chn_relu_in_rsci_vd),
      .d(chn_relu_in_rsci_d),
      .lz(chn_relu_in_rsc_lz),
      .vz(chn_relu_in_rsc_vz),
      .z(chn_relu_in_rsc_z)
    );
  SDP_X_X_relu_core_chn_relu_in_rsci_chn_relu_in_wait_ctrl X_relu_core_chn_relu_in_rsci_chn_relu_in_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_relu_in_rsci_oswt(chn_relu_in_rsci_oswt),
      .core_wen(core_wen),
      .chn_relu_in_rsci_iswt0(chn_relu_in_rsci_iswt0),
      .chn_relu_in_rsci_ld_core_psct(chn_relu_in_rsci_ld_core_psct),
      .core_wten(core_wten),
      .chn_relu_in_rsci_biwt(chn_relu_in_rsci_biwt),
      .chn_relu_in_rsci_bdwt(chn_relu_in_rsci_bdwt),
      .chn_relu_in_rsci_ld_core_sct(chn_relu_in_rsci_ld_core_sct),
      .chn_relu_in_rsci_vd(chn_relu_in_rsci_vd)
    );
  SDP_X_X_relu_core_chn_relu_in_rsci_chn_relu_in_wait_dp X_relu_core_chn_relu_in_rsci_chn_relu_in_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_relu_in_rsci_oswt(chn_relu_in_rsci_oswt),
      .chn_relu_in_rsci_bawt(chn_relu_in_rsci_bawt),
      .chn_relu_in_rsci_wen_comp(chn_relu_in_rsci_wen_comp),
      .chn_relu_in_rsci_d_mxwt(chn_relu_in_rsci_d_mxwt),
      .chn_relu_in_rsci_biwt(chn_relu_in_rsci_biwt),
      .chn_relu_in_rsci_bdwt(chn_relu_in_rsci_bdwt),
      .chn_relu_in_rsci_d(chn_relu_in_rsci_d)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu_core
// ------------------------------------------------------------------
module SDP_X_X_alu_core (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_in_rsc_z, chn_alu_in_rsc_vz, chn_alu_in_rsc_lz,
      chn_alu_op_rsc_z, chn_alu_op_rsc_vz, chn_alu_op_rsc_lz, cfg_alu_op_rsc_triosy_lz,
      cfg_alu_bypass_rsc_triosy_lz, cfg_alu_algo_rsc_triosy_lz, cfg_alu_src_rsc_triosy_lz,
      cfg_alu_shift_value_rsc_triosy_lz, cfg_nan_to_zero, cfg_precision, chn_alu_out_rsc_z,
      chn_alu_out_rsc_vz, chn_alu_out_rsc_lz, chn_alu_in_rsci_oswt, chn_alu_in_rsci_oswt_unreg,
      chn_alu_op_rsci_oswt, chn_alu_op_rsci_oswt_unreg, cfg_alu_op_rsci_d, cfg_alu_bypass_rsci_d,
      cfg_alu_algo_rsci_d, cfg_alu_src_rsci_d, cfg_alu_shift_value_rsci_d, chn_alu_out_rsci_oswt,
      chn_alu_out_rsci_oswt_unreg, cfg_alu_op_rsc_triosy_obj_oswt, cfg_alu_bypass_rsc_triosy_obj_oswt,
      cfg_alu_algo_rsc_triosy_obj_oswt, cfg_alu_src_rsc_triosy_obj_oswt, cfg_alu_shift_value_rsc_triosy_obj_oswt,
      cfg_alu_op_rsc_triosy_obj_oswt_unreg_pff
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [511:0] chn_alu_in_rsc_z;
  input chn_alu_in_rsc_vz;
  output chn_alu_in_rsc_lz;
  input [255:0] chn_alu_op_rsc_z;
  input chn_alu_op_rsc_vz;
  output chn_alu_op_rsc_lz;
  output cfg_alu_op_rsc_triosy_lz;
  output cfg_alu_bypass_rsc_triosy_lz;
  output cfg_alu_algo_rsc_triosy_lz;
  output cfg_alu_src_rsc_triosy_lz;
  output cfg_alu_shift_value_rsc_triosy_lz;
  input cfg_nan_to_zero;
  input [1:0] cfg_precision;
  output [527:0] chn_alu_out_rsc_z;
  input chn_alu_out_rsc_vz;
  output chn_alu_out_rsc_lz;
  input chn_alu_in_rsci_oswt;
  output chn_alu_in_rsci_oswt_unreg;
  input chn_alu_op_rsci_oswt;
  output chn_alu_op_rsci_oswt_unreg;
  input [15:0] cfg_alu_op_rsci_d;
  input cfg_alu_bypass_rsci_d;
  input [1:0] cfg_alu_algo_rsci_d;
  input cfg_alu_src_rsci_d;
  input [5:0] cfg_alu_shift_value_rsci_d;
  input chn_alu_out_rsci_oswt;
  output chn_alu_out_rsci_oswt_unreg;
  input cfg_alu_op_rsc_triosy_obj_oswt;
  input cfg_alu_bypass_rsc_triosy_obj_oswt;
  input cfg_alu_algo_rsc_triosy_obj_oswt;
  input cfg_alu_src_rsc_triosy_obj_oswt;
  input cfg_alu_shift_value_rsc_triosy_obj_oswt;
  output cfg_alu_op_rsc_triosy_obj_oswt_unreg_pff;
// Interconnect Declarations
  wire core_wen;
  reg chn_alu_in_rsci_iswt0;
  wire chn_alu_in_rsci_bawt;
  wire chn_alu_in_rsci_wen_comp;
  reg chn_alu_in_rsci_ld_core_psct;
  wire [511:0] chn_alu_in_rsci_d_mxwt;
  wire core_wten;
  reg chn_alu_op_rsci_iswt0;
  wire chn_alu_op_rsci_bawt;
  wire chn_alu_op_rsci_wen_comp;
  reg chn_alu_op_rsci_ld_core_psct;
  wire [255:0] chn_alu_op_rsci_d_mxwt;
  reg chn_alu_out_rsci_iswt0;
  wire chn_alu_out_rsci_bawt;
  wire chn_alu_out_rsci_wen_comp;
  wire cfg_alu_op_rsc_triosy_obj_bawt;
  wire cfg_alu_bypass_rsc_triosy_obj_bawt;
  wire cfg_alu_algo_rsc_triosy_obj_bawt;
  wire cfg_alu_src_rsc_triosy_obj_bawt;
  wire cfg_alu_shift_value_rsc_triosy_obj_bawt;
  reg [1:0] chn_alu_out_rsci_d_527_526;
  reg [3:0] chn_alu_out_rsci_d_525_522;
  reg [3:0] chn_alu_out_rsci_d_521_518;
  reg [21:0] chn_alu_out_rsci_d_517_496;
  reg chn_alu_out_rsci_d_495;
  reg [1:0] chn_alu_out_rsci_d_494_493;
  reg [3:0] chn_alu_out_rsci_d_492_489;
  reg [3:0] chn_alu_out_rsci_d_488_485;
  reg [21:0] chn_alu_out_rsci_d_484_463;
  reg chn_alu_out_rsci_d_462;
  reg [1:0] chn_alu_out_rsci_d_461_460;
  reg [3:0] chn_alu_out_rsci_d_459_456;
  reg [3:0] chn_alu_out_rsci_d_455_452;
  reg [21:0] chn_alu_out_rsci_d_451_430;
  reg chn_alu_out_rsci_d_429;
  reg [1:0] chn_alu_out_rsci_d_428_427;
  reg [3:0] chn_alu_out_rsci_d_426_423;
  reg [3:0] chn_alu_out_rsci_d_422_419;
  reg [21:0] chn_alu_out_rsci_d_418_397;
  reg chn_alu_out_rsci_d_396;
  reg [1:0] chn_alu_out_rsci_d_395_394;
  reg [3:0] chn_alu_out_rsci_d_393_390;
  reg [3:0] chn_alu_out_rsci_d_389_386;
  reg [21:0] chn_alu_out_rsci_d_385_364;
  reg chn_alu_out_rsci_d_363;
  reg [1:0] chn_alu_out_rsci_d_362_361;
  reg [3:0] chn_alu_out_rsci_d_360_357;
  reg [3:0] chn_alu_out_rsci_d_356_353;
  reg [21:0] chn_alu_out_rsci_d_352_331;
  reg chn_alu_out_rsci_d_330;
  reg [1:0] chn_alu_out_rsci_d_329_328;
  reg [3:0] chn_alu_out_rsci_d_327_324;
  reg [3:0] chn_alu_out_rsci_d_323_320;
  reg [21:0] chn_alu_out_rsci_d_319_298;
  reg chn_alu_out_rsci_d_297;
  reg [1:0] chn_alu_out_rsci_d_296_295;
  reg [3:0] chn_alu_out_rsci_d_294_291;
  reg [3:0] chn_alu_out_rsci_d_290_287;
  reg [21:0] chn_alu_out_rsci_d_286_265;
  reg chn_alu_out_rsci_d_264;
  reg [1:0] chn_alu_out_rsci_d_263_262;
  reg [3:0] chn_alu_out_rsci_d_261_258;
  reg [3:0] chn_alu_out_rsci_d_257_254;
  reg [21:0] chn_alu_out_rsci_d_253_232;
  reg chn_alu_out_rsci_d_231;
  reg [1:0] chn_alu_out_rsci_d_230_229;
  reg [3:0] chn_alu_out_rsci_d_228_225;
  reg [3:0] chn_alu_out_rsci_d_224_221;
  reg [21:0] chn_alu_out_rsci_d_220_199;
  reg chn_alu_out_rsci_d_198;
  reg [1:0] chn_alu_out_rsci_d_197_196;
  reg [3:0] chn_alu_out_rsci_d_195_192;
  reg [3:0] chn_alu_out_rsci_d_191_188;
  reg [21:0] chn_alu_out_rsci_d_187_166;
  reg chn_alu_out_rsci_d_165;
  reg [1:0] chn_alu_out_rsci_d_164_163;
  reg [3:0] chn_alu_out_rsci_d_162_159;
  reg [3:0] chn_alu_out_rsci_d_158_155;
  reg [21:0] chn_alu_out_rsci_d_154_133;
  reg chn_alu_out_rsci_d_132;
  reg [1:0] chn_alu_out_rsci_d_131_130;
  reg [3:0] chn_alu_out_rsci_d_129_126;
  reg [3:0] chn_alu_out_rsci_d_125_122;
  reg [21:0] chn_alu_out_rsci_d_121_100;
  reg chn_alu_out_rsci_d_99;
  reg [1:0] chn_alu_out_rsci_d_98_97;
  reg [3:0] chn_alu_out_rsci_d_96_93;
  reg [3:0] chn_alu_out_rsci_d_92_89;
  reg [21:0] chn_alu_out_rsci_d_88_67;
  reg chn_alu_out_rsci_d_66;
  reg [1:0] chn_alu_out_rsci_d_65_64;
  reg [3:0] chn_alu_out_rsci_d_63_60;
  reg [3:0] chn_alu_out_rsci_d_59_56;
  reg [21:0] chn_alu_out_rsci_d_55_34;
  reg chn_alu_out_rsci_d_33;
  reg [1:0] chn_alu_out_rsci_d_32_31;
  reg [3:0] chn_alu_out_rsci_d_30_27;
  reg [3:0] chn_alu_out_rsci_d_26_23;
  reg [21:0] chn_alu_out_rsci_d_22_1;
  reg chn_alu_out_rsci_d_0;
  wire [1:0] fsm_output;
  wire and_91_tmp;
  wire IsNaN_5U_23U_nor_15_tmp;
  wire IsNaN_5U_23U_nor_14_tmp;
  wire IsNaN_5U_23U_nor_13_tmp;
  wire IsNaN_5U_23U_nor_12_tmp;
  wire IsNaN_5U_23U_nor_11_tmp;
  wire IsNaN_5U_23U_nor_10_tmp;
  wire IsNaN_5U_23U_nor_9_tmp;
  wire IsNaN_5U_23U_nor_8_tmp;
  wire IsNaN_5U_23U_nor_7_tmp;
  wire IsNaN_5U_23U_nor_6_tmp;
  wire IsNaN_5U_23U_nor_5_tmp;
  wire IsNaN_5U_23U_nor_4_tmp;
  wire IsNaN_5U_23U_nor_3_tmp;
  wire IsNaN_5U_23U_nor_2_tmp;
  wire IsNaN_5U_23U_nor_1_tmp;
  wire IsNaN_5U_23U_nor_tmp;
  wire IsNaN_5U_10U_nor_15_tmp;
  wire IsNaN_5U_10U_nor_14_tmp;
  wire IsNaN_5U_10U_nor_13_tmp;
  wire IsNaN_5U_10U_nor_12_tmp;
  wire IsNaN_5U_10U_nor_11_tmp;
  wire IsNaN_5U_10U_nor_10_tmp;
  wire IsNaN_5U_10U_nor_9_tmp;
  wire IsNaN_5U_10U_nor_8_tmp;
  wire IsNaN_5U_10U_nor_7_tmp;
  wire IsNaN_5U_10U_nor_6_tmp;
  wire IsNaN_5U_10U_nor_5_tmp;
  wire IsNaN_5U_10U_nor_4_tmp;
  wire IsNaN_5U_10U_nor_3_tmp;
  wire IsNaN_5U_10U_nor_2_tmp;
  wire IsNaN_5U_10U_nor_1_tmp;
  wire IsNaN_5U_10U_nor_tmp;
  wire [4:0] else_mux_47_tmp;
  wire [4:0] else_mux_44_tmp;
  wire [4:0] else_mux_41_tmp;
  wire [4:0] else_mux_38_tmp;
  wire [4:0] else_mux_35_tmp;
  wire [4:0] else_mux_32_tmp;
  wire [4:0] else_mux_29_tmp;
  wire [4:0] else_mux_26_tmp;
  wire [4:0] else_mux_23_tmp;
  wire [4:0] else_mux_20_tmp;
  wire [4:0] else_mux_17_tmp;
  wire [4:0] else_mux_14_tmp;
  wire [4:0] else_mux_11_tmp;
  wire [4:0] else_mux_8_tmp;
  wire [4:0] else_mux_5_tmp;
  wire [4:0] else_mux_2_tmp;
  wire and_89_tmp;
  wire alu_loop_op_16_FpMantRNE_49U_24U_else_and_1_tmp;
  wire alu_loop_op_15_FpMantRNE_49U_24U_else_and_tmp;
  wire alu_loop_op_14_FpMantRNE_49U_24U_else_and_1_tmp;
  wire alu_loop_op_13_FpMantRNE_49U_24U_else_and_tmp;
  wire alu_loop_op_12_FpMantRNE_49U_24U_else_and_1_tmp;
  wire alu_loop_op_11_FpMantRNE_49U_24U_else_and_tmp;
  wire alu_loop_op_10_FpMantRNE_49U_24U_else_and_1_tmp;
  wire alu_loop_op_9_FpMantRNE_49U_24U_else_and_tmp;
  wire alu_loop_op_8_FpMantRNE_49U_24U_else_and_1_tmp;
  wire alu_loop_op_7_FpMantRNE_49U_24U_else_and_tmp;
  wire alu_loop_op_6_FpMantRNE_49U_24U_else_and_1_tmp;
  wire alu_loop_op_5_FpMantRNE_49U_24U_else_and_tmp;
  wire alu_loop_op_4_FpMantRNE_49U_24U_else_and_1_tmp;
  wire alu_loop_op_3_FpMantRNE_49U_24U_else_and_tmp;
  wire alu_loop_op_2_FpMantRNE_49U_24U_else_and_1_tmp;
  wire alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp;
  wire not_tmp_4;
  wire or_tmp_20;
  wire or_tmp_24;
  wire or_tmp_39;
  wire or_tmp_55;
  wire or_tmp_76;
  wire or_tmp_97;
  wire or_tmp_263;
  wire or_tmp_327;
  wire or_tmp_329;
  wire mux_tmp_149;
  wire not_tmp_79;
  wire mux_tmp_156;
  wire or_tmp_670;
  wire mux_tmp_339;
  wire mux_tmp_392;
  wire mux_tmp_393;
  wire or_tmp_1848;
  wire or_tmp_1857;
  wire mux_tmp_778;
  wire mux_tmp_779;
  wire or_tmp_1865;
  wire mux_tmp_781;
  wire or_tmp_1868;
  wire mux_tmp_782;
  wire mux_tmp_783;
  wire mux_tmp_785;
  wire mux_tmp_786;
  wire mux_tmp_787;
  wire mux_tmp_788;
  wire mux_tmp_789;
  wire mux_tmp_790;
  wire mux_tmp_791;
  wire mux_tmp_792;
  wire mux_tmp_793;
  wire mux_tmp_795;
  wire mux_tmp_796;
  wire or_tmp_1915;
  wire mux_tmp_823;
  wire mux_tmp_1077;
  wire or_tmp_2842;
  wire and_dcpl_7;
  wire and_dcpl_8;
  wire and_dcpl_10;
  wire and_dcpl_11;
  wire or_dcpl_3;
  wire and_dcpl_14;
  wire and_dcpl_21;
  wire and_dcpl_22;
  wire and_dcpl_23;
  wire and_dcpl_28;
  wire and_dcpl_29;
  wire or_dcpl_13;
  wire or_dcpl_14;
  wire and_dcpl_30;
  wire and_dcpl_34;
  wire and_dcpl_36;
  wire and_dcpl_122;
  wire and_dcpl_126;
  wire and_dcpl_127;
  wire and_dcpl_241;
  wire and_dcpl_256;
  wire and_dcpl_263;
  wire and_dcpl_294;
  wire and_dcpl_309;
  wire and_dcpl_316;
  wire and_dcpl_347;
  wire and_dcpl_354;
  wire and_dcpl_361;
  wire or_dcpl_112;
  wire and_dcpl_369;
  wire or_dcpl_113;
  wire and_dcpl_372;
  wire or_dcpl_116;
  wire and_dcpl_375;
  wire and_dcpl_379;
  wire and_dcpl_394;
  wire and_dcpl_395;
  wire and_dcpl_397;
  wire and_dcpl_398;
  wire and_dcpl_401;
  wire and_dcpl_402;
  wire and_dcpl_404;
  wire and_dcpl_406;
  wire and_dcpl_407;
  wire or_dcpl_131;
  wire and_dcpl_408;
  wire or_dcpl_137;
  wire mux_tmp_1500;
  wire and_dcpl_416;
  wire and_dcpl_417;
  wire and_dcpl_419;
  wire and_dcpl_421;
  wire and_dcpl_422;
  wire and_dcpl_431;
  wire and_dcpl_432;
  wire and_dcpl_434;
  wire and_dcpl_436;
  wire and_dcpl_437;
  wire and_dcpl_446;
  wire and_dcpl_447;
  wire and_dcpl_449;
  wire and_dcpl_451;
  wire and_dcpl_452;
  wire and_dcpl_473;
  wire and_dcpl_474;
  wire and_dcpl_476;
  wire and_dcpl_478;
  wire and_dcpl_479;
  wire and_dcpl_504;
  wire and_dcpl_505;
  wire and_dcpl_507;
  wire and_dcpl_509;
  wire and_dcpl_510;
  wire and_dcpl_519;
  wire and_dcpl_520;
  wire and_dcpl_522;
  wire and_dcpl_524;
  wire and_dcpl_525;
  wire and_dcpl_534;
  wire and_dcpl_535;
  wire and_dcpl_537;
  wire and_dcpl_539;
  wire and_dcpl_540;
  wire and_dcpl_549;
  wire and_dcpl_550;
  wire and_dcpl_552;
  wire and_dcpl_554;
  wire and_dcpl_555;
  wire or_dcpl_219;
  wire and_dcpl_564;
  wire and_dcpl_565;
  wire and_dcpl_567;
  wire and_dcpl_569;
  wire and_dcpl_570;
  wire and_dcpl_575;
  wire and_dcpl_576;
  wire and_dcpl_578;
  wire and_dcpl_580;
  wire and_dcpl_581;
  wire and_dcpl_586;
  wire and_dcpl_587;
  wire and_dcpl_589;
  wire and_dcpl_591;
  wire and_dcpl_592;
  wire and_dcpl_597;
  wire and_dcpl_598;
  wire and_dcpl_600;
  wire and_dcpl_602;
  wire and_dcpl_603;
  wire and_dcpl_608;
  wire and_dcpl_609;
  wire and_dcpl_611;
  wire and_dcpl_613;
  wire and_dcpl_614;
  wire and_dcpl_619;
  wire and_dcpl_620;
  wire and_dcpl_622;
  wire and_dcpl_624;
  wire and_dcpl_625;
  wire and_dcpl_630;
  wire and_dcpl_631;
  wire and_dcpl_633;
  wire and_dcpl_635;
  wire and_dcpl_636;
  wire and_dcpl_638;
  wire or_dcpl_295;
  wire and_dcpl_676;
  wire and_dcpl_695;
  wire and_dcpl_698;
  wire and_dcpl_701;
  wire and_dcpl_704;
  wire and_dcpl_707;
  wire and_dcpl_711;
  wire and_dcpl_714;
  wire and_dcpl_722;
  wire and_dcpl_725;
  wire and_dcpl_733;
  wire and_dcpl_736;
  wire and_dcpl_744;
  wire and_dcpl_747;
  wire and_dcpl_755;
  wire and_dcpl_758;
  wire and_dcpl_766;
  wire and_dcpl_769;
  wire and_dcpl_777;
  wire and_dcpl_780;
  wire and_dcpl_788;
  wire and_dcpl_791;
  wire and_dcpl_799;
  wire and_dcpl_802;
  wire and_dcpl_810;
  wire and_dcpl_813;
  wire and_dcpl_821;
  wire and_dcpl_824;
  wire and_dcpl_830;
  wire nor_tmp_847;
  wire and_dcpl_832;
  wire and_dcpl_834;
  wire and_dcpl_840;
  wire and_dcpl_843;
  wire and_dcpl_844;
  wire and_dcpl_846;
  wire and_dcpl_848;
  wire and_dcpl_856;
  wire and_dcpl_858;
  wire and_dcpl_879;
  wire and_dcpl_884;
  wire and_dcpl_886;
  wire and_dcpl_897;
  wire and_dcpl_899;
  wire and_dcpl_924;
  wire and_dcpl_926;
  wire and_dcpl_946;
  wire and_dcpl_948;
  wire and_dcpl_971;
  wire and_dcpl_1036;
  wire and_dcpl_1038;
  wire mux_tmp_1541;
  wire and_dcpl_1044;
  wire and_dcpl_1046;
  wire and_dcpl_1048;
  wire and_dcpl_1050;
  wire mux_tmp_1542;
  wire and_dcpl_1052;
  wire and_dcpl_1054;
  wire mux_tmp_1543;
  wire and_dcpl_1060;
  wire and_dcpl_1062;
  wire and_dcpl_1070;
  wire and_dcpl_1073;
  wire or_dcpl_391;
  wire or_dcpl_393;
  wire and_dcpl_1079;
  wire and_dcpl_1080;
  wire or_dcpl_394;
  wire and_dcpl_1084;
  wire and_dcpl_1087;
  wire or_dcpl_411;
  wire and_dcpl_1093;
  wire and_dcpl_1094;
  wire or_dcpl_413;
  wire or_dcpl_414;
  wire and_dcpl_1098;
  wire and_dcpl_1101;
  wire or_dcpl_429;
  wire and_dcpl_1107;
  wire and_dcpl_1108;
  wire and_dcpl_1112;
  wire and_dcpl_1115;
  wire or_dcpl_447;
  wire and_dcpl_1121;
  wire and_dcpl_1122;
  wire and_dcpl_1123;
  wire and_dcpl_1126;
  wire and_dcpl_1129;
  wire or_dcpl_465;
  wire and_dcpl_1134;
  wire and_dcpl_1135;
  wire or_dcpl_477;
  wire or_dcpl_483;
  wire and_dcpl_1152;
  wire and_dcpl_1153;
  wire or_dcpl_495;
  wire or_dcpl_501;
  wire and_dcpl_1170;
  wire and_dcpl_1171;
  wire or_dcpl_513;
  wire or_dcpl_519;
  wire and_dcpl_1188;
  wire and_dcpl_1189;
  wire or_dcpl_520;
  wire or_dcpl_531;
  wire or_dcpl_537;
  wire and_dcpl_1206;
  wire and_dcpl_1207;
  wire and_dcpl_1211;
  wire and_dcpl_1214;
  wire or_dcpl_555;
  wire and_dcpl_1220;
  wire and_dcpl_1221;
  wire or_dcpl_567;
  wire or_dcpl_573;
  wire and_dcpl_1238;
  wire and_dcpl_1239;
  wire or_dcpl_585;
  wire or_dcpl_591;
  wire and_dcpl_1256;
  wire and_dcpl_1257;
  wire or_dcpl_603;
  wire or_dcpl_609;
  wire and_dcpl_1274;
  wire and_dcpl_1275;
  wire and_dcpl_1279;
  wire and_dcpl_1283;
  wire or_dcpl_627;
  wire and_dcpl_1289;
  wire and_dcpl_1290;
  wire or_dcpl_639;
  wire or_dcpl_645;
  wire and_dcpl_1307;
  wire and_dcpl_1308;
  wire or_dcpl_657;
  wire or_dcpl_663;
  wire and_dcpl_1325;
  wire and_dcpl_1326;
  wire or_dcpl_675;
  wire and_dcpl_1329;
  wire and_dcpl_1333;
  wire and_dcpl_1335;
  wire and_dcpl_1341;
  wire and_dcpl_1347;
  wire and_dcpl_1353;
  wire and_dcpl_1359;
  wire and_dcpl_1365;
  wire and_dcpl_1371;
  wire and_dcpl_1377;
  wire and_dcpl_1383;
  wire and_dcpl_1389;
  wire and_dcpl_1395;
  wire and_dcpl_1401;
  wire and_dcpl_1407;
  wire and_dcpl_1413;
  wire and_dcpl_1419;
  wire and_dcpl_1425;
  wire or_dcpl_677;
  wire or_dcpl_678;
  wire and_dcpl_1426;
  wire or_dcpl_679;
  wire or_dcpl_681;
  wire or_dcpl_683;
  wire or_dcpl_686;
  wire or_dcpl_688;
  wire or_dcpl_692;
  wire or_dcpl_694;
  wire or_dcpl_696;
  wire or_dcpl_699;
  wire and_dcpl_1468;
  wire and_dcpl_1471;
  wire and_dcpl_1472;
  wire and_dcpl_1476;
  wire and_dcpl_1477;
  wire and_dcpl_1483;
  wire and_dcpl_1490;
  wire and_dcpl_1497;
  wire and_dcpl_1504;
  wire and_dcpl_1511;
  wire and_dcpl_1518;
  wire and_dcpl_1525;
  wire and_dcpl_1532;
  wire and_dcpl_1539;
  wire and_dcpl_1546;
  wire and_dcpl_1553;
  wire and_dcpl_1560;
  wire and_dcpl_1567;
  wire and_dcpl_1574;
  wire and_dcpl_1581;
  wire and_dcpl_1588;
  wire and_dcpl_1595;
  wire and_dcpl_1602;
  wire and_dcpl_1609;
  wire and_dcpl_1616;
  wire and_dcpl_1623;
  wire and_dcpl_1630;
  wire and_dcpl_1637;
  wire and_dcpl_1644;
  wire and_dcpl_1651;
  wire and_dcpl_1658;
  wire and_dcpl_1665;
  wire and_dcpl_1672;
  wire and_dcpl_1679;
  wire and_dcpl_1682;
  wire and_dcpl_1686;
  wire and_dcpl_1691;
  wire and_dcpl_1692;
  wire or_dcpl_775;
  wire or_dcpl_777;
  wire or_dcpl_780;
  wire or_dcpl_783;
  wire or_dcpl_785;
  wire or_dcpl_787;
  wire or_dcpl_790;
  wire or_dcpl_823;
  wire or_dcpl_830;
  wire or_dcpl_837;
  wire or_dcpl_844;
  wire or_dcpl_851;
  wire or_dcpl_859;
  wire or_dcpl_872;
  wire or_dcpl_879;
  wire or_dcpl_893;
  wire or_dcpl_901;
  wire or_tmp_3044;
  wire or_tmp_3045;
  wire or_tmp_3048;
  wire or_tmp_3190;
  wire or_tmp_3201;
  wire or_tmp_3212;
  wire or_tmp_3223;
  wire or_tmp_3234;
  wire or_tmp_3245;
  wire or_tmp_3256;
  wire or_tmp_3267;
  wire or_tmp_3278;
  wire or_tmp_3289;
  wire or_tmp_3300;
  wire or_tmp_3311;
  wire or_tmp_3322;
  wire or_tmp_3333;
  wire or_tmp_3344;
  wire or_tmp_3355;
  wire or_tmp_3479;
  reg alu_nan_to_zero_op_sign_1_lpi_1_dfm;
  reg alu_nan_to_zero_op_sign_2_lpi_1_dfm;
  reg alu_nan_to_zero_op_sign_3_lpi_1_dfm;
  reg alu_nan_to_zero_op_sign_4_lpi_1_dfm;
  reg alu_nan_to_zero_op_sign_5_lpi_1_dfm;
  reg alu_nan_to_zero_op_sign_6_lpi_1_dfm;
  reg alu_nan_to_zero_op_sign_7_lpi_1_dfm;
  reg alu_nan_to_zero_op_sign_8_lpi_1_dfm;
  reg alu_nan_to_zero_op_sign_9_lpi_1_dfm;
  reg alu_nan_to_zero_op_sign_10_lpi_1_dfm;
  reg alu_nan_to_zero_op_sign_11_lpi_1_dfm;
  reg alu_nan_to_zero_op_sign_12_lpi_1_dfm;
  reg alu_nan_to_zero_op_sign_13_lpi_1_dfm;
  reg alu_nan_to_zero_op_sign_14_lpi_1_dfm;
  reg alu_nan_to_zero_op_sign_15_lpi_1_dfm;
  reg alu_nan_to_zero_op_sign_lpi_1_dfm;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3;
  reg alu_loop_op_1_FpAdd_8U_23U_is_a_greater_slc_8_svs;
  reg alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_svs;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_1_sva;
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm;
  reg FpAlu_8U_23U_equal_tmp;
  reg alu_loop_op_1_FpCmp_8U_23U_true_else_slc_8_svs;
  reg FpAlu_8U_23U_equal_tmp_1;
  reg FpAlu_8U_23U_equal_tmp_2;
  reg alu_loop_op_1_FpCmp_8U_23U_false_else_slc_8_svs;
  reg FpAlu_8U_23U_nor_dfs;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3;
  reg alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_2_sva;
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm;
  reg alu_loop_op_2_FpCmp_8U_23U_true_else_slc_8_1_svs;
  reg alu_loop_op_2_FpCmp_8U_23U_false_else_slc_8_1_svs;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3;
  reg alu_loop_op_3_FpAdd_8U_23U_is_a_greater_slc_8_svs;
  reg alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_svs;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_3_sva;
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm;
  reg alu_loop_op_3_FpCmp_8U_23U_true_else_slc_8_svs;
  reg alu_loop_op_3_FpCmp_8U_23U_false_else_slc_8_svs;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3;
  reg alu_loop_op_4_FpAdd_8U_23U_is_a_greater_slc_8_1_svs;
  reg alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_4_sva;
  reg IsNaN_8U_23U_1_land_4_lpi_1_dfm;
  reg alu_loop_op_4_FpCmp_8U_23U_true_else_slc_8_1_svs;
  reg alu_loop_op_4_FpCmp_8U_23U_false_else_slc_8_1_svs;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3;
  reg alu_loop_op_5_FpAdd_8U_23U_is_a_greater_slc_8_svs;
  reg alu_loop_op_5_FpAdd_8U_23U_is_a_greater_oif_equal_svs;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_5_sva;
  reg IsNaN_8U_23U_1_land_5_lpi_1_dfm;
  reg alu_loop_op_5_FpCmp_8U_23U_true_else_slc_8_svs;
  reg alu_loop_op_5_FpCmp_8U_23U_false_else_slc_8_svs;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3;
  reg alu_loop_op_6_FpAdd_8U_23U_is_a_greater_slc_8_1_svs;
  reg alu_loop_op_6_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_6_sva;
  reg IsNaN_8U_23U_1_land_6_lpi_1_dfm;
  reg alu_loop_op_6_FpCmp_8U_23U_true_else_slc_8_1_svs;
  reg alu_loop_op_6_FpCmp_8U_23U_false_else_slc_8_1_svs;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3;
  reg alu_loop_op_7_FpAdd_8U_23U_is_a_greater_slc_8_svs;
  reg alu_loop_op_7_FpAdd_8U_23U_is_a_greater_oif_equal_svs;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_7_sva;
  reg IsNaN_8U_23U_1_land_7_lpi_1_dfm;
  reg alu_loop_op_7_FpCmp_8U_23U_true_else_slc_8_svs;
  reg alu_loop_op_7_FpCmp_8U_23U_false_else_slc_8_svs;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3;
  reg alu_loop_op_8_FpAdd_8U_23U_is_a_greater_slc_8_1_svs;
  reg alu_loop_op_8_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_8_sva;
  reg IsNaN_8U_23U_1_land_8_lpi_1_dfm;
  reg alu_loop_op_8_FpCmp_8U_23U_true_else_slc_8_1_svs;
  reg alu_loop_op_8_FpCmp_8U_23U_false_else_slc_8_1_svs;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3;
  reg alu_loop_op_9_FpAdd_8U_23U_is_a_greater_slc_8_svs;
  reg alu_loop_op_9_FpAdd_8U_23U_is_a_greater_oif_equal_svs;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_9_sva;
  reg IsNaN_8U_23U_1_land_9_lpi_1_dfm;
  reg alu_loop_op_9_FpCmp_8U_23U_true_else_slc_8_svs;
  reg alu_loop_op_9_FpCmp_8U_23U_false_else_slc_8_svs;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3;
  reg alu_loop_op_10_FpAdd_8U_23U_is_a_greater_slc_8_1_svs;
  reg alu_loop_op_10_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_10_sva;
  reg IsNaN_8U_23U_1_land_10_lpi_1_dfm;
  reg alu_loop_op_10_FpCmp_8U_23U_true_else_slc_8_1_svs;
  reg alu_loop_op_10_FpCmp_8U_23U_false_else_slc_8_1_svs;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3;
  reg alu_loop_op_11_FpAdd_8U_23U_is_a_greater_slc_8_svs;
  reg alu_loop_op_11_FpAdd_8U_23U_is_a_greater_oif_equal_svs;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_11_sva;
  reg IsNaN_8U_23U_1_land_11_lpi_1_dfm;
  reg alu_loop_op_11_FpCmp_8U_23U_true_else_slc_8_svs;
  reg alu_loop_op_11_FpCmp_8U_23U_false_else_slc_8_svs;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3;
  reg alu_loop_op_12_FpAdd_8U_23U_is_a_greater_slc_8_1_svs;
  reg alu_loop_op_12_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_12_sva;
  reg IsNaN_8U_23U_1_land_12_lpi_1_dfm;
  reg alu_loop_op_12_FpCmp_8U_23U_true_else_slc_8_1_svs;
  reg alu_loop_op_12_FpCmp_8U_23U_false_else_slc_8_1_svs;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3;
  reg alu_loop_op_13_FpAdd_8U_23U_is_a_greater_slc_8_svs;
  reg alu_loop_op_13_FpAdd_8U_23U_is_a_greater_oif_equal_svs;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_13_sva;
  reg IsNaN_8U_23U_1_land_13_lpi_1_dfm;
  reg alu_loop_op_13_FpCmp_8U_23U_true_else_slc_8_svs;
  reg alu_loop_op_13_FpCmp_8U_23U_false_else_slc_8_svs;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3;
  reg alu_loop_op_14_FpAdd_8U_23U_is_a_greater_slc_8_1_svs;
  reg alu_loop_op_14_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_14_sva;
  reg IsNaN_8U_23U_1_land_14_lpi_1_dfm;
  reg alu_loop_op_14_FpCmp_8U_23U_true_else_slc_8_1_svs;
  reg alu_loop_op_14_FpCmp_8U_23U_false_else_slc_8_1_svs;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3;
  reg alu_loop_op_15_FpAdd_8U_23U_is_a_greater_slc_8_svs;
  reg alu_loop_op_15_FpAdd_8U_23U_is_a_greater_oif_equal_svs;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_15_sva;
  reg IsNaN_8U_23U_1_land_15_lpi_1_dfm;
  reg alu_loop_op_15_FpCmp_8U_23U_true_else_slc_8_svs;
  reg alu_loop_op_15_FpCmp_8U_23U_false_else_slc_8_svs;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3;
  reg alu_loop_op_16_FpAdd_8U_23U_is_a_greater_slc_8_1_svs;
  reg alu_loop_op_16_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_lpi_1_dfm;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_sva;
  reg IsNaN_8U_23U_1_land_lpi_1_dfm;
  reg alu_loop_op_16_FpCmp_8U_23U_true_else_slc_8_1_svs;
  reg alu_loop_op_16_FpCmp_8U_23U_false_else_slc_8_1_svs;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_1_sva;
  reg IntShiftLeft_16U_6U_32U_return_0_1_sva;
  reg IntShiftLeft_16U_6U_32U_return_31_1_sva;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_2_sva;
  reg IntShiftLeft_16U_6U_32U_return_0_2_sva;
  reg IntShiftLeft_16U_6U_32U_return_31_2_sva;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_3_sva;
  reg IntShiftLeft_16U_6U_32U_return_0_3_sva;
  reg IntShiftLeft_16U_6U_32U_return_31_3_sva;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_4_sva;
  reg IntShiftLeft_16U_6U_32U_return_0_4_sva;
  reg IntShiftLeft_16U_6U_32U_return_31_4_sva;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_5_sva;
  reg IntShiftLeft_16U_6U_32U_return_0_5_sva;
  reg IntShiftLeft_16U_6U_32U_return_31_5_sva;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_6_sva;
  reg IntShiftLeft_16U_6U_32U_return_0_6_sva;
  reg IntShiftLeft_16U_6U_32U_return_31_6_sva;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_7_sva;
  reg IntShiftLeft_16U_6U_32U_return_0_7_sva;
  reg IntShiftLeft_16U_6U_32U_return_31_7_sva;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_8_sva;
  reg IntShiftLeft_16U_6U_32U_return_0_8_sva;
  reg IntShiftLeft_16U_6U_32U_return_31_8_sva;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_9_sva;
  reg IntShiftLeft_16U_6U_32U_return_0_9_sva;
  reg IntShiftLeft_16U_6U_32U_return_31_9_sva;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_10_sva;
  reg IntShiftLeft_16U_6U_32U_return_0_10_sva;
  reg IntShiftLeft_16U_6U_32U_return_31_10_sva;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_11_sva;
  reg IntShiftLeft_16U_6U_32U_return_0_11_sva;
  reg IntShiftLeft_16U_6U_32U_return_31_11_sva;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_12_sva;
  reg IntShiftLeft_16U_6U_32U_return_0_12_sva;
  reg IntShiftLeft_16U_6U_32U_return_31_12_sva;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_13_sva;
  reg IntShiftLeft_16U_6U_32U_return_0_13_sva;
  reg IntShiftLeft_16U_6U_32U_return_31_13_sva;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_14_sva;
  reg IntShiftLeft_16U_6U_32U_return_0_14_sva;
  reg IntShiftLeft_16U_6U_32U_return_31_14_sva;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_15_sva;
  reg IntShiftLeft_16U_6U_32U_return_0_15_sva;
  reg IntShiftLeft_16U_6U_32U_return_31_15_sva;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_sva;
  reg IntShiftLeft_16U_6U_32U_return_0_sva;
  reg IntShiftLeft_16U_6U_32U_return_31_sva;
  reg main_stage_v_1;
  reg main_stage_v_2;
  reg main_stage_v_3;
  reg main_stage_v_4;
  reg FpCmp_8U_23U_false_is_a_greater_lpi_1_dfm_7;
  reg IsNaN_8U_23U_3_land_lpi_1_dfm_6;
  reg IsNaN_8U_23U_3_land_lpi_1_dfm_7;
  reg FpCmp_8U_23U_false_is_a_greater_15_lpi_1_dfm_7;
  reg IsNaN_8U_23U_3_land_15_lpi_1_dfm_6;
  reg IsNaN_8U_23U_3_land_15_lpi_1_dfm_7;
  reg FpCmp_8U_23U_false_is_a_greater_14_lpi_1_dfm_7;
  reg IsNaN_8U_23U_3_land_14_lpi_1_dfm_6;
  reg IsNaN_8U_23U_3_land_14_lpi_1_dfm_7;
  reg FpCmp_8U_23U_false_is_a_greater_13_lpi_1_dfm_7;
  reg IsNaN_8U_23U_3_land_13_lpi_1_dfm_6;
  reg IsNaN_8U_23U_3_land_13_lpi_1_dfm_7;
  reg FpCmp_8U_23U_false_is_a_greater_12_lpi_1_dfm_7;
  reg IsNaN_8U_23U_3_land_12_lpi_1_dfm_6;
  reg IsNaN_8U_23U_3_land_12_lpi_1_dfm_7;
  reg FpCmp_8U_23U_false_is_a_greater_11_lpi_1_dfm_7;
  reg IsNaN_8U_23U_3_land_11_lpi_1_dfm_6;
  reg IsNaN_8U_23U_3_land_11_lpi_1_dfm_7;
  reg FpCmp_8U_23U_false_is_a_greater_10_lpi_1_dfm_7;
  reg IsNaN_8U_23U_3_land_10_lpi_1_dfm_6;
  reg IsNaN_8U_23U_3_land_10_lpi_1_dfm_7;
  reg FpCmp_8U_23U_false_is_a_greater_9_lpi_1_dfm_7;
  reg IsNaN_8U_23U_3_land_9_lpi_1_dfm_6;
  reg IsNaN_8U_23U_3_land_9_lpi_1_dfm_7;
  reg FpCmp_8U_23U_false_is_a_greater_8_lpi_1_dfm_7;
  reg IsNaN_8U_23U_3_land_8_lpi_1_dfm_6;
  reg IsNaN_8U_23U_3_land_8_lpi_1_dfm_7;
  reg FpCmp_8U_23U_false_is_a_greater_7_lpi_1_dfm_7;
  reg IsNaN_8U_23U_3_land_7_lpi_1_dfm_6;
  reg IsNaN_8U_23U_3_land_7_lpi_1_dfm_7;
  reg FpCmp_8U_23U_false_is_a_greater_6_lpi_1_dfm_7;
  reg IsNaN_8U_23U_3_land_6_lpi_1_dfm_6;
  reg IsNaN_8U_23U_3_land_6_lpi_1_dfm_7;
  reg FpCmp_8U_23U_false_is_a_greater_5_lpi_1_dfm_7;
  reg IsNaN_8U_23U_3_land_5_lpi_1_dfm_6;
  reg IsNaN_8U_23U_3_land_5_lpi_1_dfm_7;
  reg FpCmp_8U_23U_false_is_a_greater_4_lpi_1_dfm_7;
  reg IsNaN_8U_23U_3_land_4_lpi_1_dfm_6;
  reg IsNaN_8U_23U_3_land_4_lpi_1_dfm_7;
  reg FpCmp_8U_23U_false_is_a_greater_3_lpi_1_dfm_7;
  reg IsNaN_8U_23U_3_land_3_lpi_1_dfm_6;
  reg IsNaN_8U_23U_3_land_3_lpi_1_dfm_7;
  reg FpCmp_8U_23U_false_is_a_greater_2_lpi_1_dfm_7;
  reg IsNaN_8U_23U_3_land_2_lpi_1_dfm_6;
  reg IsNaN_8U_23U_3_land_2_lpi_1_dfm_7;
  reg FpCmp_8U_23U_false_is_a_greater_1_lpi_1_dfm_7;
  reg IsNaN_8U_23U_3_land_1_lpi_1_dfm_6;
  reg IsNaN_8U_23U_3_land_1_lpi_1_dfm_7;
  reg IsNaN_8U_23U_4_land_lpi_1_dfm_4;
  reg IsNaN_8U_23U_4_land_lpi_1_dfm_6;
  reg IsNaN_8U_23U_land_lpi_1_dfm_4;
  reg IsNaN_8U_23U_land_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_lpi_1_dfm_10;
  reg IsNaN_8U_23U_4_land_15_lpi_1_dfm_4;
  reg IsNaN_8U_23U_4_land_15_lpi_1_dfm_6;
  reg IsNaN_8U_23U_land_15_lpi_1_dfm_4;
  reg IsNaN_8U_23U_land_15_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_15_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_15_lpi_1_dfm_10;
  reg IsNaN_8U_23U_4_land_14_lpi_1_dfm_4;
  reg IsNaN_8U_23U_4_land_14_lpi_1_dfm_6;
  reg IsNaN_8U_23U_2_land_14_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_14_lpi_1_dfm_4;
  reg IsNaN_8U_23U_land_14_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_14_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_14_lpi_1_dfm_10;
  reg IsNaN_8U_23U_4_land_13_lpi_1_dfm_4;
  reg IsNaN_8U_23U_4_land_13_lpi_1_dfm_6;
  reg IsNaN_8U_23U_2_land_13_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_13_lpi_1_dfm_4;
  reg IsNaN_8U_23U_land_13_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_13_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_13_lpi_1_dfm_10;
  reg IsNaN_8U_23U_4_land_12_lpi_1_dfm_4;
  reg IsNaN_8U_23U_4_land_12_lpi_1_dfm_6;
  reg IsNaN_8U_23U_2_land_12_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_12_lpi_1_dfm_4;
  reg IsNaN_8U_23U_land_12_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_12_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_12_lpi_1_dfm_10;
  reg IsNaN_8U_23U_4_land_11_lpi_1_dfm_4;
  reg IsNaN_8U_23U_4_land_11_lpi_1_dfm_6;
  reg IsNaN_8U_23U_2_land_11_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_11_lpi_1_dfm_4;
  reg IsNaN_8U_23U_land_11_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_11_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_11_lpi_1_dfm_10;
  reg IsNaN_8U_23U_4_land_10_lpi_1_dfm_4;
  reg IsNaN_8U_23U_4_land_10_lpi_1_dfm_6;
  reg IsNaN_8U_23U_2_land_10_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_10_lpi_1_dfm_4;
  reg IsNaN_8U_23U_land_10_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_10_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_10_lpi_1_dfm_10;
  reg IsNaN_8U_23U_4_land_9_lpi_1_dfm_4;
  reg IsNaN_8U_23U_4_land_9_lpi_1_dfm_6;
  reg IsNaN_8U_23U_2_land_9_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_9_lpi_1_dfm_4;
  reg IsNaN_8U_23U_land_9_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_9_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_9_lpi_1_dfm_10;
  reg IsNaN_8U_23U_4_land_8_lpi_1_dfm_4;
  reg IsNaN_8U_23U_4_land_8_lpi_1_dfm_6;
  reg IsNaN_8U_23U_land_8_lpi_1_dfm_4;
  reg IsNaN_8U_23U_land_8_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_8_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_8_lpi_1_dfm_10;
  reg IsNaN_8U_23U_4_land_7_lpi_1_dfm_4;
  reg IsNaN_8U_23U_4_land_7_lpi_1_dfm_6;
  reg IsNaN_8U_23U_land_7_lpi_1_dfm_4;
  reg IsNaN_8U_23U_land_7_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_7_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_7_lpi_1_dfm_10;
  reg IsNaN_8U_23U_4_land_6_lpi_1_dfm_4;
  reg IsNaN_8U_23U_4_land_6_lpi_1_dfm_6;
  reg IsNaN_8U_23U_2_land_6_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_6_lpi_1_dfm_4;
  reg IsNaN_8U_23U_land_6_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_6_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_6_lpi_1_dfm_10;
  reg IsNaN_8U_23U_4_land_5_lpi_1_dfm_4;
  reg IsNaN_8U_23U_4_land_5_lpi_1_dfm_6;
  reg IsNaN_8U_23U_2_land_5_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_5_lpi_1_dfm_4;
  reg IsNaN_8U_23U_land_5_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_5_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_5_lpi_1_dfm_10;
  reg IsNaN_8U_23U_4_land_4_lpi_1_dfm_4;
  reg IsNaN_8U_23U_4_land_4_lpi_1_dfm_6;
  reg IsNaN_8U_23U_2_land_4_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_4_lpi_1_dfm_4;
  reg IsNaN_8U_23U_land_4_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_4_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_4_lpi_1_dfm_10;
  reg IsNaN_8U_23U_4_land_3_lpi_1_dfm_4;
  reg IsNaN_8U_23U_4_land_3_lpi_1_dfm_6;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_4;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_10;
  reg IsNaN_8U_23U_4_land_2_lpi_1_dfm_4;
  reg IsNaN_8U_23U_4_land_2_lpi_1_dfm_6;
  reg IsNaN_8U_23U_2_land_2_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_4;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_10;
  reg IsNaN_8U_23U_4_land_1_lpi_1_dfm_4;
  reg IsNaN_8U_23U_4_land_1_lpi_1_dfm_6;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_4;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_10;
  reg alu_loop_op_else_nor_tmp_16;
  reg alu_loop_op_else_nor_tmp_80;
  reg alu_loop_op_else_nor_tmp_81;
  reg alu_loop_op_else_nor_tmp_82;
  reg [32:0] AluOut_data_15_sva_7;
  wire [33:0] nl_AluOut_data_15_sva_7;
  reg [32:0] AluOut_data_15_sva_8;
  reg [32:0] AluOut_data_14_sva_7;
  wire [33:0] nl_AluOut_data_14_sva_7;
  reg [32:0] AluOut_data_14_sva_8;
  reg [32:0] AluOut_data_13_sva_7;
  wire [33:0] nl_AluOut_data_13_sva_7;
  reg [32:0] AluOut_data_13_sva_8;
  reg [32:0] AluOut_data_12_sva_7;
  wire [33:0] nl_AluOut_data_12_sva_7;
  reg [32:0] AluOut_data_12_sva_8;
  reg [32:0] AluOut_data_11_sva_7;
  wire [33:0] nl_AluOut_data_11_sva_7;
  reg [32:0] AluOut_data_11_sva_8;
  reg [32:0] AluOut_data_10_sva_7;
  wire [33:0] nl_AluOut_data_10_sva_7;
  reg [32:0] AluOut_data_10_sva_8;
  reg [32:0] AluOut_data_9_sva_7;
  wire [33:0] nl_AluOut_data_9_sva_7;
  reg [32:0] AluOut_data_9_sva_8;
  reg [32:0] AluOut_data_8_sva_7;
  wire [33:0] nl_AluOut_data_8_sva_7;
  reg [32:0] AluOut_data_8_sva_8;
  reg [32:0] AluOut_data_7_sva_7;
  wire [33:0] nl_AluOut_data_7_sva_7;
  reg [32:0] AluOut_data_7_sva_8;
  reg [32:0] AluOut_data_6_sva_7;
  wire [33:0] nl_AluOut_data_6_sva_7;
  reg [32:0] AluOut_data_6_sva_8;
  reg [32:0] AluOut_data_5_sva_7;
  wire [33:0] nl_AluOut_data_5_sva_7;
  reg [32:0] AluOut_data_5_sva_8;
  reg [32:0] AluOut_data_4_sva_7;
  wire [33:0] nl_AluOut_data_4_sva_7;
  reg [32:0] AluOut_data_4_sva_8;
  reg [32:0] AluOut_data_3_sva_7;
  wire [33:0] nl_AluOut_data_3_sva_7;
  reg [32:0] AluOut_data_3_sva_8;
  reg [32:0] AluOut_data_2_sva_7;
  wire [33:0] nl_AluOut_data_2_sva_7;
  reg [32:0] AluOut_data_2_sva_8;
  reg [32:0] AluOut_data_1_sva_7;
  wire [33:0] nl_AluOut_data_1_sva_7;
  reg [32:0] AluOut_data_1_sva_8;
  reg [32:0] AluOut_data_0_sva_7;
  wire [33:0] nl_AluOut_data_0_sva_7;
  reg [32:0] AluOut_data_0_sva_8;
  reg [22:0] FpCmp_8U_23U_false_o_22_0_lpi_1_dfm_6;
  reg FpAlu_8U_23U_o_0_sva_6;
  reg FpAlu_8U_23U_o_0_sva_7;
  reg [22:0] FpCmp_8U_23U_true_o_22_0_lpi_1_dfm_6;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_2;
  reg [22:0] FpCmp_8U_23U_false_o_22_0_15_lpi_1_dfm_6;
  reg FpAlu_8U_23U_o_0_15_sva_6;
  reg FpAlu_8U_23U_o_0_15_sva_7;
  reg [22:0] FpCmp_8U_23U_true_o_22_0_15_lpi_1_dfm_6;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_15_sva_2;
  reg [22:0] FpCmp_8U_23U_false_o_22_0_14_lpi_1_dfm_6;
  reg FpAlu_8U_23U_o_0_14_sva_6;
  reg FpAlu_8U_23U_o_0_14_sva_7;
  reg [22:0] FpCmp_8U_23U_true_o_22_0_14_lpi_1_dfm_6;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_14_sva_2;
  reg [22:0] FpCmp_8U_23U_false_o_22_0_13_lpi_1_dfm_6;
  reg FpAlu_8U_23U_o_0_13_sva_6;
  reg FpAlu_8U_23U_o_0_13_sva_7;
  reg [22:0] FpCmp_8U_23U_true_o_22_0_13_lpi_1_dfm_6;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_13_sva_2;
  reg [22:0] FpCmp_8U_23U_false_o_22_0_12_lpi_1_dfm_6;
  reg FpAlu_8U_23U_o_0_12_sva_6;
  reg FpAlu_8U_23U_o_0_12_sva_7;
  reg [22:0] FpCmp_8U_23U_true_o_22_0_12_lpi_1_dfm_6;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_12_sva_2;
  reg [22:0] FpCmp_8U_23U_false_o_22_0_11_lpi_1_dfm_6;
  reg FpAlu_8U_23U_o_0_11_sva_6;
  reg FpAlu_8U_23U_o_0_11_sva_7;
  reg [22:0] FpCmp_8U_23U_true_o_22_0_11_lpi_1_dfm_6;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_11_sva_2;
  reg [22:0] FpCmp_8U_23U_false_o_22_0_10_lpi_1_dfm_6;
  reg FpAlu_8U_23U_o_0_10_sva_6;
  reg FpAlu_8U_23U_o_0_10_sva_7;
  reg [22:0] FpCmp_8U_23U_true_o_22_0_10_lpi_1_dfm_6;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_10_sva_2;
  reg [22:0] FpCmp_8U_23U_false_o_22_0_9_lpi_1_dfm_6;
  reg FpAlu_8U_23U_o_0_9_sva_6;
  reg FpAlu_8U_23U_o_0_9_sva_7;
  reg [22:0] FpCmp_8U_23U_true_o_22_0_9_lpi_1_dfm_6;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_9_sva_2;
  reg [22:0] FpCmp_8U_23U_false_o_22_0_8_lpi_1_dfm_6;
  reg FpAlu_8U_23U_o_0_8_sva_6;
  reg FpAlu_8U_23U_o_0_8_sva_7;
  reg [22:0] FpCmp_8U_23U_true_o_22_0_8_lpi_1_dfm_6;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_8_sva_2;
  reg [22:0] FpCmp_8U_23U_false_o_22_0_7_lpi_1_dfm_6;
  reg FpAlu_8U_23U_o_0_7_sva_6;
  reg FpAlu_8U_23U_o_0_7_sva_7;
  reg [22:0] FpCmp_8U_23U_true_o_22_0_7_lpi_1_dfm_6;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_7_sva_2;
  reg [22:0] FpCmp_8U_23U_false_o_22_0_6_lpi_1_dfm_6;
  reg FpAlu_8U_23U_o_0_6_sva_6;
  reg FpAlu_8U_23U_o_0_6_sva_7;
  reg [22:0] FpCmp_8U_23U_true_o_22_0_6_lpi_1_dfm_6;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_6_sva_2;
  reg [22:0] FpCmp_8U_23U_false_o_22_0_5_lpi_1_dfm_6;
  reg FpAlu_8U_23U_o_0_5_sva_6;
  reg FpAlu_8U_23U_o_0_5_sva_7;
  reg [22:0] FpCmp_8U_23U_true_o_22_0_5_lpi_1_dfm_6;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_5_sva_2;
  reg [22:0] FpCmp_8U_23U_false_o_22_0_4_lpi_1_dfm_6;
  reg FpAlu_8U_23U_o_0_4_sva_6;
  reg FpAlu_8U_23U_o_0_4_sva_7;
  reg [22:0] FpCmp_8U_23U_true_o_22_0_4_lpi_1_dfm_6;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_4_sva_2;
  reg [22:0] FpCmp_8U_23U_false_o_22_0_3_lpi_1_dfm_6;
  reg FpAlu_8U_23U_o_0_3_sva_6;
  reg FpAlu_8U_23U_o_0_3_sva_7;
  reg [22:0] FpCmp_8U_23U_true_o_22_0_3_lpi_1_dfm_6;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_2;
  reg [22:0] FpCmp_8U_23U_false_o_22_0_2_lpi_1_dfm_6;
  reg FpAlu_8U_23U_o_0_2_sva_6;
  reg FpAlu_8U_23U_o_0_2_sva_7;
  reg [22:0] FpCmp_8U_23U_true_o_22_0_2_lpi_1_dfm_6;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_2;
  reg [22:0] FpCmp_8U_23U_false_o_22_0_1_lpi_1_dfm_6;
  reg FpAlu_8U_23U_o_0_1_sva_6;
  reg FpAlu_8U_23U_o_0_1_sva_7;
  reg [22:0] FpCmp_8U_23U_true_o_22_0_1_lpi_1_dfm_6;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_2;
  reg [15:0] cfg_alu_op_1_sva_1;
  reg [1:0] cfg_alu_algo_1_sva_1;
  reg [1:0] cfg_alu_algo_1_sva_5;
  reg [1:0] cfg_alu_algo_1_sva_6;
  reg [1:0] cfg_alu_algo_1_sva_7;
  reg [5:0] cfg_alu_shift_value_1_sva_1;
  reg [511:0] AluIn_data_sva_1;
  reg [511:0] AluIn_data_sva_501;
  reg [511:0] AluIn_data_sva_502;
  reg [511:0] AluIn_data_sva_503;
  reg io_read_cfg_alu_bypass_rsc_svs_7;
  reg alu_nan_to_zero_op_sign_1_lpi_1_dfm_4;
  reg alu_nan_to_zero_op_sign_2_lpi_1_dfm_4;
  reg alu_nan_to_zero_op_sign_3_lpi_1_dfm_4;
  reg alu_nan_to_zero_op_sign_4_lpi_1_dfm_4;
  reg alu_nan_to_zero_op_sign_5_lpi_1_dfm_4;
  reg alu_nan_to_zero_op_sign_6_lpi_1_dfm_4;
  reg alu_nan_to_zero_op_sign_7_lpi_1_dfm_4;
  reg alu_nan_to_zero_op_sign_8_lpi_1_dfm_3;
  reg alu_nan_to_zero_op_sign_9_lpi_1_dfm_3;
  reg alu_nan_to_zero_op_sign_10_lpi_1_dfm_3;
  reg alu_nan_to_zero_op_sign_11_lpi_1_dfm_3;
  reg alu_nan_to_zero_op_sign_12_lpi_1_dfm_3;
  reg alu_nan_to_zero_op_sign_13_lpi_1_dfm_3;
  reg alu_nan_to_zero_op_sign_14_lpi_1_dfm_3;
  reg alu_nan_to_zero_op_sign_15_lpi_1_dfm_3;
  reg alu_nan_to_zero_op_sign_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_11;
  reg FpAlu_8U_23U_equal_tmp_144;
  reg FpAlu_8U_23U_equal_tmp_146;
  reg FpAlu_8U_23U_equal_tmp_148;
  reg alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2;
  reg alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_1_sva_2;
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_9;
  reg alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_2;
  reg FpAlu_8U_23U_nor_dfs_48;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_11;
  reg alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2;
  reg alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_2_sva_2;
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_9;
  reg alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_2;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_11;
  reg alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2;
  reg alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_3_sva_2;
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_9;
  reg alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_2;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_11;
  reg alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2;
  reg alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_5;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_4_sva_2;
  reg IsNaN_8U_23U_1_land_4_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_4_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_4_lpi_1_dfm_9;
  reg alu_loop_op_4_FpCmp_8U_23U_false_slc_8_1_svs_2;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_11;
  reg alu_loop_op_5_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2;
  reg alu_loop_op_5_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_5;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_5_sva_2;
  reg IsNaN_8U_23U_1_land_5_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_5_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_5_lpi_1_dfm_9;
  reg alu_loop_op_5_FpCmp_8U_23U_false_slc_8_svs_2;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_11;
  reg alu_loop_op_6_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2;
  reg alu_loop_op_6_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_5;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_6_sva_2;
  reg IsNaN_8U_23U_1_land_6_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_6_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_6_lpi_1_dfm_9;
  reg alu_loop_op_6_FpCmp_8U_23U_false_slc_8_1_svs_2;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_11;
  reg alu_loop_op_7_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2;
  reg alu_loop_op_7_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_5;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_7_sva_2;
  reg IsNaN_8U_23U_1_land_7_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_7_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_7_lpi_1_dfm_9;
  reg alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_2;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_11;
  reg alu_loop_op_8_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2;
  reg alu_loop_op_8_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_5;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_8_sva_2;
  reg IsNaN_8U_23U_1_land_8_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_8_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_8_lpi_1_dfm_9;
  reg alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_2;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_11;
  reg alu_loop_op_9_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2;
  reg alu_loop_op_9_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_5;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_9_sva_2;
  reg IsNaN_8U_23U_1_land_9_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_9_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_9_lpi_1_dfm_9;
  reg alu_loop_op_9_FpCmp_8U_23U_false_slc_8_svs_2;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_11;
  reg alu_loop_op_10_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2;
  reg alu_loop_op_10_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_5;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_10_sva_2;
  reg IsNaN_8U_23U_1_land_10_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_10_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_10_lpi_1_dfm_9;
  reg alu_loop_op_10_FpCmp_8U_23U_false_slc_8_1_svs_2;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_11;
  reg alu_loop_op_11_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2;
  reg alu_loop_op_11_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_5;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_11_sva_2;
  reg IsNaN_8U_23U_1_land_11_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_11_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_11_lpi_1_dfm_9;
  reg alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_2;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_11;
  reg alu_loop_op_12_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2;
  reg alu_loop_op_12_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_5;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_12_sva_2;
  reg IsNaN_8U_23U_1_land_12_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_12_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_12_lpi_1_dfm_9;
  reg alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_2;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_11;
  reg alu_loop_op_13_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2;
  reg alu_loop_op_13_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_5;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_13_sva_2;
  reg IsNaN_8U_23U_1_land_13_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_13_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_13_lpi_1_dfm_9;
  reg alu_loop_op_13_FpCmp_8U_23U_false_slc_8_svs_2;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_11;
  reg alu_loop_op_14_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2;
  reg alu_loop_op_14_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_5;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_14_sva_2;
  reg IsNaN_8U_23U_1_land_14_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_14_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_14_lpi_1_dfm_9;
  reg alu_loop_op_14_FpCmp_8U_23U_false_slc_8_1_svs_2;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_11;
  reg alu_loop_op_15_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2;
  reg alu_loop_op_15_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_5;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_15_sva_2;
  reg IsNaN_8U_23U_1_land_15_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_15_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_15_lpi_1_dfm_9;
  reg alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_2;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_11;
  reg FpAlu_8U_23U_equal_tmp_235;
  reg FpAlu_8U_23U_equal_tmp_237;
  reg FpAlu_8U_23U_equal_tmp_239;
  reg alu_loop_op_16_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2;
  reg alu_loop_op_16_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5;
  reg [5:0] IntLeadZero_49U_leading_sign_49_0_rtn_sva_2;
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_9;
  reg alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_2;
  reg FpAlu_8U_23U_nor_dfs_79;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_1_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_0_1_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_31_1_sva_2;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_2_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_0_2_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_31_2_sva_2;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_3_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_0_3_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_31_3_sva_2;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_4_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_0_4_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_31_4_sva_2;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_5_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_0_5_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_31_5_sva_2;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_6_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_0_6_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_31_6_sva_2;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_7_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_0_7_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_31_7_sva_2;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_8_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_0_8_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_31_8_sva_2;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_9_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_0_9_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_31_9_sva_2;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_10_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_0_10_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_31_10_sva_2;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_11_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_0_11_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_31_11_sva_2;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_12_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_0_12_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_31_12_sva_2;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_13_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_0_13_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_31_13_sva_2;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_14_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_0_14_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_31_14_sva_2;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_15_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_0_15_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_31_15_sva_2;
  reg [29:0] IntShiftLeft_16U_6U_32U_return_30_1_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_0_sva_2;
  reg IntShiftLeft_16U_6U_32U_return_31_sva_2;
  reg cfg_alu_src_1_sva_st;
  reg alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm;
  reg alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
  reg alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  reg alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  reg [7:0] alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_itm;
  reg [7:0] alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_itm_2;
  reg alu_loop_op_1_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm;
  reg alu_loop_op_1_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2;
  reg alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm;
  reg alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3;
  reg alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4;
  reg [7:0] alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_itm;
  reg [7:0] alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_itm_2;
  reg alu_loop_op_1_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm;
  reg alu_loop_op_1_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2;
  reg alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st;
  reg alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_st_2;
  reg FpNormalize_8U_49U_if_or_itm;
  reg FpNormalize_8U_49U_if_or_itm_2;
  reg alu_loop_op_1_FpCmp_8U_23U_true_slc_8_svs_st;
  reg IsNaN_8U_23U_2_land_1_lpi_1_dfm_st;
  reg alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_st;
  reg FpAlu_8U_23U_and_itm;
  reg FpAlu_8U_23U_and_itm_3;
  reg FpAlu_8U_23U_and_itm_4;
  reg FpAlu_8U_23U_or_831_itm_3;
  reg FpAlu_8U_23U_or_831_itm_4;
  reg FpAlu_8U_23U_or_752_itm_3;
  reg FpAlu_8U_23U_or_832_itm;
  reg FpAlu_8U_23U_or_753_itm;
  reg alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_st;
  reg alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm;
  reg alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
  reg alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  reg alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  reg [7:0] alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_1_itm;
  reg [7:0] alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_1_itm_2;
  reg alu_loop_op_2_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm;
  reg alu_loop_op_2_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2;
  reg alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm;
  reg alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2;
  reg [7:0] alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_1_itm;
  reg [7:0] alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_1_itm_2;
  reg alu_loop_op_2_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm;
  reg alu_loop_op_2_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2;
  reg alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st;
  reg alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_st_2;
  reg FpNormalize_8U_49U_if_or_1_itm;
  reg FpNormalize_8U_49U_if_or_1_itm_2;
  reg alu_loop_op_2_FpCmp_8U_23U_true_slc_8_1_svs_st;
  reg IsNaN_8U_23U_2_land_2_lpi_1_dfm_st;
  reg alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_st;
  reg FpAlu_8U_23U_and_4_itm;
  reg FpAlu_8U_23U_and_4_itm_3;
  reg FpAlu_8U_23U_and_4_itm_4;
  reg FpAlu_8U_23U_or_833_itm_3;
  reg FpAlu_8U_23U_or_833_itm_4;
  reg FpAlu_8U_23U_or_755_itm_3;
  reg FpAlu_8U_23U_or_834_itm;
  reg FpAlu_8U_23U_or_756_itm;
  reg alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm;
  reg alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
  reg alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  reg alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  reg [7:0] alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_itm;
  reg [7:0] alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_itm_2;
  reg alu_loop_op_3_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm;
  reg alu_loop_op_3_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2;
  reg alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm;
  reg alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3;
  reg alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4;
  reg [7:0] alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_itm;
  reg [7:0] alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_itm_2;
  reg alu_loop_op_3_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm;
  reg alu_loop_op_3_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2;
  reg alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st;
  reg alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_st_2;
  reg FpNormalize_8U_49U_if_or_2_itm;
  reg FpNormalize_8U_49U_if_or_2_itm_2;
  reg alu_loop_op_3_FpCmp_8U_23U_true_slc_8_svs_st;
  reg IsNaN_8U_23U_2_land_3_lpi_1_dfm_st;
  reg alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_st;
  reg FpAlu_8U_23U_and_8_itm;
  reg FpAlu_8U_23U_and_8_itm_3;
  reg FpAlu_8U_23U_and_8_itm_4;
  reg FpAlu_8U_23U_or_835_itm_3;
  reg FpAlu_8U_23U_or_835_itm_4;
  reg FpAlu_8U_23U_or_758_itm_3;
  reg FpAlu_8U_23U_or_836_itm;
  reg FpAlu_8U_23U_or_759_itm;
  reg alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm;
  reg alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
  reg alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  reg alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  reg [7:0] alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_1_itm;
  reg [7:0] alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_1_itm_2;
  reg alu_loop_op_4_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm;
  reg alu_loop_op_4_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2;
  reg alu_loop_op_4_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm;
  reg alu_loop_op_4_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm_2;
  reg alu_loop_op_4_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm;
  reg alu_loop_op_4_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm_2;
  reg alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm;
  reg [7:0] alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_1_itm;
  reg [7:0] alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_1_itm_2;
  reg alu_loop_op_4_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm;
  reg alu_loop_op_4_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2;
  reg alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st;
  reg alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_4_sva_st_2;
  reg FpNormalize_8U_49U_if_or_3_itm;
  reg FpNormalize_8U_49U_if_or_3_itm_2;
  reg alu_loop_op_4_FpCmp_8U_23U_true_slc_8_1_svs_st;
  reg IsNaN_8U_23U_2_land_4_lpi_1_dfm_st;
  reg alu_loop_op_4_FpCmp_8U_23U_false_slc_8_1_svs_st;
  reg FpAlu_8U_23U_and_12_itm;
  reg FpAlu_8U_23U_and_12_itm_3;
  reg FpAlu_8U_23U_and_12_itm_4;
  reg FpAlu_8U_23U_or_837_itm_3;
  reg FpAlu_8U_23U_or_837_itm_4;
  reg FpAlu_8U_23U_or_761_itm_3;
  reg FpAlu_8U_23U_or_838_itm;
  reg FpAlu_8U_23U_or_762_itm;
  reg alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_or_itm;
  reg alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
  reg alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  reg alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  reg [7:0] alu_loop_op_5_FpAdd_8U_23U_a_left_shift_acc_itm;
  reg [7:0] alu_loop_op_5_FpAdd_8U_23U_a_left_shift_acc_itm_2;
  reg alu_loop_op_5_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm;
  reg alu_loop_op_5_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2;
  reg alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm;
  reg alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2;
  reg [7:0] alu_loop_op_5_FpAdd_8U_23U_b_left_shift_acc_itm;
  reg [7:0] alu_loop_op_5_FpAdd_8U_23U_b_left_shift_acc_itm_2;
  reg alu_loop_op_5_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm;
  reg alu_loop_op_5_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2;
  reg alu_loop_op_5_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st;
  reg alu_loop_op_5_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_5_sva_st_2;
  reg FpNormalize_8U_49U_if_or_4_itm;
  reg FpNormalize_8U_49U_if_or_4_itm_2;
  reg alu_loop_op_5_FpCmp_8U_23U_true_slc_8_svs_st;
  reg IsNaN_8U_23U_2_land_5_lpi_1_dfm_st;
  reg alu_loop_op_5_FpCmp_8U_23U_false_slc_8_svs_st;
  reg FpAlu_8U_23U_and_16_itm;
  reg FpAlu_8U_23U_and_16_itm_3;
  reg FpAlu_8U_23U_and_16_itm_4;
  reg FpAlu_8U_23U_or_839_itm_3;
  reg FpAlu_8U_23U_or_839_itm_4;
  reg FpAlu_8U_23U_or_764_itm_3;
  reg FpAlu_8U_23U_or_840_itm;
  reg FpAlu_8U_23U_or_765_itm;
  reg alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_or_itm;
  reg alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
  reg alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  reg alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  reg [7:0] alu_loop_op_6_FpAdd_8U_23U_a_left_shift_acc_1_itm;
  reg [7:0] alu_loop_op_6_FpAdd_8U_23U_a_left_shift_acc_1_itm_2;
  reg alu_loop_op_6_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm;
  reg alu_loop_op_6_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2;
  reg alu_loop_op_6_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm;
  reg alu_loop_op_6_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm_2;
  reg alu_loop_op_6_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm;
  reg alu_loop_op_6_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm_2;
  reg alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm;
  reg [7:0] alu_loop_op_6_FpAdd_8U_23U_b_left_shift_acc_1_itm;
  reg [7:0] alu_loop_op_6_FpAdd_8U_23U_b_left_shift_acc_1_itm_2;
  reg alu_loop_op_6_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm;
  reg alu_loop_op_6_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2;
  reg alu_loop_op_6_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st;
  reg alu_loop_op_6_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_6_sva_st_2;
  reg FpNormalize_8U_49U_if_or_5_itm;
  reg FpNormalize_8U_49U_if_or_5_itm_2;
  reg alu_loop_op_6_FpCmp_8U_23U_true_slc_8_1_svs_st;
  reg IsNaN_8U_23U_2_land_6_lpi_1_dfm_st;
  reg alu_loop_op_6_FpCmp_8U_23U_false_slc_8_1_svs_st;
  reg FpAlu_8U_23U_and_20_itm;
  reg FpAlu_8U_23U_and_20_itm_3;
  reg FpAlu_8U_23U_and_20_itm_4;
  reg FpAlu_8U_23U_or_841_itm_3;
  reg FpAlu_8U_23U_or_841_itm_4;
  reg FpAlu_8U_23U_or_767_itm_3;
  reg FpAlu_8U_23U_or_842_itm;
  reg FpAlu_8U_23U_or_768_itm;
  reg alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_or_itm;
  reg alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
  reg alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  reg alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  reg [7:0] alu_loop_op_7_FpAdd_8U_23U_a_left_shift_acc_itm;
  reg [7:0] alu_loop_op_7_FpAdd_8U_23U_a_left_shift_acc_itm_2;
  reg alu_loop_op_7_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm;
  reg alu_loop_op_7_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2;
  reg alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm;
  reg alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3;
  reg alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4;
  reg [7:0] alu_loop_op_7_FpAdd_8U_23U_b_left_shift_acc_itm;
  reg [7:0] alu_loop_op_7_FpAdd_8U_23U_b_left_shift_acc_itm_2;
  reg alu_loop_op_7_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm;
  reg alu_loop_op_7_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2;
  reg alu_loop_op_7_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st;
  reg alu_loop_op_7_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_7_sva_st_2;
  reg FpNormalize_8U_49U_if_or_6_itm;
  reg FpNormalize_8U_49U_if_or_6_itm_2;
  reg alu_loop_op_7_FpCmp_8U_23U_true_slc_8_svs_st;
  reg IsNaN_8U_23U_2_land_7_lpi_1_dfm_st;
  reg alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_st;
  reg FpAlu_8U_23U_and_24_itm;
  reg FpAlu_8U_23U_and_24_itm_3;
  reg FpAlu_8U_23U_and_24_itm_4;
  reg FpAlu_8U_23U_or_843_itm_3;
  reg FpAlu_8U_23U_or_843_itm_4;
  reg FpAlu_8U_23U_or_770_itm_3;
  reg FpAlu_8U_23U_or_844_itm;
  reg FpAlu_8U_23U_or_771_itm;
  reg alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_or_itm;
  reg alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
  reg alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  reg alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  reg [7:0] alu_loop_op_8_FpAdd_8U_23U_a_left_shift_acc_1_itm;
  reg [7:0] alu_loop_op_8_FpAdd_8U_23U_a_left_shift_acc_1_itm_2;
  reg alu_loop_op_8_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm;
  reg alu_loop_op_8_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2;
  reg alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm;
  reg alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3;
  reg alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4;
  reg [7:0] alu_loop_op_8_FpAdd_8U_23U_b_left_shift_acc_1_itm;
  reg [7:0] alu_loop_op_8_FpAdd_8U_23U_b_left_shift_acc_1_itm_2;
  reg alu_loop_op_8_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm;
  reg alu_loop_op_8_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2;
  reg alu_loop_op_8_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st;
  reg alu_loop_op_8_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_8_sva_st_2;
  reg FpNormalize_8U_49U_if_or_7_itm;
  reg FpNormalize_8U_49U_if_or_7_itm_2;
  reg alu_loop_op_8_FpCmp_8U_23U_true_slc_8_1_svs_st;
  reg IsNaN_8U_23U_2_land_8_lpi_1_dfm_st;
  reg alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_st;
  reg FpAlu_8U_23U_and_28_itm;
  reg FpAlu_8U_23U_and_28_itm_3;
  reg FpAlu_8U_23U_and_28_itm_4;
  reg FpAlu_8U_23U_or_845_itm_3;
  reg FpAlu_8U_23U_or_845_itm_4;
  reg FpAlu_8U_23U_or_773_itm_3;
  reg FpAlu_8U_23U_or_846_itm;
  reg FpAlu_8U_23U_or_774_itm;
  reg alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_or_itm;
  reg alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
  reg alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  reg alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  reg [7:0] alu_loop_op_9_FpAdd_8U_23U_a_left_shift_acc_itm;
  reg [7:0] alu_loop_op_9_FpAdd_8U_23U_a_left_shift_acc_itm_2;
  reg alu_loop_op_9_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm;
  reg alu_loop_op_9_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2;
  reg alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm;
  reg alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2;
  reg [7:0] alu_loop_op_9_FpAdd_8U_23U_b_left_shift_acc_itm;
  reg [7:0] alu_loop_op_9_FpAdd_8U_23U_b_left_shift_acc_itm_2;
  reg alu_loop_op_9_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm;
  reg alu_loop_op_9_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2;
  reg alu_loop_op_9_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st;
  reg alu_loop_op_9_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_9_sva_st_2;
  reg FpNormalize_8U_49U_if_or_8_itm;
  reg FpNormalize_8U_49U_if_or_8_itm_2;
  reg alu_loop_op_9_FpCmp_8U_23U_true_slc_8_svs_st;
  reg IsNaN_8U_23U_2_land_9_lpi_1_dfm_st;
  reg alu_loop_op_9_FpCmp_8U_23U_false_slc_8_svs_st;
  reg FpAlu_8U_23U_and_32_itm;
  reg FpAlu_8U_23U_and_32_itm_3;
  reg FpAlu_8U_23U_and_32_itm_4;
  reg FpAlu_8U_23U_or_847_itm_3;
  reg FpAlu_8U_23U_or_847_itm_4;
  reg FpAlu_8U_23U_or_776_itm_3;
  reg FpAlu_8U_23U_or_848_itm;
  reg FpAlu_8U_23U_or_777_itm;
  reg alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_or_itm;
  reg alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
  reg alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  reg alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  reg [7:0] alu_loop_op_10_FpAdd_8U_23U_a_left_shift_acc_1_itm;
  reg [7:0] alu_loop_op_10_FpAdd_8U_23U_a_left_shift_acc_1_itm_2;
  reg alu_loop_op_10_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm;
  reg alu_loop_op_10_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2;
  reg alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm;
  reg alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2;
  reg [7:0] alu_loop_op_10_FpAdd_8U_23U_b_left_shift_acc_1_itm;
  reg [7:0] alu_loop_op_10_FpAdd_8U_23U_b_left_shift_acc_1_itm_2;
  reg alu_loop_op_10_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm;
  reg alu_loop_op_10_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2;
  reg alu_loop_op_10_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st;
  reg alu_loop_op_10_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_10_sva_st_2;
  reg FpNormalize_8U_49U_if_or_9_itm;
  reg FpNormalize_8U_49U_if_or_9_itm_2;
  reg alu_loop_op_10_FpCmp_8U_23U_true_slc_8_1_svs_st;
  reg IsNaN_8U_23U_2_land_10_lpi_1_dfm_st;
  reg alu_loop_op_10_FpCmp_8U_23U_false_slc_8_1_svs_st;
  reg FpAlu_8U_23U_and_36_itm;
  reg FpAlu_8U_23U_and_36_itm_3;
  reg FpAlu_8U_23U_and_36_itm_4;
  reg FpAlu_8U_23U_or_849_itm_3;
  reg FpAlu_8U_23U_or_849_itm_4;
  reg FpAlu_8U_23U_or_779_itm_3;
  reg FpAlu_8U_23U_or_850_itm;
  reg FpAlu_8U_23U_or_780_itm;
  reg alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_or_itm;
  reg alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
  reg alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  reg alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  reg [7:0] alu_loop_op_11_FpAdd_8U_23U_a_left_shift_acc_itm;
  reg [7:0] alu_loop_op_11_FpAdd_8U_23U_a_left_shift_acc_itm_2;
  reg alu_loop_op_11_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm;
  reg alu_loop_op_11_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2;
  reg alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm;
  reg alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2;
  reg [7:0] alu_loop_op_11_FpAdd_8U_23U_b_left_shift_acc_itm;
  reg [7:0] alu_loop_op_11_FpAdd_8U_23U_b_left_shift_acc_itm_2;
  reg alu_loop_op_11_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm;
  reg alu_loop_op_11_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2;
  reg alu_loop_op_11_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st;
  reg alu_loop_op_11_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_11_sva_st_2;
  reg FpNormalize_8U_49U_if_or_10_itm;
  reg FpNormalize_8U_49U_if_or_10_itm_2;
  reg alu_loop_op_11_FpCmp_8U_23U_true_slc_8_svs_st;
  reg IsNaN_8U_23U_2_land_11_lpi_1_dfm_st;
  reg alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_st;
  reg FpAlu_8U_23U_and_40_itm;
  reg FpAlu_8U_23U_and_40_itm_3;
  reg FpAlu_8U_23U_and_40_itm_4;
  reg FpAlu_8U_23U_or_851_itm_3;
  reg FpAlu_8U_23U_or_851_itm_4;
  reg FpAlu_8U_23U_or_782_itm_3;
  reg FpAlu_8U_23U_or_852_itm;
  reg FpAlu_8U_23U_or_783_itm;
  reg alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_or_itm;
  reg alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
  reg alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  reg alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  reg [7:0] alu_loop_op_12_FpAdd_8U_23U_a_left_shift_acc_1_itm;
  reg [7:0] alu_loop_op_12_FpAdd_8U_23U_a_left_shift_acc_1_itm_2;
  reg alu_loop_op_12_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm;
  reg alu_loop_op_12_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2;
  reg alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm;
  reg alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2;
  reg [7:0] alu_loop_op_12_FpAdd_8U_23U_b_left_shift_acc_1_itm;
  reg [7:0] alu_loop_op_12_FpAdd_8U_23U_b_left_shift_acc_1_itm_2;
  reg alu_loop_op_12_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm;
  reg alu_loop_op_12_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2;
  reg alu_loop_op_12_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st;
  reg alu_loop_op_12_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_12_sva_st_2;
  reg FpNormalize_8U_49U_if_or_11_itm;
  reg FpNormalize_8U_49U_if_or_11_itm_2;
  reg alu_loop_op_12_FpCmp_8U_23U_true_slc_8_1_svs_st;
  reg IsNaN_8U_23U_2_land_12_lpi_1_dfm_st;
  reg alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_st;
  reg FpAlu_8U_23U_and_44_itm;
  reg FpAlu_8U_23U_and_44_itm_3;
  reg FpAlu_8U_23U_and_44_itm_4;
  reg FpAlu_8U_23U_or_853_itm_3;
  reg FpAlu_8U_23U_or_853_itm_4;
  reg FpAlu_8U_23U_or_785_itm_3;
  reg FpAlu_8U_23U_or_854_itm;
  reg FpAlu_8U_23U_or_786_itm;
  reg alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_or_itm;
  reg alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
  reg alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  reg alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  reg [7:0] alu_loop_op_13_FpAdd_8U_23U_a_left_shift_acc_itm;
  reg [7:0] alu_loop_op_13_FpAdd_8U_23U_a_left_shift_acc_itm_2;
  reg alu_loop_op_13_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm;
  reg alu_loop_op_13_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2;
  reg alu_loop_op_13_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_itm;
  reg alu_loop_op_13_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_itm_2;
  reg alu_loop_op_13_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_itm;
  reg alu_loop_op_13_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_itm_2;
  reg alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm;
  reg [7:0] alu_loop_op_13_FpAdd_8U_23U_b_left_shift_acc_itm;
  reg [7:0] alu_loop_op_13_FpAdd_8U_23U_b_left_shift_acc_itm_2;
  reg alu_loop_op_13_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm;
  reg alu_loop_op_13_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2;
  reg alu_loop_op_13_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st;
  reg alu_loop_op_13_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_13_sva_st_2;
  reg FpNormalize_8U_49U_if_or_12_itm;
  reg FpNormalize_8U_49U_if_or_12_itm_2;
  reg alu_loop_op_13_FpCmp_8U_23U_true_slc_8_svs_st;
  reg IsNaN_8U_23U_2_land_13_lpi_1_dfm_st;
  reg alu_loop_op_13_FpCmp_8U_23U_false_slc_8_svs_st;
  reg FpAlu_8U_23U_and_48_itm;
  reg FpAlu_8U_23U_and_48_itm_3;
  reg FpAlu_8U_23U_and_48_itm_4;
  reg FpAlu_8U_23U_or_855_itm_3;
  reg FpAlu_8U_23U_or_855_itm_4;
  reg FpAlu_8U_23U_or_788_itm_3;
  reg FpAlu_8U_23U_or_856_itm;
  reg FpAlu_8U_23U_or_789_itm;
  reg alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_or_itm;
  reg alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
  reg alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  reg alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  reg [7:0] alu_loop_op_14_FpAdd_8U_23U_a_left_shift_acc_1_itm;
  reg [7:0] alu_loop_op_14_FpAdd_8U_23U_a_left_shift_acc_1_itm_2;
  reg alu_loop_op_14_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm;
  reg alu_loop_op_14_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2;
  reg alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm;
  reg alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2;
  reg [7:0] alu_loop_op_14_FpAdd_8U_23U_b_left_shift_acc_1_itm;
  reg [7:0] alu_loop_op_14_FpAdd_8U_23U_b_left_shift_acc_1_itm_2;
  reg alu_loop_op_14_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm;
  reg alu_loop_op_14_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2;
  reg alu_loop_op_14_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st;
  reg alu_loop_op_14_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_14_sva_st_2;
  reg FpNormalize_8U_49U_if_or_13_itm;
  reg FpNormalize_8U_49U_if_or_13_itm_2;
  reg alu_loop_op_14_FpCmp_8U_23U_true_slc_8_1_svs_st;
  reg IsNaN_8U_23U_2_land_14_lpi_1_dfm_st;
  reg alu_loop_op_14_FpCmp_8U_23U_false_slc_8_1_svs_st;
  reg FpAlu_8U_23U_and_52_itm;
  reg FpAlu_8U_23U_and_52_itm_3;
  reg FpAlu_8U_23U_and_52_itm_4;
  reg FpAlu_8U_23U_or_857_itm_3;
  reg FpAlu_8U_23U_or_857_itm_4;
  reg FpAlu_8U_23U_or_791_itm_3;
  reg FpAlu_8U_23U_or_858_itm;
  reg FpAlu_8U_23U_or_792_itm;
  reg alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_or_itm;
  reg alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
  reg alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  reg alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  reg [7:0] alu_loop_op_15_FpAdd_8U_23U_a_left_shift_acc_itm;
  reg [7:0] alu_loop_op_15_FpAdd_8U_23U_a_left_shift_acc_itm_2;
  reg alu_loop_op_15_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm;
  reg alu_loop_op_15_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2;
  reg alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm;
  reg alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3;
  reg alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4;
  reg [7:0] alu_loop_op_15_FpAdd_8U_23U_b_left_shift_acc_itm;
  reg [7:0] alu_loop_op_15_FpAdd_8U_23U_b_left_shift_acc_itm_2;
  reg alu_loop_op_15_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm;
  reg alu_loop_op_15_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2;
  reg alu_loop_op_15_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st;
  reg alu_loop_op_15_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_15_sva_st_2;
  reg FpNormalize_8U_49U_if_or_14_itm;
  reg FpNormalize_8U_49U_if_or_14_itm_2;
  reg alu_loop_op_15_FpCmp_8U_23U_true_slc_8_svs_st;
  reg IsNaN_8U_23U_2_land_15_lpi_1_dfm_st;
  reg alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_st;
  reg FpAlu_8U_23U_and_56_itm;
  reg FpAlu_8U_23U_and_56_itm_3;
  reg FpAlu_8U_23U_and_56_itm_4;
  reg FpAlu_8U_23U_or_859_itm_3;
  reg FpAlu_8U_23U_or_859_itm_4;
  reg FpAlu_8U_23U_or_794_itm_3;
  reg FpAlu_8U_23U_or_860_itm;
  reg FpAlu_8U_23U_or_795_itm;
  reg [1:0] cfg_alu_algo_1_sva_st_15;
  reg alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_or_itm;
  reg alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
  reg alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  reg alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  reg [7:0] alu_loop_op_16_FpAdd_8U_23U_a_left_shift_acc_1_itm;
  reg [7:0] alu_loop_op_16_FpAdd_8U_23U_a_left_shift_acc_1_itm_2;
  reg alu_loop_op_16_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm;
  reg alu_loop_op_16_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2;
  reg alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm;
  reg alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3;
  reg alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4;
  reg [7:0] alu_loop_op_16_FpAdd_8U_23U_b_left_shift_acc_1_itm;
  reg [7:0] alu_loop_op_16_FpAdd_8U_23U_b_left_shift_acc_1_itm_2;
  reg alu_loop_op_16_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm;
  reg alu_loop_op_16_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2;
  reg alu_loop_op_16_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st;
  reg alu_loop_op_16_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_st_2;
  reg FpNormalize_8U_49U_if_or_15_itm;
  reg FpNormalize_8U_49U_if_or_15_itm_2;
  reg alu_loop_op_16_FpCmp_8U_23U_true_slc_8_1_svs_st;
  reg IsNaN_8U_23U_2_land_lpi_1_dfm_st;
  reg alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_st;
  reg FpAlu_8U_23U_and_60_itm;
  reg FpAlu_8U_23U_and_60_itm_3;
  reg FpAlu_8U_23U_and_60_itm_4;
  reg FpAlu_8U_23U_or_861_itm_3;
  reg FpAlu_8U_23U_or_861_itm_4;
  reg FpAlu_8U_23U_or_797_itm_3;
  reg FpAlu_8U_23U_or_862_itm;
  reg FpAlu_8U_23U_or_798_itm;
  reg alu_loop_op_else_if_mux_itm;
  reg [29:0] alu_loop_op_else_if_mux_1_itm;
  reg alu_loop_op_else_if_mux_2_itm;
  reg alu_loop_op_else_else_if_mux_itm;
  reg alu_loop_op_else_else_if_mux_itm_2;
  reg [29:0] alu_loop_op_else_else_if_mux_1_itm;
  reg [29:0] alu_loop_op_else_else_if_mux_1_itm_2;
  reg alu_loop_op_else_else_if_mux_2_itm;
  reg alu_loop_op_else_else_if_mux_2_itm_2;
  reg alu_loop_op_else_if_mux_3_itm;
  reg [29:0] alu_loop_op_else_if_mux_4_itm;
  reg alu_loop_op_else_if_mux_5_itm;
  reg alu_loop_op_else_else_if_mux_3_itm;
  reg alu_loop_op_else_else_if_mux_3_itm_2;
  reg [29:0] alu_loop_op_else_else_if_mux_4_itm;
  reg [29:0] alu_loop_op_else_else_if_mux_4_itm_2;
  reg alu_loop_op_else_else_if_mux_5_itm;
  reg alu_loop_op_else_else_if_mux_5_itm_2;
  reg alu_loop_op_else_if_mux_6_itm;
  reg [29:0] alu_loop_op_else_if_mux_7_itm;
  reg alu_loop_op_else_if_mux_8_itm;
  reg alu_loop_op_else_else_if_mux_6_itm;
  reg alu_loop_op_else_else_if_mux_6_itm_3;
  reg alu_loop_op_else_else_if_mux_6_itm_4;
  reg [29:0] alu_loop_op_else_else_if_mux_7_itm;
  reg [29:0] alu_loop_op_else_else_if_mux_7_itm_3;
  reg [29:0] alu_loop_op_else_else_if_mux_7_itm_4;
  reg alu_loop_op_else_else_if_mux_8_itm;
  reg alu_loop_op_else_else_if_mux_8_itm_3;
  reg alu_loop_op_else_else_if_mux_8_itm_4;
  reg alu_loop_op_else_if_mux_9_itm;
  reg [29:0] alu_loop_op_else_if_mux_10_itm;
  reg alu_loop_op_else_if_mux_11_itm;
  reg alu_loop_op_else_else_if_mux_9_itm;
  reg alu_loop_op_else_else_if_mux_9_itm_2;
  reg [29:0] alu_loop_op_else_else_if_mux_10_itm;
  reg [29:0] alu_loop_op_else_else_if_mux_10_itm_2;
  reg alu_loop_op_else_else_if_mux_11_itm;
  reg alu_loop_op_else_else_if_mux_11_itm_2;
  reg alu_loop_op_else_if_mux_12_itm;
  reg [29:0] alu_loop_op_else_if_mux_13_itm;
  reg alu_loop_op_else_if_mux_14_itm;
  reg alu_loop_op_else_else_if_mux_12_itm;
  reg alu_loop_op_else_else_if_mux_12_itm_3;
  reg alu_loop_op_else_else_if_mux_12_itm_4;
  reg [29:0] alu_loop_op_else_else_if_mux_13_itm;
  reg [29:0] alu_loop_op_else_else_if_mux_13_itm_3;
  reg [29:0] alu_loop_op_else_else_if_mux_13_itm_4;
  reg alu_loop_op_else_else_if_mux_14_itm;
  reg alu_loop_op_else_else_if_mux_14_itm_3;
  reg alu_loop_op_else_else_if_mux_14_itm_4;
  reg alu_loop_op_else_if_mux_15_itm;
  reg [29:0] alu_loop_op_else_if_mux_16_itm;
  reg alu_loop_op_else_if_mux_17_itm;
  reg alu_loop_op_else_else_if_mux_15_itm;
  reg alu_loop_op_else_else_if_mux_15_itm_3;
  reg alu_loop_op_else_else_if_mux_15_itm_4;
  reg [29:0] alu_loop_op_else_else_if_mux_16_itm;
  reg [29:0] alu_loop_op_else_else_if_mux_16_itm_3;
  reg [29:0] alu_loop_op_else_else_if_mux_16_itm_4;
  reg alu_loop_op_else_else_if_mux_17_itm;
  reg alu_loop_op_else_else_if_mux_17_itm_3;
  reg alu_loop_op_else_else_if_mux_17_itm_4;
  reg alu_loop_op_else_if_mux_18_itm;
  reg [29:0] alu_loop_op_else_if_mux_19_itm;
  reg alu_loop_op_else_if_mux_20_itm;
  reg alu_loop_op_else_else_if_mux_18_itm;
  reg alu_loop_op_else_else_if_mux_18_itm_3;
  reg alu_loop_op_else_else_if_mux_18_itm_4;
  reg [29:0] alu_loop_op_else_else_if_mux_19_itm;
  reg [29:0] alu_loop_op_else_else_if_mux_19_itm_3;
  reg [29:0] alu_loop_op_else_else_if_mux_19_itm_4;
  reg alu_loop_op_else_else_if_mux_20_itm;
  reg alu_loop_op_else_else_if_mux_20_itm_3;
  reg alu_loop_op_else_else_if_mux_20_itm_4;
  reg alu_loop_op_else_if_mux_21_itm;
  reg [29:0] alu_loop_op_else_if_mux_22_itm;
  reg alu_loop_op_else_if_mux_23_itm;
  reg alu_loop_op_else_else_if_mux_21_itm;
  reg alu_loop_op_else_else_if_mux_21_itm_3;
  reg alu_loop_op_else_else_if_mux_21_itm_4;
  reg [29:0] alu_loop_op_else_else_if_mux_22_itm;
  reg [29:0] alu_loop_op_else_else_if_mux_22_itm_3;
  reg [29:0] alu_loop_op_else_else_if_mux_22_itm_4;
  reg alu_loop_op_else_else_if_mux_23_itm;
  reg alu_loop_op_else_else_if_mux_23_itm_3;
  reg alu_loop_op_else_else_if_mux_23_itm_4;
  reg alu_loop_op_else_if_mux_24_itm;
  reg [29:0] alu_loop_op_else_if_mux_25_itm;
  reg alu_loop_op_else_if_mux_26_itm;
  reg alu_loop_op_else_else_if_mux_24_itm;
  reg alu_loop_op_else_else_if_mux_24_itm_3;
  reg alu_loop_op_else_else_if_mux_24_itm_4;
  reg [29:0] alu_loop_op_else_else_if_mux_25_itm;
  reg [29:0] alu_loop_op_else_else_if_mux_25_itm_3;
  reg [29:0] alu_loop_op_else_else_if_mux_25_itm_4;
  reg alu_loop_op_else_else_if_mux_26_itm;
  reg alu_loop_op_else_else_if_mux_26_itm_3;
  reg alu_loop_op_else_else_if_mux_26_itm_4;
  reg alu_loop_op_else_if_mux_27_itm;
  reg [29:0] alu_loop_op_else_if_mux_28_itm;
  reg alu_loop_op_else_if_mux_29_itm;
  reg alu_loop_op_else_else_if_mux_27_itm;
  reg alu_loop_op_else_else_if_mux_27_itm_3;
  reg alu_loop_op_else_else_if_mux_27_itm_4;
  reg [29:0] alu_loop_op_else_else_if_mux_28_itm;
  reg [29:0] alu_loop_op_else_else_if_mux_28_itm_3;
  reg [29:0] alu_loop_op_else_else_if_mux_28_itm_4;
  reg alu_loop_op_else_else_if_mux_29_itm;
  reg alu_loop_op_else_else_if_mux_29_itm_3;
  reg alu_loop_op_else_else_if_mux_29_itm_4;
  reg alu_loop_op_else_if_mux_30_itm;
  reg [29:0] alu_loop_op_else_if_mux_31_itm;
  reg alu_loop_op_else_if_mux_32_itm;
  reg alu_loop_op_else_else_if_mux_30_itm;
  reg alu_loop_op_else_else_if_mux_30_itm_3;
  reg alu_loop_op_else_else_if_mux_30_itm_4;
  reg [29:0] alu_loop_op_else_else_if_mux_31_itm;
  reg [29:0] alu_loop_op_else_else_if_mux_31_itm_3;
  reg [29:0] alu_loop_op_else_else_if_mux_31_itm_4;
  reg alu_loop_op_else_else_if_mux_32_itm;
  reg alu_loop_op_else_else_if_mux_32_itm_3;
  reg alu_loop_op_else_else_if_mux_32_itm_4;
  reg alu_loop_op_else_if_mux_33_itm;
  reg [29:0] alu_loop_op_else_if_mux_34_itm;
  reg alu_loop_op_else_if_mux_35_itm;
  reg alu_loop_op_else_else_if_mux_33_itm;
  reg alu_loop_op_else_else_if_mux_33_itm_3;
  reg alu_loop_op_else_else_if_mux_33_itm_4;
  reg [29:0] alu_loop_op_else_else_if_mux_34_itm;
  reg [29:0] alu_loop_op_else_else_if_mux_34_itm_3;
  reg [29:0] alu_loop_op_else_else_if_mux_34_itm_4;
  reg alu_loop_op_else_else_if_mux_35_itm;
  reg alu_loop_op_else_else_if_mux_35_itm_3;
  reg alu_loop_op_else_else_if_mux_35_itm_4;
  reg alu_loop_op_else_if_mux_36_itm;
  reg [29:0] alu_loop_op_else_if_mux_37_itm;
  reg alu_loop_op_else_if_mux_38_itm;
  reg alu_loop_op_else_else_if_mux_36_itm;
  reg alu_loop_op_else_else_if_mux_36_itm_3;
  reg alu_loop_op_else_else_if_mux_36_itm_4;
  reg [29:0] alu_loop_op_else_else_if_mux_37_itm;
  reg [29:0] alu_loop_op_else_else_if_mux_37_itm_3;
  reg [29:0] alu_loop_op_else_else_if_mux_37_itm_4;
  reg alu_loop_op_else_else_if_mux_38_itm;
  reg alu_loop_op_else_else_if_mux_38_itm_3;
  reg alu_loop_op_else_else_if_mux_38_itm_4;
  reg alu_loop_op_else_if_mux_39_itm;
  reg [29:0] alu_loop_op_else_if_mux_40_itm;
  reg alu_loop_op_else_if_mux_41_itm;
  reg alu_loop_op_else_else_if_mux_39_itm;
  reg alu_loop_op_else_else_if_mux_39_itm_3;
  reg alu_loop_op_else_else_if_mux_39_itm_4;
  reg [29:0] alu_loop_op_else_else_if_mux_40_itm;
  reg [29:0] alu_loop_op_else_else_if_mux_40_itm_3;
  reg [29:0] alu_loop_op_else_else_if_mux_40_itm_4;
  reg alu_loop_op_else_else_if_mux_41_itm;
  reg alu_loop_op_else_else_if_mux_41_itm_3;
  reg alu_loop_op_else_else_if_mux_41_itm_4;
  reg alu_loop_op_else_if_mux_42_itm;
  reg [29:0] alu_loop_op_else_if_mux_43_itm;
  reg alu_loop_op_else_if_mux_44_itm;
  reg alu_loop_op_else_else_if_mux_42_itm;
  reg alu_loop_op_else_else_if_mux_42_itm_3;
  reg alu_loop_op_else_else_if_mux_42_itm_4;
  reg [29:0] alu_loop_op_else_else_if_mux_43_itm;
  reg [29:0] alu_loop_op_else_else_if_mux_43_itm_3;
  reg [29:0] alu_loop_op_else_else_if_mux_43_itm_4;
  reg alu_loop_op_else_else_if_mux_44_itm;
  reg alu_loop_op_else_else_if_mux_44_itm_3;
  reg alu_loop_op_else_else_if_mux_44_itm_4;
  reg [1:0] cfg_alu_algo_1_sva_st_31;
  reg alu_loop_op_else_if_mux_45_itm;
  reg [29:0] alu_loop_op_else_if_mux_46_itm;
  reg alu_loop_op_else_if_mux_47_itm;
  reg alu_loop_op_else_else_if_mux_45_itm;
  reg alu_loop_op_else_else_if_mux_45_itm_3;
  reg alu_loop_op_else_else_if_mux_45_itm_4;
  reg [29:0] alu_loop_op_else_else_if_mux_46_itm;
  reg [29:0] alu_loop_op_else_else_if_mux_46_itm_3;
  reg [29:0] alu_loop_op_else_else_if_mux_46_itm_4;
  reg alu_loop_op_else_else_if_mux_47_itm;
  reg alu_loop_op_else_else_if_mux_47_itm_3;
  reg alu_loop_op_else_else_if_mux_47_itm_4;
  reg io_read_cfg_alu_bypass_rsc_svs_st_1;
  reg cfg_alu_src_1_sva_st_1;
  reg io_read_cfg_alu_bypass_rsc_svs_st_5;
  reg io_read_cfg_alu_bypass_rsc_svs_st_6;
  reg alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_st_3;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_2_land_1_lpi_1_dfm_st_1;
  reg alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_st_2;
  reg alu_loop_op_2_FpAdd_8U_23U_is_a_greater_slc_8_1_svs_st_2;
  reg alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_st_2;
  reg alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_st_3;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_2_land_2_lpi_1_dfm_st_1;
  reg alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_st_2;
  reg alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_st_3;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_2_land_3_lpi_1_dfm_st_1;
  reg alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_st_2;
  reg alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_4_sva_st_3;
  reg IsNaN_8U_23U_land_4_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_2_land_4_lpi_1_dfm_st_1;
  reg alu_loop_op_4_FpCmp_8U_23U_false_slc_8_1_svs_st_2;
  reg alu_loop_op_5_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_5_sva_st_3;
  reg IsNaN_8U_23U_land_5_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_2_land_5_lpi_1_dfm_st_1;
  reg alu_loop_op_5_FpCmp_8U_23U_false_slc_8_svs_st_2;
  reg alu_loop_op_6_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_6_sva_st_3;
  reg IsNaN_8U_23U_land_6_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_2_land_6_lpi_1_dfm_st_1;
  reg alu_loop_op_6_FpCmp_8U_23U_false_slc_8_1_svs_st_2;
  reg alu_loop_op_7_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_7_sva_st_3;
  reg IsNaN_8U_23U_land_7_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_2_land_7_lpi_1_dfm_st_1;
  reg alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_st_2;
  reg alu_loop_op_8_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_8_sva_st_3;
  reg IsNaN_8U_23U_land_8_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_2_land_8_lpi_1_dfm_st_1;
  reg alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_st_2;
  reg alu_loop_op_9_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_9_sva_st_3;
  reg IsNaN_8U_23U_land_9_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_2_land_9_lpi_1_dfm_st_1;
  reg alu_loop_op_9_FpCmp_8U_23U_false_slc_8_svs_st_2;
  reg alu_loop_op_10_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_10_sva_st_3;
  reg IsNaN_8U_23U_land_10_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_2_land_10_lpi_1_dfm_st_1;
  reg alu_loop_op_10_FpCmp_8U_23U_false_slc_8_1_svs_st_2;
  reg alu_loop_op_11_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_11_sva_st_3;
  reg IsNaN_8U_23U_land_11_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_2_land_11_lpi_1_dfm_st_1;
  reg alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_st_2;
  reg alu_loop_op_12_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_12_sva_st_3;
  reg IsNaN_8U_23U_land_12_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_2_land_12_lpi_1_dfm_st_1;
  reg alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_st_2;
  reg alu_loop_op_13_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_13_sva_st_3;
  reg IsNaN_8U_23U_land_13_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_2_land_13_lpi_1_dfm_st_1;
  reg alu_loop_op_13_FpCmp_8U_23U_false_slc_8_svs_st_2;
  reg alu_loop_op_14_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_14_sva_st_3;
  reg IsNaN_8U_23U_land_14_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_2_land_14_lpi_1_dfm_st_1;
  reg alu_loop_op_14_FpCmp_8U_23U_false_slc_8_1_svs_st_2;
  reg alu_loop_op_15_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_15_sva_st_3;
  reg IsNaN_8U_23U_land_15_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_2_land_15_lpi_1_dfm_st_1;
  reg alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_st_2;
  reg [1:0] cfg_alu_algo_1_sva_st_92;
  reg [1:0] cfg_alu_algo_1_sva_st_204;
  reg [1:0] cfg_alu_algo_1_sva_st_205;
  reg alu_loop_op_16_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_st_3;
  reg IsNaN_8U_23U_land_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_2_land_lpi_1_dfm_st_1;
  reg alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_st_2;
  reg [1:0] cfg_alu_algo_1_sva_st_96;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_9_0;
  reg [3:0] FpAdd_8U_23U_qr_2_lpi_1_dfm_7_4;
  reg [3:0] FpAdd_8U_23U_qr_2_lpi_1_dfm_3_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_9_0;
  reg [3:0] FpAdd_8U_23U_qr_3_lpi_1_dfm_7_4;
  reg [3:0] FpAdd_8U_23U_qr_3_lpi_1_dfm_3_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_9_0;
  reg [3:0] FpAdd_8U_23U_qr_4_lpi_1_dfm_7_4;
  reg [3:0] FpAdd_8U_23U_qr_4_lpi_1_dfm_3_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_9_0;
  reg [3:0] FpAdd_8U_23U_qr_5_lpi_1_dfm_7_4;
  reg [3:0] FpAdd_8U_23U_qr_5_lpi_1_dfm_3_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_9_0;
  reg [3:0] FpAdd_8U_23U_qr_6_lpi_1_dfm_7_4;
  reg [3:0] FpAdd_8U_23U_qr_6_lpi_1_dfm_3_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_9_0;
  reg [3:0] FpAdd_8U_23U_qr_7_lpi_1_dfm_7_4;
  reg [3:0] FpAdd_8U_23U_qr_7_lpi_1_dfm_3_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_9_0;
  reg [3:0] FpAdd_8U_23U_qr_8_lpi_1_dfm_7_4;
  reg [3:0] FpAdd_8U_23U_qr_8_lpi_1_dfm_3_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_9_0;
  reg [3:0] FpAdd_8U_23U_qr_9_lpi_1_dfm_7_4;
  reg [3:0] FpAdd_8U_23U_qr_9_lpi_1_dfm_3_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_9_0;
  reg [3:0] FpAdd_8U_23U_qr_10_lpi_1_dfm_7_4;
  reg [3:0] FpAdd_8U_23U_qr_10_lpi_1_dfm_3_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_9_0;
  reg [3:0] FpAdd_8U_23U_qr_11_lpi_1_dfm_7_4;
  reg [3:0] FpAdd_8U_23U_qr_11_lpi_1_dfm_3_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_9_0;
  reg [3:0] FpAdd_8U_23U_qr_12_lpi_1_dfm_7_4;
  reg [3:0] FpAdd_8U_23U_qr_12_lpi_1_dfm_3_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_9_0;
  reg [3:0] FpAdd_8U_23U_qr_13_lpi_1_dfm_7_4;
  reg [3:0] FpAdd_8U_23U_qr_13_lpi_1_dfm_3_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_9_0;
  reg [3:0] FpAdd_8U_23U_qr_14_lpi_1_dfm_7_4;
  reg [3:0] FpAdd_8U_23U_qr_14_lpi_1_dfm_3_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_9_0;
  reg [3:0] FpAdd_8U_23U_qr_15_lpi_1_dfm_7_4;
  reg [3:0] FpAdd_8U_23U_qr_15_lpi_1_dfm_3_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_9_0;
  reg [3:0] FpAdd_8U_23U_qr_16_lpi_1_dfm_7_4;
  reg [3:0] FpAdd_8U_23U_qr_16_lpi_1_dfm_3_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_9_0;
  reg [3:0] FpAdd_8U_23U_qr_lpi_1_dfm_7_4;
  reg [3:0] FpAdd_8U_23U_qr_lpi_1_dfm_3_0;
  reg [3:0] FpAdd_8U_23U_qr_2_lpi_1_dfm_4_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_2_lpi_1_dfm_4_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_2_lpi_1_dfm_5_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_2_lpi_1_dfm_5_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_3_lpi_1_dfm_4_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_3_lpi_1_dfm_4_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_3_lpi_1_dfm_5_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_3_lpi_1_dfm_5_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_4_lpi_1_dfm_4_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_4_lpi_1_dfm_4_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_4_lpi_1_dfm_5_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_4_lpi_1_dfm_5_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_5_lpi_1_dfm_4_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_5_lpi_1_dfm_4_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_5_lpi_1_dfm_5_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_5_lpi_1_dfm_5_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_6_lpi_1_dfm_4_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_6_lpi_1_dfm_4_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_6_lpi_1_dfm_5_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_6_lpi_1_dfm_5_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_7_lpi_1_dfm_4_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_7_lpi_1_dfm_4_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_7_lpi_1_dfm_5_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_7_lpi_1_dfm_5_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_8_lpi_1_dfm_4_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_8_lpi_1_dfm_4_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_8_lpi_1_dfm_5_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_8_lpi_1_dfm_5_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_9_lpi_1_dfm_4_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_9_lpi_1_dfm_4_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_9_lpi_1_dfm_5_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_9_lpi_1_dfm_5_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_10_lpi_1_dfm_4_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_10_lpi_1_dfm_4_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_10_lpi_1_dfm_5_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_10_lpi_1_dfm_5_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_11_lpi_1_dfm_4_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_11_lpi_1_dfm_4_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_11_lpi_1_dfm_5_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_11_lpi_1_dfm_5_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_12_lpi_1_dfm_4_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_12_lpi_1_dfm_4_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_12_lpi_1_dfm_5_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_12_lpi_1_dfm_5_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_13_lpi_1_dfm_4_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_13_lpi_1_dfm_4_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_13_lpi_1_dfm_5_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_13_lpi_1_dfm_5_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_14_lpi_1_dfm_4_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_14_lpi_1_dfm_4_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_14_lpi_1_dfm_5_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_14_lpi_1_dfm_5_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_15_lpi_1_dfm_4_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_15_lpi_1_dfm_4_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_15_lpi_1_dfm_5_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_15_lpi_1_dfm_5_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_16_lpi_1_dfm_4_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_16_lpi_1_dfm_4_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_16_lpi_1_dfm_5_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_16_lpi_1_dfm_5_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_lpi_1_dfm_4_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_lpi_1_dfm_4_3_0_1;
  reg [3:0] FpAdd_8U_23U_qr_lpi_1_dfm_5_7_4_1;
  reg [3:0] FpAdd_8U_23U_qr_lpi_1_dfm_5_3_0_1;
  reg alu_loop_op_1_else_if_conc_itm_31;
  reg [29:0] alu_loop_op_1_else_if_conc_itm_30_1;
  reg alu_loop_op_1_else_if_conc_itm_0;
  reg alu_loop_op_1_else_else_if_conc_itm_31;
  reg [29:0] alu_loop_op_1_else_else_if_conc_itm_30_1;
  reg alu_loop_op_1_else_else_if_conc_itm_0;
  reg alu_loop_op_1_else_else_if_conc_itm_1_31_1;
  reg [29:0] alu_loop_op_1_else_else_if_conc_itm_1_30_1_1;
  reg alu_loop_op_1_else_else_if_conc_itm_1_0_1;
  reg alu_loop_op_2_else_if_conc_1_itm_31;
  reg [29:0] alu_loop_op_2_else_if_conc_1_itm_30_1;
  reg alu_loop_op_2_else_if_conc_1_itm_0;
  reg alu_loop_op_2_else_else_if_conc_1_itm_31;
  reg [29:0] alu_loop_op_2_else_else_if_conc_1_itm_30_1;
  reg alu_loop_op_2_else_else_if_conc_1_itm_0;
  reg alu_loop_op_2_else_else_if_conc_1_itm_1_31_1;
  reg [29:0] alu_loop_op_2_else_else_if_conc_1_itm_1_30_1_1;
  reg alu_loop_op_2_else_else_if_conc_1_itm_1_0_1;
  reg alu_loop_op_4_else_if_conc_1_itm_31;
  reg [29:0] alu_loop_op_4_else_if_conc_1_itm_30_1;
  reg alu_loop_op_4_else_if_conc_1_itm_0;
  reg alu_loop_op_4_else_else_if_conc_1_itm_31;
  reg [29:0] alu_loop_op_4_else_else_if_conc_1_itm_30_1;
  reg alu_loop_op_4_else_else_if_conc_1_itm_0;
  reg alu_loop_op_4_else_else_if_conc_1_itm_1_31_1;
  reg [29:0] alu_loop_op_4_else_else_if_conc_1_itm_1_30_1_1;
  reg alu_loop_op_4_else_else_if_conc_1_itm_1_0_1;
  wire FpAdd_8U_23U_mux_242_tmp_49;
  wire FpAdd_8U_23U_mux_226_tmp_49;
  wire FpAdd_8U_23U_mux_210_tmp_49;
  wire FpAdd_8U_23U_mux_194_tmp_49;
  wire FpAdd_8U_23U_mux_178_tmp_49;
  wire FpAdd_8U_23U_mux_162_tmp_49;
  wire FpAdd_8U_23U_mux_146_tmp_49;
  wire FpAdd_8U_23U_mux_130_tmp_49;
  wire FpAdd_8U_23U_mux_114_tmp_49;
  wire FpAdd_8U_23U_mux_98_tmp_49;
  wire FpAdd_8U_23U_mux_82_tmp_49;
  wire FpAdd_8U_23U_mux_66_tmp_49;
  wire FpAdd_8U_23U_mux_50_tmp_49;
  wire FpAdd_8U_23U_mux_34_tmp_49;
  wire FpAdd_8U_23U_mux_18_tmp_49;
  wire FpAdd_8U_23U_mux_2_tmp_49;
  wire IsDenorm_5U_23U_land_lpi_1_dfm;
  wire IsInf_5U_23U_land_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_15_cse;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_sva;
  wire IsDenorm_5U_23U_land_15_lpi_1_dfm;
  wire IsInf_5U_23U_land_15_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_14_cse;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_15_sva;
  wire IsDenorm_5U_23U_land_14_lpi_1_dfm;
  wire IsInf_5U_23U_land_14_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_13_cse;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_14_sva;
  wire IsDenorm_5U_23U_land_13_lpi_1_dfm;
  wire IsInf_5U_23U_land_13_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_12_cse;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_13_sva;
  wire IsDenorm_5U_23U_land_12_lpi_1_dfm;
  wire IsInf_5U_23U_land_12_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_11_cse;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_12_sva;
  wire IsDenorm_5U_23U_land_11_lpi_1_dfm;
  wire IsInf_5U_23U_land_11_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_10_cse;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_11_sva;
  wire IsDenorm_5U_23U_land_10_lpi_1_dfm;
  wire IsInf_5U_23U_land_10_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_9_cse;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_10_sva;
  wire IsDenorm_5U_23U_land_9_lpi_1_dfm;
  wire IsInf_5U_23U_land_9_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_8_cse;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_9_sva;
  wire IsDenorm_5U_23U_land_8_lpi_1_dfm;
  wire IsInf_5U_23U_land_8_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_7_cse;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_8_sva;
  wire IsDenorm_5U_23U_land_7_lpi_1_dfm;
  wire IsInf_5U_23U_land_7_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_6_cse;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_7_sva;
  wire IsDenorm_5U_23U_land_6_lpi_1_dfm;
  wire IsInf_5U_23U_land_6_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_5_cse;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_6_sva;
  wire IsDenorm_5U_23U_land_5_lpi_1_dfm;
  wire IsInf_5U_23U_land_5_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_4_cse;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_5_sva;
  wire IsDenorm_5U_23U_land_4_lpi_1_dfm;
  wire IsInf_5U_23U_land_4_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_3_cse;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_4_sva;
  wire IsDenorm_5U_23U_land_3_lpi_1_dfm;
  wire IsInf_5U_23U_land_3_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_2_cse;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_3_sva;
  wire IsDenorm_5U_23U_land_2_lpi_1_dfm;
  wire IsInf_5U_23U_land_2_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_1_cse;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_2_sva;
  wire IsDenorm_5U_23U_land_1_lpi_1_dfm;
  wire IsInf_5U_23U_land_1_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_cse;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_1_sva;
  wire [4:0] else_AluOp_data_15_14_10_lpi_1_dfm_mx0;
  wire [4:0] else_AluOp_data_14_14_10_lpi_1_dfm_mx0;
  wire [4:0] else_AluOp_data_13_14_10_lpi_1_dfm_mx0;
  wire [4:0] else_AluOp_data_12_14_10_lpi_1_dfm_mx0;
  wire [4:0] else_AluOp_data_11_14_10_lpi_1_dfm_mx0;
  wire [4:0] else_AluOp_data_10_14_10_lpi_1_dfm_mx0;
  wire [4:0] else_AluOp_data_9_14_10_lpi_1_dfm_mx0;
  wire [4:0] else_AluOp_data_8_14_10_lpi_1_dfm_mx0;
  wire [4:0] else_AluOp_data_7_14_10_lpi_1_dfm_mx0;
  wire [4:0] else_AluOp_data_6_14_10_lpi_1_dfm_mx0;
  wire [4:0] else_AluOp_data_5_14_10_lpi_1_dfm_mx0;
  wire [4:0] else_AluOp_data_4_14_10_lpi_1_dfm_mx0;
  wire [4:0] else_AluOp_data_3_14_10_lpi_1_dfm_mx0;
  wire [4:0] else_AluOp_data_2_14_10_lpi_1_dfm_mx0;
  wire [4:0] else_AluOp_data_1_14_10_lpi_1_dfm_mx0;
  wire [4:0] else_AluOp_data_0_14_10_lpi_1_dfm_mx0;
  wire and_1_m1c;
  wire alu_loop_op_else_equal_tmp;
  wire else_unequal_tmp;
  wire FpAdd_8U_23U_and_143_ssc;
  wire FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_and_47_tmp;
  wire FpAdd_8U_23U_is_inf_lpi_1_dfm;
  wire FpAdd_8U_23U_and_141_ssc;
  wire FpAdd_8U_23U_is_inf_15_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_and_46_tmp;
  wire FpAdd_8U_23U_is_inf_15_lpi_1_dfm;
  wire FpAdd_8U_23U_and_139_ssc;
  wire FpAdd_8U_23U_is_inf_14_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_and_45_tmp;
  wire FpAdd_8U_23U_is_inf_14_lpi_1_dfm;
  wire FpAdd_8U_23U_and_137_ssc;
  wire FpAdd_8U_23U_is_inf_13_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_and_44_tmp;
  wire FpAdd_8U_23U_is_inf_13_lpi_1_dfm;
  wire FpAdd_8U_23U_and_135_ssc;
  wire FpAdd_8U_23U_is_inf_12_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_and_43_tmp;
  wire FpAdd_8U_23U_is_inf_12_lpi_1_dfm;
  wire FpAdd_8U_23U_and_133_ssc;
  wire FpAdd_8U_23U_is_inf_11_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_and_42_tmp;
  wire FpAdd_8U_23U_is_inf_11_lpi_1_dfm;
  wire FpAdd_8U_23U_and_131_ssc;
  wire FpAdd_8U_23U_is_inf_10_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_and_41_tmp;
  wire FpAdd_8U_23U_is_inf_10_lpi_1_dfm;
  wire FpAdd_8U_23U_and_129_ssc;
  wire FpAdd_8U_23U_is_inf_9_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_and_40_tmp;
  wire FpAdd_8U_23U_is_inf_9_lpi_1_dfm;
  wire FpAdd_8U_23U_and_127_ssc;
  wire FpAdd_8U_23U_is_inf_8_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_and_39_tmp;
  wire FpAdd_8U_23U_is_inf_8_lpi_1_dfm;
  wire FpAdd_8U_23U_and_125_ssc;
  wire FpAdd_8U_23U_is_inf_7_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_and_38_tmp;
  wire FpAdd_8U_23U_is_inf_7_lpi_1_dfm;
  wire FpAdd_8U_23U_and_123_ssc;
  wire FpAdd_8U_23U_is_inf_6_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_and_37_tmp;
  wire FpAdd_8U_23U_is_inf_6_lpi_1_dfm;
  wire FpAdd_8U_23U_and_121_ssc;
  wire FpAdd_8U_23U_is_inf_5_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_and_36_tmp;
  wire FpAdd_8U_23U_is_inf_5_lpi_1_dfm;
  wire FpAdd_8U_23U_and_119_ssc;
  wire FpAdd_8U_23U_is_inf_4_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_and_35_tmp;
  wire FpAdd_8U_23U_is_inf_4_lpi_1_dfm;
  wire FpAdd_8U_23U_and_117_ssc;
  wire FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_and_34_tmp;
  wire FpAdd_8U_23U_is_inf_3_lpi_1_dfm;
  wire FpAdd_8U_23U_and_115_ssc;
  wire FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_and_33_tmp;
  wire FpAdd_8U_23U_is_inf_2_lpi_1_dfm;
  wire FpAdd_8U_23U_and_113_ssc;
  wire FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_and_32_tmp;
  wire FpAdd_8U_23U_is_inf_1_lpi_1_dfm;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w0;
  wire alu_nan_to_zero_op_sign_lpi_1_dfm_mx0w0;
  wire alu_nan_to_zero_op_sign_15_lpi_1_dfm_mx0w0;
  wire alu_nan_to_zero_op_sign_14_lpi_1_dfm_mx0w0;
  wire alu_nan_to_zero_op_sign_13_lpi_1_dfm_mx0w0;
  wire alu_nan_to_zero_op_sign_12_lpi_1_dfm_mx0w0;
  wire alu_nan_to_zero_op_sign_11_lpi_1_dfm_mx0w0;
  wire alu_nan_to_zero_op_sign_10_lpi_1_dfm_mx0w0;
  wire alu_nan_to_zero_op_sign_9_lpi_1_dfm_mx0w0;
  wire alu_nan_to_zero_op_sign_8_lpi_1_dfm_mx0w0;
  wire alu_nan_to_zero_op_sign_7_lpi_1_dfm_mx0w0;
  wire alu_nan_to_zero_op_sign_6_lpi_1_dfm_mx0w0;
  wire alu_nan_to_zero_op_sign_5_lpi_1_dfm_mx0w0;
  wire alu_nan_to_zero_op_sign_4_lpi_1_dfm_mx0w0;
  wire alu_nan_to_zero_op_sign_3_lpi_1_dfm_mx0w0;
  wire alu_nan_to_zero_op_sign_2_lpi_1_dfm_mx0w0;
  wire alu_nan_to_zero_op_sign_1_lpi_1_dfm_mx0w0;
  wire FpCmp_8U_23U_true_else_3_and_45_tmp;
  wire FpAlu_8U_23U_and_276_m1c;
  wire FpAlu_8U_23U_and_277_cse;
  wire FpAlu_8U_23U_and_279_cse;
  wire FpCmp_8U_23U_false_else_3_or_45_tmp;
  wire FpAlu_8U_23U_and_278_m1c;
  wire FpAlu_8U_23U_equal_tmp_2_mx0w0;
  wire FpAlu_8U_23U_equal_tmp_mx0w0;
  wire FpCmp_8U_23U_false_is_a_greater_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_is_a_greater_lpi_1_dfm_2_mx0;
  wire FpAlu_8U_23U_nor_dfs_mx0w0;
  wire FpCmp_8U_23U_true_else_3_and_42_tmp;
  wire FpAlu_8U_23U_and_262_m1c;
  wire FpAlu_8U_23U_and_263_cse;
  wire FpAlu_8U_23U_and_265_cse;
  wire FpCmp_8U_23U_false_else_3_or_42_tmp;
  wire FpAlu_8U_23U_and_264_m1c;
  wire FpCmp_8U_23U_false_is_a_greater_15_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_is_a_greater_15_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_else_3_and_39_tmp;
  wire FpAlu_8U_23U_and_248_m1c;
  wire FpAlu_8U_23U_and_249_cse;
  wire FpAlu_8U_23U_and_251_cse;
  wire FpCmp_8U_23U_false_else_3_or_39_tmp;
  wire FpAlu_8U_23U_and_250_m1c;
  wire FpCmp_8U_23U_false_is_a_greater_14_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_is_a_greater_14_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_else_3_and_36_tmp;
  wire FpAlu_8U_23U_and_234_m1c;
  wire FpAlu_8U_23U_and_235_cse;
  wire FpAlu_8U_23U_and_237_cse;
  wire FpCmp_8U_23U_false_else_3_or_36_tmp;
  wire FpAlu_8U_23U_and_236_m1c;
  wire FpCmp_8U_23U_false_is_a_greater_13_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_is_a_greater_13_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_else_3_and_33_tmp;
  wire FpAlu_8U_23U_and_220_m1c;
  wire FpAlu_8U_23U_and_221_cse;
  wire FpAlu_8U_23U_and_223_cse;
  wire FpCmp_8U_23U_false_else_3_or_33_tmp;
  wire FpAlu_8U_23U_and_222_m1c;
  wire FpCmp_8U_23U_false_is_a_greater_12_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_is_a_greater_12_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_else_3_and_30_tmp;
  wire FpAlu_8U_23U_and_206_m1c;
  wire FpAlu_8U_23U_and_207_cse;
  wire FpAlu_8U_23U_and_209_cse;
  wire FpCmp_8U_23U_false_else_3_or_30_tmp;
  wire FpAlu_8U_23U_and_208_m1c;
  wire FpCmp_8U_23U_false_is_a_greater_11_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_is_a_greater_11_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_else_3_and_27_tmp;
  wire FpAlu_8U_23U_and_192_m1c;
  wire FpAlu_8U_23U_and_193_cse;
  wire FpAlu_8U_23U_and_195_cse;
  wire FpCmp_8U_23U_false_else_3_or_27_tmp;
  wire FpAlu_8U_23U_and_194_m1c;
  wire FpCmp_8U_23U_false_is_a_greater_10_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_is_a_greater_10_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_else_3_and_24_tmp;
  wire FpAlu_8U_23U_and_178_m1c;
  wire FpAlu_8U_23U_and_179_cse;
  wire FpAlu_8U_23U_and_181_cse;
  wire FpCmp_8U_23U_false_else_3_or_24_tmp;
  wire FpAlu_8U_23U_and_180_m1c;
  wire FpCmp_8U_23U_false_is_a_greater_9_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_is_a_greater_9_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_else_3_and_21_tmp;
  wire FpAlu_8U_23U_and_164_m1c;
  wire FpAlu_8U_23U_and_165_cse;
  wire FpAlu_8U_23U_and_167_cse;
  wire FpCmp_8U_23U_false_else_3_or_21_tmp;
  wire FpAlu_8U_23U_and_166_m1c;
  wire FpCmp_8U_23U_false_is_a_greater_8_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_is_a_greater_8_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_else_3_and_18_tmp;
  wire FpAlu_8U_23U_and_150_m1c;
  wire FpAlu_8U_23U_and_151_cse;
  wire FpAlu_8U_23U_and_153_cse;
  wire FpCmp_8U_23U_false_else_3_or_18_tmp;
  wire FpAlu_8U_23U_and_152_m1c;
  wire FpCmp_8U_23U_false_is_a_greater_7_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_is_a_greater_7_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_else_3_and_15_tmp;
  wire FpAlu_8U_23U_and_136_m1c;
  wire FpAlu_8U_23U_and_137_cse;
  wire FpAlu_8U_23U_and_139_cse;
  wire FpCmp_8U_23U_false_else_3_or_15_tmp;
  wire FpAlu_8U_23U_and_138_m1c;
  wire FpCmp_8U_23U_false_is_a_greater_6_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_is_a_greater_6_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_else_3_and_12_tmp;
  wire FpAlu_8U_23U_and_122_m1c;
  wire FpAlu_8U_23U_and_123_cse;
  wire FpAlu_8U_23U_and_125_cse;
  wire FpCmp_8U_23U_false_else_3_or_12_tmp;
  wire FpAlu_8U_23U_and_124_m1c;
  wire FpCmp_8U_23U_false_is_a_greater_5_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_is_a_greater_5_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_else_3_and_9_tmp;
  wire FpAlu_8U_23U_and_108_m1c;
  wire FpAlu_8U_23U_and_109_cse;
  wire FpAlu_8U_23U_and_111_cse;
  wire FpCmp_8U_23U_false_else_3_or_9_tmp;
  wire FpAlu_8U_23U_and_110_m1c;
  wire FpCmp_8U_23U_false_is_a_greater_4_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_is_a_greater_4_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_else_3_and_6_tmp;
  wire FpAlu_8U_23U_and_94_m1c;
  wire FpAlu_8U_23U_and_95_cse;
  wire FpAlu_8U_23U_and_97_cse;
  wire FpCmp_8U_23U_false_else_3_or_6_tmp;
  wire FpAlu_8U_23U_and_96_m1c;
  wire FpCmp_8U_23U_false_is_a_greater_3_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_is_a_greater_3_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_else_3_and_3_tmp;
  wire FpAlu_8U_23U_and_80_m1c;
  wire FpAlu_8U_23U_and_81_cse;
  wire FpAlu_8U_23U_and_83_cse;
  wire FpCmp_8U_23U_false_else_3_or_3_tmp;
  wire FpAlu_8U_23U_and_82_m1c;
  wire FpCmp_8U_23U_false_is_a_greater_2_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_is_a_greater_2_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_else_3_and_tmp;
  wire FpAlu_8U_23U_and_66_m1c;
  wire FpAlu_8U_23U_and_67_cse;
  wire FpAlu_8U_23U_and_69_cse;
  wire FpCmp_8U_23U_false_else_3_or_tmp;
  wire FpAlu_8U_23U_and_68_m1c;
  wire FpCmp_8U_23U_false_is_a_greater_1_lpi_1_dfm_2_mx0;
  wire FpCmp_8U_23U_true_is_a_greater_1_lpi_1_dfm_2_mx0;
  wire else_AluOp_data_15_15_lpi_1_dfm_mx0;
  wire else_AluOp_data_14_15_lpi_1_dfm_mx0;
  wire else_AluOp_data_13_15_lpi_1_dfm_mx0;
  wire else_AluOp_data_12_15_lpi_1_dfm_mx0;
  wire else_AluOp_data_11_15_lpi_1_dfm_mx0;
  wire else_AluOp_data_10_15_lpi_1_dfm_mx0;
  wire else_AluOp_data_9_15_lpi_1_dfm_mx0;
  wire else_AluOp_data_8_15_lpi_1_dfm_mx0;
  wire else_AluOp_data_7_15_lpi_1_dfm_mx0;
  wire else_AluOp_data_6_15_lpi_1_dfm_mx0;
  wire else_AluOp_data_5_15_lpi_1_dfm_mx0;
  wire else_AluOp_data_4_15_lpi_1_dfm_mx0;
  wire else_AluOp_data_3_15_lpi_1_dfm_mx0;
  wire else_AluOp_data_2_15_lpi_1_dfm_mx0;
  wire else_AluOp_data_1_15_lpi_1_dfm_mx0;
  wire else_AluOp_data_0_15_lpi_1_dfm_mx0;
  wire [9:0] else_AluOp_data_15_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_AluOp_data_14_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_AluOp_data_13_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_AluOp_data_12_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_AluOp_data_11_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_AluOp_data_10_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_AluOp_data_9_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_AluOp_data_8_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_AluOp_data_7_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_AluOp_data_6_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_AluOp_data_5_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_AluOp_data_4_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_AluOp_data_3_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_AluOp_data_2_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_AluOp_data_1_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_AluOp_data_0_9_0_lpi_1_dfm_mx0;
  wire [3:0] FpAdd_8U_23U_o_expo_lpi_1_dfm_2_7_4;
  wire [3:0] FpAdd_8U_23U_o_expo_15_lpi_1_dfm_2_7_4;
  wire [3:0] FpAdd_8U_23U_o_expo_14_lpi_1_dfm_2_7_4;
  wire [3:0] FpAdd_8U_23U_o_expo_13_lpi_1_dfm_2_7_4;
  wire [3:0] FpAdd_8U_23U_o_expo_12_lpi_1_dfm_2_7_4;
  wire [3:0] FpAdd_8U_23U_o_expo_11_lpi_1_dfm_2_7_4;
  wire [3:0] FpAdd_8U_23U_o_expo_10_lpi_1_dfm_2_7_4;
  wire [3:0] FpAdd_8U_23U_o_expo_9_lpi_1_dfm_2_7_4;
  wire [3:0] FpAdd_8U_23U_o_expo_8_lpi_1_dfm_2_7_4;
  wire [3:0] FpAdd_8U_23U_o_expo_7_lpi_1_dfm_2_7_4;
  wire [3:0] FpAdd_8U_23U_o_expo_6_lpi_1_dfm_2_7_4;
  wire [3:0] FpAdd_8U_23U_o_expo_5_lpi_1_dfm_2_7_4;
  wire [3:0] FpAdd_8U_23U_o_expo_4_lpi_1_dfm_2_7_4;
  wire [3:0] FpAdd_8U_23U_o_expo_3_lpi_1_dfm_2_7_4;
  wire [3:0] FpAdd_8U_23U_o_expo_2_lpi_1_dfm_2_7_4;
  wire [3:0] FpAdd_8U_23U_o_expo_1_lpi_1_dfm_2_7_4;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_15_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_15_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_14_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_14_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_13_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_13_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_12_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_12_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_11_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_11_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_10_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_10_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_9_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_9_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_8_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_8_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_7_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_7_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_6_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_6_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_5_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_5_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_4_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_4_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_3_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_3_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_2_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_2_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_1_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_1_lpi_1_dfm;
  wire alu_nan_to_zero_land_lpi_1_dfm;
  wire alu_nan_to_zero_land_15_lpi_1_dfm;
  wire alu_nan_to_zero_land_14_lpi_1_dfm;
  wire alu_nan_to_zero_land_13_lpi_1_dfm;
  wire alu_nan_to_zero_land_12_lpi_1_dfm;
  wire alu_nan_to_zero_land_11_lpi_1_dfm;
  wire alu_nan_to_zero_land_10_lpi_1_dfm;
  wire alu_nan_to_zero_land_9_lpi_1_dfm;
  wire alu_nan_to_zero_land_8_lpi_1_dfm;
  wire alu_nan_to_zero_land_7_lpi_1_dfm;
  wire alu_nan_to_zero_land_6_lpi_1_dfm;
  wire alu_nan_to_zero_land_5_lpi_1_dfm;
  wire alu_nan_to_zero_land_4_lpi_1_dfm;
  wire alu_nan_to_zero_land_3_lpi_1_dfm;
  wire alu_nan_to_zero_land_2_lpi_1_dfm;
  wire alu_nan_to_zero_land_1_lpi_1_dfm;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_mx2;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_mx2;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_mx2;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_mx2;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_mx2;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_mx2;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_mx2;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_mx2;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_mx2;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_mx2;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_mx2;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_mx2;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_mx2;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_mx2;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_mx2;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_mx2;
  wire [3:0] FpAdd_8U_23U_o_expo_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_8U_23U_o_expo_15_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_8U_23U_o_expo_14_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_8U_23U_o_expo_13_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_8U_23U_o_expo_12_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_8U_23U_o_expo_11_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_8U_23U_o_expo_10_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_8U_23U_o_expo_9_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_8U_23U_o_expo_8_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_8U_23U_o_expo_7_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_8U_23U_o_expo_6_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_8U_23U_o_expo_5_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_8U_23U_o_expo_4_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_8U_23U_o_expo_3_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_8U_23U_o_expo_2_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_8U_23U_o_expo_1_lpi_1_dfm_2_3_0;
  wire [9:0] alu_nan_to_zero_op_mant_lpi_1_dfm;
  wire [9:0] alu_nan_to_zero_op_mant_15_lpi_1_dfm;
  wire [9:0] alu_nan_to_zero_op_mant_14_lpi_1_dfm;
  wire [9:0] alu_nan_to_zero_op_mant_13_lpi_1_dfm;
  wire [9:0] alu_nan_to_zero_op_mant_12_lpi_1_dfm;
  wire [9:0] alu_nan_to_zero_op_mant_11_lpi_1_dfm;
  wire [9:0] alu_nan_to_zero_op_mant_10_lpi_1_dfm;
  wire [9:0] alu_nan_to_zero_op_mant_9_lpi_1_dfm;
  wire [9:0] alu_nan_to_zero_op_mant_8_lpi_1_dfm;
  wire [9:0] alu_nan_to_zero_op_mant_7_lpi_1_dfm;
  wire [9:0] alu_nan_to_zero_op_mant_6_lpi_1_dfm;
  wire [9:0] alu_nan_to_zero_op_mant_5_lpi_1_dfm;
  wire [9:0] alu_nan_to_zero_op_mant_4_lpi_1_dfm;
  wire [9:0] alu_nan_to_zero_op_mant_3_lpi_1_dfm;
  wire [9:0] alu_nan_to_zero_op_mant_2_lpi_1_dfm;
  wire [9:0] alu_nan_to_zero_op_mant_1_lpi_1_dfm;
  wire [4:0] alu_nan_to_zero_op_expo_lpi_1_dfm;
  wire [4:0] alu_nan_to_zero_op_expo_15_lpi_1_dfm;
  wire [4:0] alu_nan_to_zero_op_expo_14_lpi_1_dfm;
  wire [4:0] alu_nan_to_zero_op_expo_13_lpi_1_dfm;
  wire [4:0] alu_nan_to_zero_op_expo_12_lpi_1_dfm;
  wire [4:0] alu_nan_to_zero_op_expo_11_lpi_1_dfm;
  wire [4:0] alu_nan_to_zero_op_expo_10_lpi_1_dfm;
  wire [4:0] alu_nan_to_zero_op_expo_9_lpi_1_dfm;
  wire [4:0] alu_nan_to_zero_op_expo_8_lpi_1_dfm;
  wire [4:0] alu_nan_to_zero_op_expo_7_lpi_1_dfm;
  wire [4:0] alu_nan_to_zero_op_expo_6_lpi_1_dfm;
  wire [4:0] alu_nan_to_zero_op_expo_5_lpi_1_dfm;
  wire [4:0] alu_nan_to_zero_op_expo_4_lpi_1_dfm;
  wire [4:0] alu_nan_to_zero_op_expo_3_lpi_1_dfm;
  wire [4:0] alu_nan_to_zero_op_expo_2_lpi_1_dfm;
  wire [4:0] alu_nan_to_zero_op_expo_1_lpi_1_dfm;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_22_13_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_22_13_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_22_13_mx2;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_12_10_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_9_0_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_9_0_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_9_0_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_22_13_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_22_13_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_22_13_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_22_13_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_22_13_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_22_13_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_22_13_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_22_13_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_22_13_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_22_13_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_22_13_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_22_13_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_22_13_mx2;
  wire [78:0] IntShiftLeft_16U_6U_32U_mbits_fixed_sva;
  wire [78:0] IntShiftLeft_16U_6U_32U_mbits_fixed_15_sva;
  wire [78:0] IntShiftLeft_16U_6U_32U_mbits_fixed_14_sva;
  wire [78:0] IntShiftLeft_16U_6U_32U_mbits_fixed_13_sva;
  wire [78:0] IntShiftLeft_16U_6U_32U_mbits_fixed_12_sva;
  wire [78:0] IntShiftLeft_16U_6U_32U_mbits_fixed_11_sva;
  wire [78:0] IntShiftLeft_16U_6U_32U_mbits_fixed_10_sva;
  wire [78:0] IntShiftLeft_16U_6U_32U_mbits_fixed_9_sva;
  wire [78:0] IntShiftLeft_16U_6U_32U_mbits_fixed_8_sva;
  wire [78:0] IntShiftLeft_16U_6U_32U_mbits_fixed_7_sva;
  wire [78:0] IntShiftLeft_16U_6U_32U_mbits_fixed_6_sva;
  wire [78:0] IntShiftLeft_16U_6U_32U_mbits_fixed_5_sva;
  wire [78:0] IntShiftLeft_16U_6U_32U_mbits_fixed_4_sva;
  wire [78:0] IntShiftLeft_16U_6U_32U_mbits_fixed_3_sva;
  wire [78:0] IntShiftLeft_16U_6U_32U_mbits_fixed_2_sva;
  wire [78:0] IntShiftLeft_16U_6U_32U_mbits_fixed_1_sva;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_12_10_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_9_0_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_9_0_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_9_0_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_9_0_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_9_0_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_9_0_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_9_0_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_9_0_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_9_0_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_9_0_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_9_0_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_9_0_mx2;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_9_0_mx2;
  wire or_4809_cse;
  wire chn_alu_out_and_cse;
  reg reg_cfg_alu_shift_value_rsc_triosy_obj_ld_core_psct_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_cse;
  wire nor_1748_cse;
  wire nor_1720_cse;
  wire nor_1724_cse;
  wire nor_333_cse;
  wire or_899_cse;
  wire nor_1693_cse;
  wire nor_1697_cse;
  wire nor_1666_cse;
  wire nor_1670_cse;
  wire nor_1639_cse;
  wire nor_1643_cse;
  wire nor_1612_cse;
  wire nor_1616_cse;
  wire nor_1585_cse;
  wire nor_1589_cse;
  wire nor_1559_cse;
  wire nor_1563_cse;
  wire nor_1533_cse;
  wire nor_1537_cse;
  wire nor_1507_cse;
  wire nor_1511_cse;
  wire nor_1481_cse;
  wire nor_1485_cse;
  wire nor_1455_cse;
  wire nor_1459_cse;
  wire nor_1429_cse;
  wire nor_1433_cse;
  wire nor_1403_cse;
  wire nor_1407_cse;
  wire nor_1378_cse;
  wire nor_1353_cse;
  reg reg_chn_alu_out_rsci_ld_core_psct_cse;
  wire IsNaN_8U_23U_2_aelse_and_cse;
  wire AluIn_data_and_cse;
  wire FpAdd_8U_23U_int_mant_p1_and_cse;
  wire alu_loop_op_else_if_and_cse;
  wire alu_loop_op_else_else_if_and_cse;
  wire FpAdd_8U_23U_b_left_shift_and_cse;
  wire nor_1317_cse;
  wire or_1935_cse;
  wire and_3689_cse;
  wire nor_1813_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_14_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_15_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_17_cse;
  reg reg_alu_loop_op_2_FpAdd_8U_23U_is_a_greater_slc_8_1_svs_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_20_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_23_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_26_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_29_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_32_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_35_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_38_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_41_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_44_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_47_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_50_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_53_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_56_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_59_cse;
  wire and_3707_cse;
  wire FpAdd_8U_23U_and_144_cse;
  wire FpAdd_8U_23U_and_146_cse;
  wire FpAdd_8U_23U_and_148_cse;
  wire FpAdd_8U_23U_and_150_cse;
  wire FpAdd_8U_23U_and_152_cse;
  wire FpAdd_8U_23U_and_154_cse;
  wire FpAdd_8U_23U_and_156_cse;
  wire FpAdd_8U_23U_and_158_cse;
  wire FpAdd_8U_23U_and_160_cse;
  wire FpAdd_8U_23U_and_162_cse;
  wire FpAdd_8U_23U_and_164_cse;
  wire FpAdd_8U_23U_and_166_cse;
  wire FpAdd_8U_23U_and_168_cse;
  wire FpAdd_8U_23U_and_170_cse;
  wire FpAdd_8U_23U_and_172_cse;
  wire FpAdd_8U_23U_and_174_cse;
  wire FpAlu_8U_23U_and_692_cse;
  wire alu_loop_op_else_if_and_9_cse;
  wire alu_loop_op_else_else_if_and_9_cse;
  wire alu_loop_op_else_if_and_12_cse;
  wire alu_loop_op_else_else_if_and_12_cse;
  wire alu_loop_op_else_if_and_15_cse;
  wire alu_loop_op_else_else_if_and_15_cse;
  wire alu_loop_op_else_if_and_18_cse;
  wire alu_loop_op_else_else_if_and_18_cse;
  wire alu_loop_op_else_if_and_21_cse;
  wire alu_loop_op_else_else_if_and_21_cse;
  wire alu_loop_op_else_if_and_24_cse;
  wire alu_loop_op_else_else_if_and_24_cse;
  wire alu_loop_op_else_if_and_27_cse;
  wire alu_loop_op_else_else_if_and_27_cse;
  wire alu_loop_op_else_if_and_30_cse;
  wire alu_loop_op_else_else_if_and_30_cse;
  wire alu_loop_op_else_if_and_33_cse;
  wire alu_loop_op_else_else_if_and_33_cse;
  wire alu_loop_op_else_if_and_36_cse;
  wire alu_loop_op_else_else_if_and_36_cse;
  wire alu_loop_op_else_if_and_39_cse;
  wire alu_loop_op_else_else_if_and_39_cse;
  wire alu_loop_op_else_if_and_42_cse;
  wire alu_loop_op_else_else_if_and_42_cse;
  wire alu_loop_op_else_if_and_45_cse;
  wire alu_loop_op_else_else_if_and_45_cse;
  wire alu_loop_op_else_if_and_48_cse;
  wire alu_loop_op_else_else_if_and_48_cse;
  wire alu_loop_op_else_if_and_51_cse;
  wire alu_loop_op_else_else_if_and_51_cse;
  wire alu_loop_op_else_if_and_54_cse;
  wire alu_loop_op_else_else_if_and_54_cse;
  wire alu_nan_to_zero_op_sign_and_cse;
  wire FpAdd_8U_23U_is_a_greater_and_cse;
  wire IsZero_8U_23U_and_cse;
  wire FpAdd_8U_23U_is_a_greater_and_1_cse;
  wire FpAdd_8U_23U_is_a_greater_and_3_cse;
  wire FpAdd_8U_23U_is_a_greater_and_8_cse;
  wire IntShiftLeft_16U_6U_32U_and_cse;
  wire IsZero_8U_23U_and_16_cse;
  wire alu_loop_op_if_alu_loop_op_if_nor_cse;
  wire alu_loop_op_if_alu_loop_op_if_nor_1_cse;
  wire alu_loop_op_if_alu_loop_op_if_nor_2_cse;
  wire alu_loop_op_if_alu_loop_op_if_nor_3_cse;
  wire alu_loop_op_if_alu_loop_op_if_nor_4_cse;
  wire alu_loop_op_if_alu_loop_op_if_nor_5_cse;
  wire alu_loop_op_if_alu_loop_op_if_nor_6_cse;
  wire alu_loop_op_if_alu_loop_op_if_nor_7_cse;
  wire alu_loop_op_if_alu_loop_op_if_nor_8_cse;
  wire alu_loop_op_if_alu_loop_op_if_nor_9_cse;
  wire alu_loop_op_if_alu_loop_op_if_nor_10_cse;
  wire alu_loop_op_if_alu_loop_op_if_nor_11_cse;
  wire alu_loop_op_if_alu_loop_op_if_nor_12_cse;
  wire alu_loop_op_if_alu_loop_op_if_nor_13_cse;
  wire alu_loop_op_if_alu_loop_op_if_nor_14_cse;
  wire alu_loop_op_if_alu_loop_op_if_nor_15_cse;
  wire or_22_cse;
  wire nor_2061_cse;
  wire or_334_cse;
  wire or_350_cse;
  wire or_1923_cse;
  wire or_3303_cse;
  wire and_dcpl_1789;
  wire or_dcpl_1047;
  wire and_dcpl_1796;
  wire or_dcpl_1052;
  wire and_dcpl_1804;
  wire or_dcpl_1057;
  wire and_dcpl_1812;
  wire or_dcpl_1062;
  wire and_dcpl_1820;
  wire or_dcpl_1067;
  wire and_dcpl_1828;
  wire or_dcpl_1072;
  wire and_dcpl_1836;
  wire or_dcpl_1077;
  wire and_dcpl_1844;
  wire or_dcpl_1082;
  wire and_dcpl_1852;
  wire or_dcpl_1087;
  wire and_dcpl_1860;
  wire or_dcpl_1092;
  wire and_dcpl_1868;
  wire or_dcpl_1097;
  wire and_dcpl_1876;
  wire or_dcpl_1102;
  wire and_dcpl_1884;
  wire or_dcpl_1107;
  wire and_dcpl_1892;
  wire or_dcpl_1112;
  wire and_dcpl_1900;
  wire or_dcpl_1117;
  wire and_dcpl_1908;
  wire or_dcpl_1122;
  wire and_dcpl_1916;
  wire FpAdd_8U_23U_and_ssc;
  wire FpAdd_8U_23U_and_2_ssc;
  wire FpAdd_8U_23U_and_4_ssc;
  wire FpAdd_8U_23U_and_6_ssc;
  wire FpAdd_8U_23U_and_8_ssc;
  wire FpAdd_8U_23U_and_10_ssc;
  wire FpAdd_8U_23U_and_12_ssc;
  wire FpAdd_8U_23U_and_14_ssc;
  wire FpAdd_8U_23U_and_16_ssc;
  wire FpAdd_8U_23U_and_18_ssc;
  wire FpAdd_8U_23U_and_20_ssc;
  wire FpAdd_8U_23U_and_22_ssc;
  wire FpAdd_8U_23U_and_24_ssc;
  wire FpAdd_8U_23U_and_26_ssc;
  wire FpAdd_8U_23U_and_28_ssc;
  wire FpAdd_8U_23U_and_30_ssc;
  wire [7:0] FpAdd_8U_23U_o_expo_1_sva_4;
  wire [8:0] nl_FpAdd_8U_23U_o_expo_1_sva_4;
  wire FpAdd_8U_23U_and_51_ssc;
  wire nor_7_ssc;
  wire [7:0] FpAdd_8U_23U_o_expo_2_sva_4;
  wire [8:0] nl_FpAdd_8U_23U_o_expo_2_sva_4;
  wire FpAdd_8U_23U_and_55_ssc;
  wire [7:0] FpAdd_8U_23U_o_expo_3_sva_4;
  wire [8:0] nl_FpAdd_8U_23U_o_expo_3_sva_4;
  wire FpAdd_8U_23U_and_59_ssc;
  wire [7:0] FpAdd_8U_23U_o_expo_4_sva_4;
  wire [8:0] nl_FpAdd_8U_23U_o_expo_4_sva_4;
  wire FpAdd_8U_23U_and_63_ssc;
  wire [7:0] FpAdd_8U_23U_o_expo_5_sva_4;
  wire [8:0] nl_FpAdd_8U_23U_o_expo_5_sva_4;
  wire FpAdd_8U_23U_and_67_ssc;
  wire [7:0] FpAdd_8U_23U_o_expo_6_sva_4;
  wire [8:0] nl_FpAdd_8U_23U_o_expo_6_sva_4;
  wire FpAdd_8U_23U_and_71_ssc;
  wire [7:0] FpAdd_8U_23U_o_expo_7_sva_4;
  wire [8:0] nl_FpAdd_8U_23U_o_expo_7_sva_4;
  wire FpAdd_8U_23U_and_75_ssc;
  wire [7:0] FpAdd_8U_23U_o_expo_8_sva_4;
  wire [8:0] nl_FpAdd_8U_23U_o_expo_8_sva_4;
  wire FpAdd_8U_23U_and_79_ssc;
  wire [7:0] FpAdd_8U_23U_o_expo_9_sva_4;
  wire [8:0] nl_FpAdd_8U_23U_o_expo_9_sva_4;
  wire FpAdd_8U_23U_and_83_ssc;
  wire [7:0] FpAdd_8U_23U_o_expo_10_sva_4;
  wire [8:0] nl_FpAdd_8U_23U_o_expo_10_sva_4;
  wire FpAdd_8U_23U_and_87_ssc;
  wire [7:0] FpAdd_8U_23U_o_expo_11_sva_4;
  wire [8:0] nl_FpAdd_8U_23U_o_expo_11_sva_4;
  wire FpAdd_8U_23U_and_91_ssc;
  wire [7:0] FpAdd_8U_23U_o_expo_12_sva_4;
  wire [8:0] nl_FpAdd_8U_23U_o_expo_12_sva_4;
  wire FpAdd_8U_23U_and_95_ssc;
  wire [7:0] FpAdd_8U_23U_o_expo_13_sva_4;
  wire [8:0] nl_FpAdd_8U_23U_o_expo_13_sva_4;
  wire FpAdd_8U_23U_and_99_ssc;
  wire [7:0] FpAdd_8U_23U_o_expo_14_sva_4;
  wire [8:0] nl_FpAdd_8U_23U_o_expo_14_sva_4;
  wire FpAdd_8U_23U_and_103_ssc;
  wire [7:0] FpAdd_8U_23U_o_expo_15_sva_4;
  wire [8:0] nl_FpAdd_8U_23U_o_expo_15_sva_4;
  wire FpAdd_8U_23U_and_107_ssc;
  wire [7:0] FpAdd_8U_23U_o_expo_sva_4;
  wire [8:0] nl_FpAdd_8U_23U_o_expo_sva_4;
  wire FpAdd_8U_23U_and_111_ssc;
  wire asn_1837;
  wire or_cse_2;
  wire and_498_rgt;
  wire and_543_rgt;
  wire and_589_rgt;
  wire and_715_rgt;
  wire and_719_rgt;
  wire and_723_rgt;
  wire and_726_rgt;
  wire and_730_rgt;
  wire and_733_rgt;
  wire and_737_rgt;
  wire and_741_rgt;
  wire and_745_rgt;
  wire and_749_rgt;
  wire and_753_rgt;
  wire and_757_rgt;
  wire and_761_rgt;
  wire and_764_rgt;
  wire and_768_rgt;
  wire and_772_rgt;
  wire and_776_rgt;
  wire and_779_rgt;
  wire and_783_rgt;
  wire and_786_rgt;
  wire and_790_rgt;
  wire and_794_rgt;
  wire and_798_rgt;
  wire and_802_rgt;
  wire and_806_rgt;
  wire and_810_rgt;
  wire and_814_rgt;
  wire and_817_rgt;
  wire and_821_rgt;
  wire and_824_rgt;
  wire and_828_rgt;
  wire and_831_rgt;
  wire and_1106_rgt;
  wire and_1108_rgt;
  wire and_1135_rgt;
  wire and_1308_rgt;
  wire and_1311_rgt;
  wire and_1313_rgt;
  wire and_1315_rgt;
  wire and_1316_rgt;
  wire and_1323_rgt;
  wire and_1325_rgt;
  wire and_1327_rgt;
  wire and_1328_rgt;
  wire and_1333_rgt;
  wire and_1335_rgt;
  wire and_1337_rgt;
  wire and_1339_rgt;
  wire and_1346_rgt;
  wire and_1347_rgt;
  wire and_1351_rgt;
  wire and_1353_rgt;
  wire and_1355_rgt;
  wire and_1356_rgt;
  wire and_1364_rgt;
  wire and_1366_rgt;
  wire and_1368_rgt;
  wire and_1369_rgt;
  wire and_1380_rgt;
  wire and_1382_rgt;
  wire and_1384_rgt;
  wire and_1386_rgt;
  wire and_1391_rgt;
  wire and_1393_rgt;
  wire and_1395_rgt;
  wire and_1396_rgt;
  wire and_1400_rgt;
  wire and_1402_rgt;
  wire and_1404_rgt;
  wire and_1406_rgt;
  wire and_1413_rgt;
  wire and_1415_rgt;
  wire and_1417_rgt;
  wire and_1418_rgt;
  wire and_1425_rgt;
  wire and_1427_rgt;
  wire and_1429_rgt;
  wire and_1431_rgt;
  wire and_1438_rgt;
  wire and_1440_rgt;
  wire and_1442_rgt;
  wire and_1444_rgt;
  wire and_1452_rgt;
  wire and_1454_rgt;
  wire and_1456_rgt;
  wire and_1458_rgt;
  wire and_1469_rgt;
  wire and_1471_rgt;
  wire and_1473_rgt;
  wire and_1475_rgt;
  wire and_1481_rgt;
  wire and_1483_rgt;
  wire and_1485_rgt;
  wire and_1487_rgt;
  wire and_1492_rgt;
  wire and_1494_rgt;
  wire and_1496_rgt;
  wire and_1498_rgt;
  wire and_1503_rgt;
  wire and_1505_rgt;
  wire and_1507_rgt;
  wire and_1508_rgt;
  wire and_1895_rgt;
  wire and_1899_rgt;
  wire and_1903_rgt;
  wire and_1907_rgt;
  wire and_1911_rgt;
  wire and_1921_rgt;
  wire and_1925_rgt;
  wire and_1929_rgt;
  wire and_1933_rgt;
  wire and_2163_rgt;
  wire and_2167_rgt;
  wire and_2171_rgt;
  wire and_2175_rgt;
  wire and_2179_rgt;
  wire and_2183_rgt;
  wire and_2185_rgt;
  wire and_2186_rgt;
  wire and_2193_rgt;
  wire and_2198_rgt;
  wire [48:0] alu_loop_op_1_FpNormalize_8U_49U_else_lshift_itm;
  wire [48:0] alu_loop_op_2_FpNormalize_8U_49U_else_lshift_1_itm;
  wire [48:0] alu_loop_op_3_FpNormalize_8U_49U_else_lshift_itm;
  wire [48:0] alu_loop_op_4_FpNormalize_8U_49U_else_lshift_1_itm;
  wire [48:0] alu_loop_op_5_FpNormalize_8U_49U_else_lshift_itm;
  wire [48:0] alu_loop_op_6_FpNormalize_8U_49U_else_lshift_1_itm;
  wire [48:0] alu_loop_op_7_FpNormalize_8U_49U_else_lshift_itm;
  wire [48:0] alu_loop_op_8_FpNormalize_8U_49U_else_lshift_1_itm;
  wire [48:0] alu_loop_op_9_FpNormalize_8U_49U_else_lshift_itm;
  wire [48:0] alu_loop_op_10_FpNormalize_8U_49U_else_lshift_1_itm;
  wire [48:0] alu_loop_op_11_FpNormalize_8U_49U_else_lshift_itm;
  wire [48:0] alu_loop_op_12_FpNormalize_8U_49U_else_lshift_1_itm;
  wire [48:0] alu_loop_op_13_FpNormalize_8U_49U_else_lshift_itm;
  wire [48:0] alu_loop_op_14_FpNormalize_8U_49U_else_lshift_1_itm;
  wire [48:0] alu_loop_op_15_FpNormalize_8U_49U_else_lshift_itm;
  wire [48:0] alu_loop_op_16_FpNormalize_8U_49U_else_lshift_1_itm;
  wire mux_16_itm;
  wire mux_127_itm;
  wire mux_393_itm;
  wire mux_415_itm;
  wire mux_478_itm;
  wire mux_604_itm;
  wire mux_782_itm;
  wire mux_1425_itm;
  wire FpNormalize_8U_49U_else_and_tmp;
  wire [7:0] z_out;
  wire FpNormalize_8U_49U_else_and_tmp_1;
  wire [7:0] z_out_1;
  wire FpNormalize_8U_49U_else_and_tmp_2;
  wire [7:0] z_out_2;
  wire FpNormalize_8U_49U_else_and_tmp_3;
  wire [7:0] z_out_3;
  wire FpNormalize_8U_49U_else_and_tmp_4;
  wire [7:0] z_out_4;
  wire FpNormalize_8U_49U_else_and_tmp_5;
  wire [7:0] z_out_5;
  wire FpNormalize_8U_49U_else_and_tmp_6;
  wire [7:0] z_out_6;
  wire FpNormalize_8U_49U_else_and_tmp_7;
  wire [7:0] z_out_7;
  wire FpNormalize_8U_49U_else_and_tmp_8;
  wire [7:0] z_out_8;
  wire FpNormalize_8U_49U_else_and_tmp_9;
  wire [7:0] z_out_9;
  wire FpNormalize_8U_49U_else_and_tmp_10;
  wire [7:0] z_out_10;
  wire FpNormalize_8U_49U_else_and_tmp_11;
  wire [7:0] z_out_11;
  wire FpNormalize_8U_49U_else_and_tmp_12;
  wire [7:0] z_out_12;
  wire FpNormalize_8U_49U_else_and_tmp_13;
  wire [7:0] z_out_13;
  wire FpNormalize_8U_49U_else_and_tmp_14;
  wire [7:0] z_out_14;
  wire FpNormalize_8U_49U_else_and_tmp_15;
  wire [7:0] z_out_15;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp;
  wire [7:0] z_out_16;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_1;
  wire [7:0] z_out_17;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_2;
  wire [7:0] z_out_18;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_3;
  wire [7:0] z_out_19;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_4;
  wire [7:0] z_out_20;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_5;
  wire [7:0] z_out_21;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_6;
  wire [7:0] z_out_22;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_7;
  wire [7:0] z_out_23;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_8;
  wire [7:0] z_out_24;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_9;
  wire [7:0] z_out_25;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_10;
  wire [7:0] z_out_26;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_11;
  wire [7:0] z_out_27;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_12;
  wire [7:0] z_out_28;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_13;
  wire [7:0] z_out_29;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_14;
  wire [7:0] z_out_30;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_15;
  wire [7:0] z_out_31;
  wire chn_alu_in_rsci_ld_core_psct_mx0c0;
  wire chn_alu_op_rsci_ld_core_psct_mx0c1;
  wire alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
  wire main_stage_v_2_mx0c1;
  wire alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0;
  wire alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0;
  wire alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0;
  wire alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0;
  wire alu_loop_op_5_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0;
  wire alu_loop_op_6_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0;
  wire alu_loop_op_7_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0;
  wire alu_loop_op_8_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0;
  wire alu_loop_op_9_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0;
  wire alu_loop_op_10_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0;
  wire alu_loop_op_11_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0;
  wire alu_loop_op_12_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0;
  wire alu_loop_op_13_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0;
  wire alu_loop_op_14_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0;
  wire alu_loop_op_15_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0;
  wire alu_loop_op_16_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0;
  wire main_stage_v_3_mx0c1;
  wire [7:0] alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
  wire [7:0] alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
  wire [7:0] alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
  wire [7:0] alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
  wire [7:0] alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
  wire [7:0] alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
  wire [7:0] alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
  wire [7:0] alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
  wire [7:0] alu_loop_op_5_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_5_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
  wire [7:0] alu_loop_op_5_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_5_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
  wire [7:0] alu_loop_op_6_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_6_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
  wire [7:0] alu_loop_op_6_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_6_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
  wire [7:0] alu_loop_op_7_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_7_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
  wire [7:0] alu_loop_op_7_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_7_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
  wire [7:0] alu_loop_op_8_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_8_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
  wire [7:0] alu_loop_op_8_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_8_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
  wire [7:0] alu_loop_op_9_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_9_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
  wire [7:0] alu_loop_op_9_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_9_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
  wire [7:0] alu_loop_op_10_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_10_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
  wire [7:0] alu_loop_op_10_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_10_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
  wire [7:0] alu_loop_op_11_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_11_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
  wire [7:0] alu_loop_op_11_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_11_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
  wire [7:0] alu_loop_op_12_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_12_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
  wire [7:0] alu_loop_op_12_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_12_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
  wire [7:0] alu_loop_op_13_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_13_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
  wire [7:0] alu_loop_op_13_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_13_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
  wire [7:0] alu_loop_op_14_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_14_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
  wire [7:0] alu_loop_op_14_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_14_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
  wire [7:0] alu_loop_op_15_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_15_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
  wire [7:0] alu_loop_op_15_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_15_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
  wire [7:0] alu_loop_op_16_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_16_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
  wire [7:0] alu_loop_op_16_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
  wire [8:0] nl_alu_loop_op_16_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
  wire main_stage_v_4_mx0c1;
  wire FpNormalize_8U_49U_if_or_itm_mx0w0;
  wire FpNormalize_8U_49U_if_or_1_itm_mx0w0;
  wire FpNormalize_8U_49U_if_or_2_itm_mx0w0;
  wire FpNormalize_8U_49U_if_or_3_itm_mx0w0;
  wire FpNormalize_8U_49U_if_or_4_itm_mx0w0;
  wire FpNormalize_8U_49U_if_or_5_itm_mx0w0;
  wire FpNormalize_8U_49U_if_or_6_itm_mx0w0;
  wire FpNormalize_8U_49U_if_or_7_itm_mx0w0;
  wire FpNormalize_8U_49U_if_or_8_itm_mx0w0;
  wire FpNormalize_8U_49U_if_or_9_itm_mx0w0;
  wire FpNormalize_8U_49U_if_or_10_itm_mx0w0;
  wire FpNormalize_8U_49U_if_or_11_itm_mx0w0;
  wire FpNormalize_8U_49U_if_or_12_itm_mx0w0;
  wire FpNormalize_8U_49U_if_or_13_itm_mx0w0;
  wire FpNormalize_8U_49U_if_or_14_itm_mx0w0;
  wire FpNormalize_8U_49U_if_or_15_itm_mx0w0;
  wire main_stage_v_1_mx0c1;
  wire cfg_alu_src_1_sva_st_1_mx0c1;
  wire [49:0] FpAdd_8U_23U_asn_76_mx1w1;
  wire [51:0] nl_FpAdd_8U_23U_asn_76_mx1w1;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_mx1;
  wire [49:0] FpAdd_8U_23U_asn_73_mx1w1;
  wire [51:0] nl_FpAdd_8U_23U_asn_73_mx1w1;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_mx1;
  wire [49:0] FpAdd_8U_23U_asn_70_mx1w1;
  wire [51:0] nl_FpAdd_8U_23U_asn_70_mx1w1;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_mx1;
  wire [49:0] FpAdd_8U_23U_asn_67_mx1w1;
  wire [51:0] nl_FpAdd_8U_23U_asn_67_mx1w1;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_mx1;
  wire [49:0] FpAdd_8U_23U_asn_64_mx1w1;
  wire [51:0] nl_FpAdd_8U_23U_asn_64_mx1w1;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_mx1;
  wire [49:0] FpAdd_8U_23U_asn_61_mx1w1;
  wire [51:0] nl_FpAdd_8U_23U_asn_61_mx1w1;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_mx1;
  wire [49:0] FpAdd_8U_23U_asn_58_mx1w1;
  wire [51:0] nl_FpAdd_8U_23U_asn_58_mx1w1;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_mx1;
  wire [49:0] FpAdd_8U_23U_asn_55_mx1w1;
  wire [51:0] nl_FpAdd_8U_23U_asn_55_mx1w1;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_mx1;
  wire [49:0] FpAdd_8U_23U_asn_52_mx1w1;
  wire [51:0] nl_FpAdd_8U_23U_asn_52_mx1w1;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_mx1;
  wire [49:0] FpAdd_8U_23U_asn_49_mx1w1;
  wire [51:0] nl_FpAdd_8U_23U_asn_49_mx1w1;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_mx1;
  wire [49:0] FpAdd_8U_23U_asn_46_mx1w1;
  wire [51:0] nl_FpAdd_8U_23U_asn_46_mx1w1;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_mx1;
  wire [49:0] FpAdd_8U_23U_asn_43_mx1w1;
  wire [51:0] nl_FpAdd_8U_23U_asn_43_mx1w1;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_mx1;
  wire [49:0] FpAdd_8U_23U_asn_40_mx1w1;
  wire [51:0] nl_FpAdd_8U_23U_asn_40_mx1w1;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_mx1;
  wire [49:0] FpAdd_8U_23U_asn_37_mx1w1;
  wire [51:0] nl_FpAdd_8U_23U_asn_37_mx1w1;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_mx1;
  wire [49:0] FpAdd_8U_23U_asn_34_mx1w1;
  wire [51:0] nl_FpAdd_8U_23U_asn_34_mx1w1;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_mx1;
  wire [49:0] FpAdd_8U_23U_asn_mx1w1;
  wire [51:0] nl_FpAdd_8U_23U_asn_mx1w1;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_mx1;
  wire alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
  wire alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
  wire alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
  wire alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
  wire alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0;
  wire alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
  wire alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0;
  wire alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
  wire alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0;
  wire alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0;
  wire alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
  wire alu_loop_op_5_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0;
  wire alu_loop_op_6_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0;
  wire alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
  wire alu_loop_op_7_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0;
  wire alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
  wire alu_loop_op_8_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0;
  wire alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
  wire alu_loop_op_9_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0;
  wire alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
  wire alu_loop_op_10_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0;
  wire alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
  wire alu_loop_op_11_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0;
  wire alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
  wire alu_loop_op_12_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0;
  wire alu_loop_op_13_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0;
  wire alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
  wire alu_loop_op_14_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0;
  wire alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
  wire alu_loop_op_15_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0;
  wire alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
  wire alu_loop_op_16_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0;
  wire alu_loop_op_4_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm_mx0w0;
  wire alu_loop_op_4_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm_mx0w0;
  wire alu_loop_op_6_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm_mx0w0;
  wire alu_loop_op_6_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm_mx0w0;
  wire alu_loop_op_13_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_itm_mx0w0;
  wire alu_loop_op_13_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_itm_mx0w0;
  wire FpAlu_8U_23U_or_831_itm_mx0w0;
  wire FpAlu_8U_23U_or_752_itm_mx0w0;
  wire FpAlu_8U_23U_or_833_itm_mx0w0;
  wire FpAlu_8U_23U_or_755_itm_mx0w0;
  wire FpAlu_8U_23U_or_835_itm_mx0w0;
  wire FpAlu_8U_23U_or_758_itm_mx0w0;
  wire FpAlu_8U_23U_or_837_itm_mx0w0;
  wire FpAlu_8U_23U_or_761_itm_mx0w0;
  wire FpAlu_8U_23U_or_839_itm_mx0w0;
  wire FpAlu_8U_23U_or_764_itm_mx0w0;
  wire FpAlu_8U_23U_or_841_itm_mx0w0;
  wire FpAlu_8U_23U_or_767_itm_mx0w0;
  wire FpAlu_8U_23U_or_843_itm_mx0w0;
  wire FpAlu_8U_23U_or_770_itm_mx0w0;
  wire FpAlu_8U_23U_or_845_itm_mx0w0;
  wire FpAlu_8U_23U_or_773_itm_mx0w0;
  wire FpAlu_8U_23U_or_847_itm_mx0w0;
  wire FpAlu_8U_23U_or_776_itm_mx0w0;
  wire FpAlu_8U_23U_or_849_itm_mx0w0;
  wire FpAlu_8U_23U_or_779_itm_mx0w0;
  wire FpAlu_8U_23U_or_851_itm_mx0w0;
  wire FpAlu_8U_23U_or_782_itm_mx0w0;
  wire FpAlu_8U_23U_or_853_itm_mx0w0;
  wire FpAlu_8U_23U_or_785_itm_mx0w0;
  wire FpAlu_8U_23U_or_855_itm_mx0w0;
  wire FpAlu_8U_23U_or_788_itm_mx0w0;
  wire FpAlu_8U_23U_or_857_itm_mx0w0;
  wire FpAlu_8U_23U_or_791_itm_mx0w0;
  wire FpAlu_8U_23U_or_859_itm_mx0w0;
  wire FpAlu_8U_23U_or_794_itm_mx0w0;
  wire FpAlu_8U_23U_or_861_itm_mx0w0;
  wire FpAlu_8U_23U_or_797_itm_mx0w0;
  wire FpAlu_8U_23U_and_itm_mx0w0;
  wire FpAlu_8U_23U_and_4_itm_mx0w0;
  wire FpAlu_8U_23U_and_8_itm_mx0w0;
  wire FpAlu_8U_23U_and_12_itm_mx0w0;
  wire FpAlu_8U_23U_and_16_itm_mx0w0;
  wire FpAlu_8U_23U_and_20_itm_mx0w0;
  wire FpAlu_8U_23U_and_24_itm_mx0w0;
  wire FpAlu_8U_23U_and_28_itm_mx0w0;
  wire FpAlu_8U_23U_and_32_itm_mx0w0;
  wire FpAlu_8U_23U_and_36_itm_mx0w0;
  wire FpAlu_8U_23U_and_40_itm_mx0w0;
  wire FpAlu_8U_23U_and_44_itm_mx0w0;
  wire FpAlu_8U_23U_and_48_itm_mx0w0;
  wire FpAlu_8U_23U_and_52_itm_mx0w0;
  wire FpAlu_8U_23U_and_56_itm_mx0w0;
  wire FpAlu_8U_23U_and_60_itm_mx0w0;
  wire FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_mx0w0;
  wire FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_mx0w1;
  wire FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_mx0w2;
  wire FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_mx0w3;
  wire FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w4;
  wire FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_1_mx0w0;
  wire FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_1_mx0w1;
  wire FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_1_mx0w2;
  wire FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_1_mx0w3;
  wire FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w4;
  wire FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_2_mx0w0;
  wire FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_2_mx0w1;
  wire FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_2_mx0w2;
  wire FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_2_mx0w3;
  wire FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w4;
  wire FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_3_mx0w0;
  wire FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_3_mx0w1;
  wire FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_3_mx0w2;
  wire FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_3_mx0w3;
  wire FpAdd_8U_23U_is_a_greater_lor_4_lpi_1_dfm_1_mx0w4;
  wire FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_4_mx0w0;
  wire FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_4_mx0w1;
  wire FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_4_mx0w2;
  wire FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_4_mx0w3;
  wire FpAdd_8U_23U_is_a_greater_lor_5_lpi_1_dfm_1_mx0w4;
  wire FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_5_mx0w0;
  wire FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_5_mx0w1;
  wire FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_5_mx0w2;
  wire FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_5_mx0w3;
  wire FpAdd_8U_23U_is_a_greater_lor_6_lpi_1_dfm_1_mx0w4;
  wire FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_6_mx0w0;
  wire FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_6_mx0w1;
  wire FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_6_mx0w2;
  wire FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_6_mx0w3;
  wire FpAdd_8U_23U_is_a_greater_lor_7_lpi_1_dfm_1_mx0w4;
  wire FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_7_mx0w0;
  wire FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_7_mx0w1;
  wire FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_7_mx0w2;
  wire FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_7_mx0w3;
  wire FpAdd_8U_23U_is_a_greater_lor_8_lpi_1_dfm_1_mx0w4;
  wire FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_8_mx0w0;
  wire FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_8_mx0w1;
  wire FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_8_mx0w2;
  wire FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_8_mx0w3;
  wire FpAdd_8U_23U_is_a_greater_lor_9_lpi_1_dfm_1_mx0w4;
  wire FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_9_mx0w0;
  wire FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_9_mx0w1;
  wire FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_9_mx0w2;
  wire FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_9_mx0w3;
  wire FpAdd_8U_23U_is_a_greater_lor_10_lpi_1_dfm_1_mx0w4;
  wire FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_10_mx0w0;
  wire FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_10_mx0w1;
  wire FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_10_mx0w2;
  wire FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_10_mx0w3;
  wire FpAdd_8U_23U_is_a_greater_lor_11_lpi_1_dfm_1_mx0w4;
  wire FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_11_mx0w0;
  wire FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_11_mx0w1;
  wire FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_11_mx0w2;
  wire FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_11_mx0w3;
  wire FpAdd_8U_23U_is_a_greater_lor_12_lpi_1_dfm_1_mx0w4;
  wire FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_12_mx0w0;
  wire FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_12_mx0w1;
  wire FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_12_mx0w2;
  wire FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_12_mx0w3;
  wire FpAdd_8U_23U_is_a_greater_lor_13_lpi_1_dfm_1_mx0w4;
  wire FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_13_mx0w0;
  wire FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_13_mx0w1;
  wire FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_13_mx0w2;
  wire FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_13_mx0w3;
  wire FpAdd_8U_23U_is_a_greater_lor_14_lpi_1_dfm_1_mx0w4;
  wire FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_14_mx0w0;
  wire FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_14_mx0w1;
  wire FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_14_mx0w2;
  wire FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_14_mx0w3;
  wire FpAdd_8U_23U_is_a_greater_lor_15_lpi_1_dfm_1_mx0w4;
  wire FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_15_mx0w0;
  wire FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_15_mx0w1;
  wire FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_15_mx0w2;
  wire FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_15_mx0w3;
  wire FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w4;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_65_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_64_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_67_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_66_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_69_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_68_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_71_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_70_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_73_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_72_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_75_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_74_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_77_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_76_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_79_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_78_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_81_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_80_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_83_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_82_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_85_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_84_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_87_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_86_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_89_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_88_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_91_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_90_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_93_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_92_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_95_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_94_mx0w1;
  wire IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_3_land_15_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_3_land_14_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_3_land_13_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_3_land_12_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_3_land_11_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_3_land_10_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_3_land_9_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_3_land_8_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_3_land_7_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_3_land_6_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_3_land_5_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_3_land_4_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_3_land_3_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_3_land_2_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_3_land_1_lpi_1_dfm_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_0_1_sva_mx0w0;
  wire [29:0] IntShiftLeft_16U_6U_32U_return_30_1_1_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_31_1_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_0_2_sva_mx0w0;
  wire [29:0] IntShiftLeft_16U_6U_32U_return_30_1_2_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_31_2_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_0_3_sva_mx0w0;
  wire [29:0] IntShiftLeft_16U_6U_32U_return_30_1_3_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_31_3_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_0_4_sva_mx0w0;
  wire [29:0] IntShiftLeft_16U_6U_32U_return_30_1_4_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_31_4_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_0_5_sva_mx0w0;
  wire [29:0] IntShiftLeft_16U_6U_32U_return_30_1_5_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_31_5_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_0_6_sva_mx0w0;
  wire [29:0] IntShiftLeft_16U_6U_32U_return_30_1_6_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_31_6_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_0_7_sva_mx0w0;
  wire [29:0] IntShiftLeft_16U_6U_32U_return_30_1_7_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_31_7_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_0_8_sva_mx0w0;
  wire [29:0] IntShiftLeft_16U_6U_32U_return_30_1_8_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_31_8_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_0_9_sva_mx0w0;
  wire [29:0] IntShiftLeft_16U_6U_32U_return_30_1_9_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_31_9_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_0_10_sva_mx0w0;
  wire [29:0] IntShiftLeft_16U_6U_32U_return_30_1_10_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_31_10_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_0_11_sva_mx0w0;
  wire [29:0] IntShiftLeft_16U_6U_32U_return_30_1_11_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_31_11_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_0_12_sva_mx0w0;
  wire [29:0] IntShiftLeft_16U_6U_32U_return_30_1_12_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_31_12_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_0_13_sva_mx0w0;
  wire [29:0] IntShiftLeft_16U_6U_32U_return_30_1_13_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_31_13_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_0_14_sva_mx0w0;
  wire [29:0] IntShiftLeft_16U_6U_32U_return_30_1_14_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_31_14_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_0_15_sva_mx0w0;
  wire [29:0] IntShiftLeft_16U_6U_32U_return_30_1_15_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_31_15_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_0_sva_mx0w0;
  wire [29:0] IntShiftLeft_16U_6U_32U_return_30_1_sva_mx0w0;
  wire IntShiftLeft_16U_6U_32U_return_31_sva_mx0w0;
  wire alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  wire alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  wire alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  wire alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  wire alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  wire alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  wire alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  wire alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  wire alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  wire alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  wire alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  wire alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  wire alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  wire alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  wire alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  wire alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  wire IsNaN_8U_23U_2_land_lpi_1_dfm_mx1w0;
  wire IsNaN_8U_23U_2_land_15_lpi_1_dfm_mx1w0;
  wire IsNaN_8U_23U_2_land_14_lpi_1_dfm_mx1w0;
  wire IsNaN_8U_23U_2_land_13_lpi_1_dfm_mx1w0;
  wire IsNaN_8U_23U_2_land_12_lpi_1_dfm_mx1w0;
  wire IsNaN_8U_23U_2_land_11_lpi_1_dfm_mx1w0;
  wire IsNaN_8U_23U_2_land_10_lpi_1_dfm_mx1w0;
  wire IsNaN_8U_23U_2_land_9_lpi_1_dfm_mx1w0;
  wire IsNaN_8U_23U_2_land_8_lpi_1_dfm_mx1w0;
  wire IsNaN_8U_23U_2_land_7_lpi_1_dfm_mx1w0;
  wire IsNaN_8U_23U_2_land_6_lpi_1_dfm_mx1w0;
  wire IsNaN_8U_23U_2_land_5_lpi_1_dfm_mx1w0;
  wire IsNaN_8U_23U_2_land_4_lpi_1_dfm_mx1w0;
  wire IsNaN_8U_23U_2_land_3_lpi_1_dfm_mx1w0;
  wire IsNaN_8U_23U_2_land_2_lpi_1_dfm_mx1w0;
  wire IsNaN_8U_23U_2_land_1_lpi_1_dfm_mx1w0;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_1_sva;
  wire [50:0] nl_FpAdd_8U_23U_int_mant_p1_1_sva;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_91_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_1_sva;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_2_sva;
  wire [50:0] nl_FpAdd_8U_23U_int_mant_p1_2_sva;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_85_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_2_sva;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_3_sva;
  wire [50:0] nl_FpAdd_8U_23U_int_mant_p1_3_sva;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_79_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_3_sva;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_4_sva;
  wire [50:0] nl_FpAdd_8U_23U_int_mant_p1_4_sva;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_73_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_4_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_4_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_4_sva;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_5_sva;
  wire [50:0] nl_FpAdd_8U_23U_int_mant_p1_5_sva;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_67_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_5_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_5_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_5_sva;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_6_sva;
  wire [50:0] nl_FpAdd_8U_23U_int_mant_p1_6_sva;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_61_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_6_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_6_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_6_sva;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_7_sva;
  wire [50:0] nl_FpAdd_8U_23U_int_mant_p1_7_sva;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_55_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_7_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_7_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_7_sva;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_8_sva;
  wire [50:0] nl_FpAdd_8U_23U_int_mant_p1_8_sva;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_49_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_8_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_8_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_8_sva;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_9_sva;
  wire [50:0] nl_FpAdd_8U_23U_int_mant_p1_9_sva;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_43_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_9_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_9_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_9_sva;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_10_sva;
  wire [50:0] nl_FpAdd_8U_23U_int_mant_p1_10_sva;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_37_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_10_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_10_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_10_sva;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_11_sva;
  wire [50:0] nl_FpAdd_8U_23U_int_mant_p1_11_sva;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_31_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_11_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_11_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_11_sva;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_12_sva;
  wire [50:0] nl_FpAdd_8U_23U_int_mant_p1_12_sva;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_25_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_12_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_12_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_12_sva;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_13_sva;
  wire [50:0] nl_FpAdd_8U_23U_int_mant_p1_13_sva;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_19_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_13_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_13_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_13_sva;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_14_sva;
  wire [50:0] nl_FpAdd_8U_23U_int_mant_p1_14_sva;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_13_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_14_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_14_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_14_sva;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_15_sva;
  wire [50:0] nl_FpAdd_8U_23U_int_mant_p1_15_sva;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_7_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_15_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_15_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_15_sva;
  wire [49:0] FpAdd_8U_23U_int_mant_p1_sva;
  wire [50:0] nl_FpAdd_8U_23U_int_mant_p1_sva;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_1_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_sva;
  wire [22:0] FpAdd_8U_23U_o_mant_1_lpi_1_dfm_2_mx0;
  wire [22:0] FpAdd_8U_23U_o_mant_2_lpi_1_dfm_2_mx0;
  wire [22:0] FpAdd_8U_23U_o_mant_3_lpi_1_dfm_2_mx0;
  wire [22:0] FpAdd_8U_23U_o_mant_4_lpi_1_dfm_2_mx0;
  wire [22:0] FpAdd_8U_23U_o_mant_5_lpi_1_dfm_2_mx0;
  wire [22:0] FpAdd_8U_23U_o_mant_6_lpi_1_dfm_2_mx0;
  wire [22:0] FpAdd_8U_23U_o_mant_7_lpi_1_dfm_2_mx0;
  wire [22:0] FpAdd_8U_23U_o_mant_8_lpi_1_dfm_2_mx0;
  wire [22:0] FpAdd_8U_23U_o_mant_9_lpi_1_dfm_2_mx0;
  wire [22:0] FpAdd_8U_23U_o_mant_10_lpi_1_dfm_2_mx0;
  wire [22:0] FpAdd_8U_23U_o_mant_11_lpi_1_dfm_2_mx0;
  wire [22:0] FpAdd_8U_23U_o_mant_12_lpi_1_dfm_2_mx0;
  wire [22:0] FpAdd_8U_23U_o_mant_13_lpi_1_dfm_2_mx0;
  wire [22:0] FpAdd_8U_23U_o_mant_14_lpi_1_dfm_2_mx0;
  wire [22:0] FpAdd_8U_23U_o_mant_15_lpi_1_dfm_2_mx0;
  wire [22:0] FpAdd_8U_23U_o_mant_lpi_1_dfm_2_mx0;
  wire [7:0] FpAdd_8U_23U_o_expo_1_lpi_1_dfm_1;
  wire [48:0] FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0;
  wire FpMantRNE_49U_24U_else_carry_1_sva;
  wire [7:0] FpAdd_8U_23U_o_expo_2_lpi_1_dfm_1;
  wire [48:0] FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0;
  wire FpMantRNE_49U_24U_else_carry_2_sva;
  wire [7:0] FpAdd_8U_23U_o_expo_3_lpi_1_dfm_1;
  wire [48:0] FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0;
  wire FpMantRNE_49U_24U_else_carry_3_sva;
  wire [7:0] FpAdd_8U_23U_o_expo_4_lpi_1_dfm_1;
  wire [48:0] FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0;
  wire FpMantRNE_49U_24U_else_carry_4_sva;
  wire [7:0] FpAdd_8U_23U_o_expo_5_lpi_1_dfm_1;
  wire [48:0] FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0;
  wire FpMantRNE_49U_24U_else_carry_5_sva;
  wire [7:0] FpAdd_8U_23U_o_expo_6_lpi_1_dfm_1;
  wire [48:0] FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0;
  wire FpMantRNE_49U_24U_else_carry_6_sva;
  wire [7:0] FpAdd_8U_23U_o_expo_7_lpi_1_dfm_1;
  wire [48:0] FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0;
  wire FpMantRNE_49U_24U_else_carry_7_sva;
  wire [7:0] FpAdd_8U_23U_o_expo_8_lpi_1_dfm_1;
  wire [48:0] FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0;
  wire FpMantRNE_49U_24U_else_carry_8_sva;
  wire [7:0] FpAdd_8U_23U_o_expo_9_lpi_1_dfm_1;
  wire [48:0] FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0;
  wire FpMantRNE_49U_24U_else_carry_9_sva;
  wire [7:0] FpAdd_8U_23U_o_expo_10_lpi_1_dfm_1;
  wire [48:0] FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0;
  wire FpMantRNE_49U_24U_else_carry_10_sva;
  wire [7:0] FpAdd_8U_23U_o_expo_11_lpi_1_dfm_1;
  wire [48:0] FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0;
  wire FpMantRNE_49U_24U_else_carry_11_sva;
  wire [7:0] FpAdd_8U_23U_o_expo_12_lpi_1_dfm_1;
  wire [48:0] FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0;
  wire FpMantRNE_49U_24U_else_carry_12_sva;
  wire [7:0] FpAdd_8U_23U_o_expo_13_lpi_1_dfm_1;
  wire [48:0] FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0;
  wire FpMantRNE_49U_24U_else_carry_13_sva;
  wire [7:0] FpAdd_8U_23U_o_expo_14_lpi_1_dfm_1;
  wire [48:0] FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0;
  wire FpMantRNE_49U_24U_else_carry_14_sva;
  wire [7:0] FpAdd_8U_23U_o_expo_15_lpi_1_dfm_1;
  wire [48:0] FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0;
  wire FpMantRNE_49U_24U_else_carry_15_sva;
  wire [7:0] FpAdd_8U_23U_o_expo_lpi_1_dfm_1;
  wire [48:0] FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0;
  wire FpMantRNE_49U_24U_else_carry_sva;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_1_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_1_sva;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_2_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_2_sva;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_3_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_3_sva;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_4_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_4_sva;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_5_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_5_sva;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_6_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_6_sva;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_7_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_7_sva;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_8_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_8_sva;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_9_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_9_sva;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_10_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_10_sva;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_11_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_11_sva;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_12_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_12_sva;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_13_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_13_sva;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_14_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_14_sva;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_15_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_15_sva;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_sva;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_30_ssc;
  wire IsNaN_5U_23U_land_lpi_1_dfm;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_28_ssc;
  wire IsNaN_5U_23U_land_15_lpi_1_dfm;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_26_ssc;
  wire IsNaN_5U_23U_land_14_lpi_1_dfm;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_24_ssc;
  wire IsNaN_5U_23U_land_13_lpi_1_dfm;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_22_ssc;
  wire IsNaN_5U_23U_land_12_lpi_1_dfm;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_20_ssc;
  wire IsNaN_5U_23U_land_11_lpi_1_dfm;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_18_ssc;
  wire IsNaN_5U_23U_land_10_lpi_1_dfm;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_16_ssc;
  wire IsNaN_5U_23U_land_9_lpi_1_dfm;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_ssc;
  wire IsNaN_5U_23U_land_8_lpi_1_dfm;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_ssc;
  wire IsNaN_5U_23U_land_7_lpi_1_dfm;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_ssc;
  wire IsNaN_5U_23U_land_6_lpi_1_dfm;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_ssc;
  wire IsNaN_5U_23U_land_5_lpi_1_dfm;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_ssc;
  wire IsNaN_5U_23U_land_4_lpi_1_dfm;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_ssc;
  wire IsNaN_5U_23U_land_3_lpi_1_dfm;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_ssc;
  wire IsNaN_5U_23U_land_2_lpi_1_dfm;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_ssc;
  wire IsNaN_5U_23U_land_1_lpi_1_dfm;
  wire or_4_cse;
  wire or_5_cse;
  wire or_6_cse;
  wire or_7_cse;
  wire or_8_cse;
  wire or_9_cse;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_4_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_4_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_5_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_5_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_6_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_6_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_7_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_7_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_8_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_8_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_9_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_9_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_10_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_10_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_11_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_11_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_12_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_12_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_13_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_13_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_14_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_14_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_15_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_15_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_sva_2;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_sva_2;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_sva_2;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_sva_2;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_sva_2;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_sva_2;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_sva_2;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_sva_2;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_sva_2;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_sva_2;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_sva_2;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_sva_2;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_sva_2;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_sva_2;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_sva_2;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_sva_2;
  wire FpCmp_8U_23U_true_is_abs_a_greater_1_lpi_1_dfm_1;
  wire FpCmp_8U_23U_false_is_abs_a_greater_1_lpi_1_dfm_1;
  wire FpCmp_8U_23U_true_is_abs_a_greater_2_lpi_1_dfm_1;
  wire FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_1;
  wire FpCmp_8U_23U_true_is_abs_a_greater_3_lpi_1_dfm_1;
  wire FpCmp_8U_23U_false_is_abs_a_greater_3_lpi_1_dfm_1;
  wire FpCmp_8U_23U_true_is_abs_a_greater_4_lpi_1_dfm_1;
  wire FpCmp_8U_23U_false_is_abs_a_greater_4_lpi_1_dfm_1;
  wire FpCmp_8U_23U_true_is_abs_a_greater_5_lpi_1_dfm_1;
  wire FpCmp_8U_23U_false_is_abs_a_greater_5_lpi_1_dfm_1;
  wire FpCmp_8U_23U_true_is_abs_a_greater_6_lpi_1_dfm_1;
  wire FpCmp_8U_23U_false_is_abs_a_greater_6_lpi_1_dfm_1;
  wire FpCmp_8U_23U_true_is_abs_a_greater_7_lpi_1_dfm_1;
  wire FpCmp_8U_23U_false_is_abs_a_greater_7_lpi_1_dfm_1;
  wire FpCmp_8U_23U_true_is_abs_a_greater_8_lpi_1_dfm_1;
  wire FpCmp_8U_23U_false_is_abs_a_greater_8_lpi_1_dfm_1;
  wire FpCmp_8U_23U_true_is_abs_a_greater_9_lpi_1_dfm_1;
  wire FpCmp_8U_23U_false_is_abs_a_greater_9_lpi_1_dfm_1;
  wire FpCmp_8U_23U_true_is_abs_a_greater_10_lpi_1_dfm_1;
  wire FpCmp_8U_23U_false_is_abs_a_greater_10_lpi_1_dfm_1;
  wire FpCmp_8U_23U_true_is_abs_a_greater_11_lpi_1_dfm_1;
  wire FpCmp_8U_23U_false_is_abs_a_greater_11_lpi_1_dfm_1;
  wire FpCmp_8U_23U_true_is_abs_a_greater_12_lpi_1_dfm_1;
  wire FpCmp_8U_23U_false_is_abs_a_greater_12_lpi_1_dfm_1;
  wire FpCmp_8U_23U_true_is_abs_a_greater_13_lpi_1_dfm_1;
  wire FpCmp_8U_23U_false_is_abs_a_greater_13_lpi_1_dfm_1;
  wire FpCmp_8U_23U_true_is_abs_a_greater_14_lpi_1_dfm_1;
  wire FpCmp_8U_23U_false_is_abs_a_greater_14_lpi_1_dfm_1;
  wire FpCmp_8U_23U_true_is_abs_a_greater_15_lpi_1_dfm_1;
  wire FpCmp_8U_23U_false_is_abs_a_greater_15_lpi_1_dfm_1;
  wire FpCmp_8U_23U_true_is_abs_a_greater_lpi_1_dfm_1;
  wire FpCmp_8U_23U_false_is_abs_a_greater_lpi_1_dfm_1;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_15_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_15_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_14_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_14_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_13_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_13_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_12_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_12_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_11_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_11_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_10_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_10_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_9_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_9_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_8_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_8_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_7_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_7_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_6_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_6_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_5_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_5_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_4_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_4_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_3_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_3_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_2_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_2_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_1_sva;
  wire IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_1_sva;
  wire FpNormalize_8U_49U_oelse_not_33;
  wire FpAdd_8U_23U_asn_256;
  wire FpAdd_8U_23U_asn_258;
  wire FpNormalize_8U_49U_oelse_not_35;
  wire FpAdd_8U_23U_asn_260;
  wire FpAdd_8U_23U_asn_262;
  wire FpNormalize_8U_49U_oelse_not_37;
  wire FpAdd_8U_23U_asn_264;
  wire FpAdd_8U_23U_asn_266;
  wire FpNormalize_8U_49U_oelse_not_39;
  wire FpAdd_8U_23U_asn_268;
  wire FpAdd_8U_23U_asn_270;
  wire FpNormalize_8U_49U_oelse_not_41;
  wire FpAdd_8U_23U_asn_272;
  wire FpAdd_8U_23U_asn_274;
  wire FpNormalize_8U_49U_oelse_not_43;
  wire FpAdd_8U_23U_asn_276;
  wire FpAdd_8U_23U_asn_278;
  wire FpNormalize_8U_49U_oelse_not_45;
  wire FpAdd_8U_23U_asn_280;
  wire FpAdd_8U_23U_asn_282;
  wire FpNormalize_8U_49U_oelse_not_47;
  wire FpAdd_8U_23U_asn_284;
  wire FpAdd_8U_23U_asn_286;
  wire FpNormalize_8U_49U_oelse_not_49;
  wire FpAdd_8U_23U_asn_288;
  wire FpAdd_8U_23U_asn_290;
  wire FpNormalize_8U_49U_oelse_not_51;
  wire FpAdd_8U_23U_asn_292;
  wire FpAdd_8U_23U_asn_294;
  wire FpNormalize_8U_49U_oelse_not_53;
  wire FpAdd_8U_23U_asn_296;
  wire FpAdd_8U_23U_asn_298;
  wire FpNormalize_8U_49U_oelse_not_55;
  wire FpAdd_8U_23U_asn_300;
  wire FpAdd_8U_23U_asn_302;
  wire FpNormalize_8U_49U_oelse_not_57;
  wire FpAdd_8U_23U_asn_304;
  wire FpAdd_8U_23U_asn_306;
  wire FpNormalize_8U_49U_oelse_not_59;
  wire FpAdd_8U_23U_asn_308;
  wire FpAdd_8U_23U_asn_310;
  wire FpNormalize_8U_49U_oelse_not_61;
  wire FpAdd_8U_23U_asn_312;
  wire FpAdd_8U_23U_asn_314;
  wire FpNormalize_8U_49U_oelse_not_63;
  wire FpAdd_8U_23U_asn_316;
  wire FpAdd_8U_23U_asn_318;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_16;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_17;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_18;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_19;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_20;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_21;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_22;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_23;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_24;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_25;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_26;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_27;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_28;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_29;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_30;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_31;
  wire [5:0] libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_16;
  wire [5:0] libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_17;
  wire [5:0] libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_18;
  wire [5:0] libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_19;
  wire [5:0] libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_20;
  wire [5:0] libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_21;
  wire [5:0] libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_22;
  wire [5:0] libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_23;
  wire [5:0] libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_24;
  wire [5:0] libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_25;
  wire [5:0] libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_26;
  wire [5:0] libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_27;
  wire [5:0] libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_28;
  wire [5:0] libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_29;
  wire [5:0] libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_30;
  wire [5:0] libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_31;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp_2;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp_2;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_95_ssc;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_tmp_2;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_94_ssc;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_tmp_2;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_93_ssc;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_tmp_2;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_92_ssc;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_tmp_2;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_91_ssc;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_tmp_2;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_90_ssc;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_tmp_2;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_89_ssc;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_tmp_2;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_88_ssc;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_tmp_2;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_87_ssc;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_tmp_2;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_86_ssc;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_tmp_2;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_85_ssc;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_tmp_2;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_84_ssc;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_tmp_2;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_83_ssc;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_tmp_2;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_82_ssc;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_tmp_2;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_81_ssc;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_tmp_2;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_80_ssc;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_tmp;
  reg [2:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_tmp_1;
  reg [9:0] reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_tmp_2;
  wire AluIn_data_and_1_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_cse;
  wire FpAdd_8U_23U_is_a_greater_oelse_FpAdd_8U_23U_is_a_greater_oelse_or_21_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_75_cse;
  wire FpAdd_8U_23U_b_left_shift_and_32_cse;
  wire IsZero_8U_23U_1_and_cse;
  wire FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_78_cse;
  wire AluIn_data_and_2_cse;
  wire alu_loop_op_else_else_if_and_57_cse;
  wire alu_loop_op_else_else_if_and_60_cse;
  wire alu_loop_op_else_else_if_and_66_cse;
  wire FpAlu_8U_23U_and_832_cse;
  wire FpAdd_8U_23U_and_176_cse;
  wire IsNaN_8U_23U_aelse_and_16_cse;
  wire FpAdd_8U_23U_and_178_cse;
  wire IsNaN_8U_23U_aelse_and_18_cse;
  wire FpAdd_8U_23U_and_180_cse;
  wire FpAdd_8U_23U_and_182_cse;
  wire FpAdd_8U_23U_and_184_cse;
  wire IsNaN_8U_23U_aelse_and_24_cse;
  wire FpAdd_8U_23U_and_186_cse;
  wire FpAdd_8U_23U_and_188_cse;
  wire FpAdd_8U_23U_and_190_cse;
  wire FpAdd_8U_23U_and_192_cse;
  wire FpAdd_8U_23U_and_194_cse;
  wire FpAdd_8U_23U_and_196_cse;
  wire IsNaN_8U_23U_aelse_and_36_cse;
  wire FpAdd_8U_23U_and_198_cse;
  wire FpAdd_8U_23U_and_200_cse;
  wire FpAdd_8U_23U_and_202_cse;
  wire FpAdd_8U_23U_and_204_cse;
  wire FpAdd_8U_23U_and_206_cse;
  wire AluIn_data_and_3_cse;
  wire FpAlu_8U_23U_and_849_cse;
  wire cfg_alu_algo_and_115_cse;
  wire FpAlu_8U_23U_and_889_cse;
  wire IsNaN_8U_23U_aelse_IsNaN_8U_23U_2_aelse_or_15_cse;
  wire FpAdd_8U_23U_and_208_cse;
  wire FpNormalize_8U_49U_if_and_31_cse;
  wire FpAdd_8U_23U_and_210_cse;
  wire FpNormalize_8U_49U_if_and_32_cse;
  wire FpAdd_8U_23U_and_212_cse;
  wire FpNormalize_8U_49U_if_and_33_cse;
  wire FpAdd_8U_23U_and_214_cse;
  wire FpNormalize_8U_49U_if_and_34_cse;
  wire FpNormalize_8U_49U_if_and_35_cse;
  wire FpNormalize_8U_49U_if_and_36_cse;
  wire FpNormalize_8U_49U_if_and_37_cse;
  wire FpAdd_8U_23U_and_216_cse;
  wire FpNormalize_8U_49U_if_and_38_cse;
  wire FpNormalize_8U_49U_if_and_39_cse;
  wire FpNormalize_8U_49U_if_and_40_cse;
  wire FpNormalize_8U_49U_if_and_41_cse;
  wire FpNormalize_8U_49U_if_and_42_cse;
  wire FpAdd_8U_23U_and_218_cse;
  wire FpNormalize_8U_49U_if_and_43_cse;
  wire FpAdd_8U_23U_and_220_cse;
  wire FpNormalize_8U_49U_if_and_44_cse;
  wire FpAdd_8U_23U_and_222_cse;
  wire FpNormalize_8U_49U_if_and_45_cse;
  wire FpAdd_8U_23U_and_224_cse;
  wire FpNormalize_8U_49U_if_and_46_cse;
  wire FpAdd_8U_23U_and_226_cse;
  wire FpAdd_8U_23U_and_228_cse;
  wire FpAdd_8U_23U_and_230_cse;
  wire FpAdd_8U_23U_and_232_cse;
  wire FpAdd_8U_23U_and_234_cse;
  wire FpAdd_8U_23U_and_236_cse;
  wire FpAdd_8U_23U_and_238_cse;
  wire IsNaN_8U_23U_1_aelse_and_34_cse;
  wire alu_loop_op_else_else_if_and_105_cse;
  wire alu_loop_op_else_else_if_and_108_cse;
  wire alu_loop_op_else_else_if_and_111_cse;
  wire alu_loop_op_else_else_if_and_114_cse;
  wire alu_loop_op_else_else_if_and_117_cse;
  wire alu_loop_op_else_else_if_and_120_cse;
  wire alu_loop_op_else_else_if_and_123_cse;
  wire alu_loop_op_else_else_if_and_126_cse;
  wire alu_loop_op_else_else_if_and_129_cse;
  wire alu_loop_op_else_else_if_and_132_cse;
  wire alu_loop_op_else_else_if_and_135_cse;
  wire alu_loop_op_else_else_if_and_138_cse;
  wire alu_loop_op_else_else_if_and_141_cse;
  wire FpAlu_8U_23U_and_1040_cse;
  wire FpAlu_8U_23U_FpAlu_8U_23U_or_79_cse;
  wire alu_loop_op_else_else_if_and_144_cse;
  wire alu_loop_op_else_else_if_and_147_cse;
  wire alu_loop_op_else_else_if_and_150_cse;
  wire IsNaN_8U_23U_2_aelse_and_74_cse;
  wire FpAlu_8U_23U_and_1120_cse;
  wire cfg_alu_src_and_cse;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_cse;
  wire FpAdd_8U_23U_int_mant_p1_and_16_cse;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_16_cse;
  wire FpAdd_8U_23U_int_mant_p1_and_17_cse;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_17_cse;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_18_cse;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_19_cse;
  wire FpAdd_8U_23U_int_mant_p1_and_20_cse;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_20_cse;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_21_cse;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_22_cse;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_23_cse;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_24_cse;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_25_cse;
  wire FpAdd_8U_23U_int_mant_p1_and_26_cse;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_26_cse;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_27_cse;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_28_cse;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_29_cse;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_30_cse;
  wire FpAdd_8U_23U_is_a_greater_and_17_cse;
  wire FpAlu_8U_23U_and_976_cse;
  wire FpAlu_8U_23U_and_1056_cse;
  wire cfg_alu_algo_and_132_cse;
  wire alu_nan_to_zero_op_sign_and_25_cse;
  wire IntShiftLeft_16U_6U_32U_and_48_cse;
  wire IntShiftLeft_16U_6U_32U_and_93_cse;
  reg [1:0] reg_cfg_alu_algo_1_sva_st_93_cse;
  reg reg_alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse;
  reg reg_alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse;
  reg reg_alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse;
  reg reg_alu_loop_op_5_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse;
  reg reg_alu_loop_op_6_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse;
  reg reg_alu_loop_op_7_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse;
  reg reg_alu_loop_op_8_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse;
  reg reg_alu_loop_op_9_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse;
  reg reg_alu_loop_op_10_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse;
  reg reg_alu_loop_op_11_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse;
  reg reg_alu_loop_op_12_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse;
  reg reg_alu_loop_op_13_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse;
  reg reg_alu_loop_op_14_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse;
  reg reg_alu_loop_op_15_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse;
  reg reg_alu_loop_op_16_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse;
  wire FpCmp_8U_23U_false_if_and_cse;
  wire FpCmp_8U_23U_true_if_and_7_cse;
  wire mux_1631_cse;
  reg [1:0] reg_cfg_alu_algo_1_sva_st_157_cse;
  reg reg_alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse;
  wire or_338_cse;
  wire mux_157_cse;
  wire nor_1930_cse;
  wire nor_1928_cse;
  wire nor_1862_cse;
  wire nor_1815_cse;
  reg reg_FpAlu_8U_23U_or_797_cse;
  reg reg_FpAlu_8U_23U_or_794_cse;
  reg reg_FpAlu_8U_23U_or_791_cse;
  reg reg_FpAlu_8U_23U_or_788_cse;
  reg reg_FpAlu_8U_23U_or_785_cse;
  reg reg_FpAlu_8U_23U_or_782_cse;
  reg reg_FpAlu_8U_23U_or_779_cse;
  reg reg_FpAlu_8U_23U_or_776_cse;
  reg reg_FpAlu_8U_23U_or_773_cse;
  reg reg_FpAlu_8U_23U_or_770_cse;
  reg reg_FpAlu_8U_23U_or_767_cse;
  reg reg_FpAlu_8U_23U_or_764_cse;
  reg reg_FpAlu_8U_23U_or_761_cse;
  reg reg_FpAlu_8U_23U_or_758_cse;
  reg reg_FpAlu_8U_23U_or_755_cse;
  reg reg_FpAlu_8U_23U_or_752_cse;
  wire IsNaN_8U_23U_2_aelse_and_48_cse;
  wire and_1105_cse;
  wire nor_577_cse;
  wire mux_818_cse;
  wire or_1938_cse;
  wire and_1141_cse;
  wire and_1307_cse;
  wire and_1318_cse;
  wire FpCmp_8U_23U_true_if_and_cse;
  wire mux_1456_cse;
  wire nor_1743_cse;
  wire and_149_cse;
  wire and_150_cse;
  wire and_151_cse;
  wire and_152_cse;
  wire FpAdd_8U_23U_is_a_greater_oelse_and_17_cse;
  wire FpCmp_8U_23U_false_if_and_32_cse;
  wire FpCmp_8U_23U_false_if_and_39_cse;
  wire or_343_cse;
  reg [1:0] reg_cfg_alu_algo_1_sva_st_110_cse;
  wire mux_250_cse;
  wire mux_251_cse;
  wire mux_285_cse;
  wire AluOut_data_and_cse;
  wire FpAlu_8U_23U_o_and_cse;
  wire nor_326_cse;
  wire nor_1742_cse;
  wire IsZero_8U_23U_1_and_25_cse;
  wire IsZero_8U_23U_1_and_24_cse;
  wire IsNaN_8U_23U_1_aelse_or_5_cse;
  wire IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_1_aelse_or_5_cse;
  wire IsNaN_8U_23U_aelse_and_47_cse;
  wire mux_819_cse;
  wire mux_823_cse;
  wire mux_805_cse;
  wire mux_807_cse;
  wire mux_811_cse;
  wire nor_1312_cse;
  wire AluOut_data_and_16_cse;
  wire FpAlu_8U_23U_o_and_16_cse;
  wire mux_980_cse;
  wire mux_1082_cse;
  wire mux_1092_cse;
  wire and_1421_cse;
  wire FpCmp_8U_23U_false_if_and_49_cse;
  wire FpCmp_8U_23U_false_if_and_48_cse;
  wire or_1827_cse;
  wire or_1128_cse;
  wire FpAlu_8U_23U_or_863_cse;
  wire FpAlu_8U_23U_or_864_cse;
  wire FpAlu_8U_23U_or_865_cse;
  wire FpAlu_8U_23U_or_866_cse;
  wire FpAlu_8U_23U_or_867_cse;
  wire FpAlu_8U_23U_or_868_cse;
  wire FpAlu_8U_23U_or_869_cse;
  wire FpAlu_8U_23U_or_870_cse;
  wire FpAlu_8U_23U_or_871_cse;
  wire FpAlu_8U_23U_or_872_cse;
  wire FpAlu_8U_23U_or_873_cse;
  wire FpAlu_8U_23U_or_874_cse;
  wire FpAlu_8U_23U_or_875_cse;
  wire FpAlu_8U_23U_or_876_cse;
  wire FpAlu_8U_23U_or_877_cse;
  wire FpAlu_8U_23U_or_878_cse;
  wire FpAdd_8U_23U_is_addition_and_33_cse;
  wire FpAdd_8U_23U_is_addition_and_cse;
  wire nor_327_cse;
  wire IsNaN_8U_23U_aelse_and_cse;
  wire IsNaN_8U_23U_1_aelse_or_3_cse;
  wire IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_1_aelse_or_3_cse;
  wire IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_15_cse;
  wire IsNaN_8U_23U_3_aelse_and_2_cse;
  wire IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_13_cse;
  wire IsNaN_8U_23U_3_aelse_or_1_cse;
  wire IsNaN_8U_23U_3_aelse_and_5_cse;
  wire mux_1349_cse;
  wire or_878_cse;
  wire or_879_cse;
  wire mux_477_cse;
  wire xor_cse;
  wire FpAdd_8U_23U_if_3_and_cse;
  wire IsNaN_8U_23U_3_aelse_and_cse;
  wire IsNaN_8U_23U_3_aelse_and_1_cse;
  wire IsNaN_8U_23U_3_aelse_and_9_cse;
  wire alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
  wire alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
  wire alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
  wire alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
  wire alu_loop_op_5_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
  wire alu_loop_op_6_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
  wire alu_loop_op_7_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
  wire alu_loop_op_8_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
  wire alu_loop_op_9_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
  wire alu_loop_op_10_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
  wire alu_loop_op_11_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
  wire alu_loop_op_12_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
  wire alu_loop_op_13_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
  wire alu_loop_op_14_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
  wire alu_loop_op_15_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
  wire alu_loop_op_16_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_5_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_7_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_9_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_11_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_12_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_13_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_14_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_15_itm_23_1;
  wire alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1;
  wire alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1;
  wire alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1;
  wire alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1;
  wire alu_loop_op_5_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1;
  wire alu_loop_op_6_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1;
  wire alu_loop_op_7_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1;
  wire alu_loop_op_8_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1;
  wire alu_loop_op_9_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1;
  wire alu_loop_op_10_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1;
  wire alu_loop_op_11_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1;
  wire alu_loop_op_12_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1;
  wire alu_loop_op_13_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1;
  wire alu_loop_op_14_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1;
  wire alu_loop_op_15_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1;
  wire alu_loop_op_16_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1;
  wire FpCmp_8U_23U_false_else_else_if_acc_16_itm_23_1;
  wire FpCmp_8U_23U_false_else_if_acc_16_itm_8_1;
  wire FpCmp_8U_23U_false_else_else_if_acc_18_itm_23_1;
  wire FpCmp_8U_23U_false_else_if_acc_18_itm_8_1;
  wire FpCmp_8U_23U_false_else_else_if_acc_20_itm_23_1;
  wire FpCmp_8U_23U_false_else_if_acc_20_itm_8_1;
  wire FpCmp_8U_23U_false_else_else_if_acc_22_itm_23_1;
  wire FpCmp_8U_23U_false_else_if_acc_22_itm_8_1;
  wire FpCmp_8U_23U_false_else_else_if_acc_24_itm_23_1;
  wire FpCmp_8U_23U_false_else_if_acc_24_itm_8_1;
  wire FpCmp_8U_23U_false_else_else_if_acc_26_itm_23_1;
  wire FpCmp_8U_23U_false_else_if_acc_26_itm_8_1;
  wire FpCmp_8U_23U_false_else_else_if_acc_28_itm_23_1;
  wire FpCmp_8U_23U_false_else_if_acc_28_itm_8_1;
  wire FpCmp_8U_23U_false_else_else_if_acc_30_itm_23_1;
  wire FpCmp_8U_23U_false_else_if_acc_30_itm_8_1;
  wire FpCmp_8U_23U_false_else_else_if_acc_32_itm_23_1;
  wire FpCmp_8U_23U_false_else_if_acc_32_itm_8_1;
  wire FpCmp_8U_23U_false_else_else_if_acc_34_itm_23_1;
  wire FpCmp_8U_23U_false_else_if_acc_34_itm_8_1;
  wire FpCmp_8U_23U_false_else_else_if_acc_36_itm_23_1;
  wire FpCmp_8U_23U_false_else_if_acc_36_itm_8_1;
  wire FpCmp_8U_23U_false_else_else_if_acc_38_itm_23_1;
  wire FpCmp_8U_23U_false_else_if_acc_38_itm_8_1;
  wire FpCmp_8U_23U_false_else_else_if_acc_40_itm_23_1;
  wire FpCmp_8U_23U_false_else_if_acc_40_itm_8_1;
  wire FpCmp_8U_23U_false_else_else_if_acc_42_itm_23_1;
  wire FpCmp_8U_23U_false_else_if_acc_42_itm_8_1;
  wire FpCmp_8U_23U_false_else_else_if_acc_44_itm_23_1;
  wire FpCmp_8U_23U_false_else_if_acc_44_itm_8_1;
  wire FpCmp_8U_23U_false_else_else_if_acc_46_itm_23_1;
  wire FpCmp_8U_23U_false_else_if_acc_46_itm_8_1;
  wire FpCmp_8U_23U_true_if_acc_16_itm_8_1;
  wire FpCmp_8U_23U_true_if_acc_18_itm_8_1;
  wire FpCmp_8U_23U_true_if_acc_20_itm_8_1;
  wire FpCmp_8U_23U_true_if_acc_22_itm_8_1;
  wire FpCmp_8U_23U_true_if_acc_24_itm_8_1;
  wire FpCmp_8U_23U_true_if_acc_26_itm_8_1;
  wire FpCmp_8U_23U_true_if_acc_28_itm_8_1;
  wire FpCmp_8U_23U_true_if_acc_30_itm_8_1;
  wire FpCmp_8U_23U_true_if_acc_32_itm_8_1;
  wire FpCmp_8U_23U_true_if_acc_34_itm_8_1;
  wire FpCmp_8U_23U_true_if_acc_36_itm_8_1;
  wire FpCmp_8U_23U_true_if_acc_38_itm_8_1;
  wire FpCmp_8U_23U_true_if_acc_40_itm_8_1;
  wire FpCmp_8U_23U_true_if_acc_42_itm_8_1;
  wire FpCmp_8U_23U_true_if_acc_44_itm_8_1;
  wire FpCmp_8U_23U_true_if_acc_46_itm_8_1;
  wire alu_loop_op_16_else_if_acc_1_itm_32_1;
  wire alu_loop_op_16_else_else_if_acc_1_itm_32_1;
  wire alu_loop_op_15_else_if_acc_itm_32_1;
  wire alu_loop_op_15_else_else_if_acc_itm_32_1;
  wire alu_loop_op_14_else_if_acc_1_itm_32_1;
  wire alu_loop_op_14_else_else_if_acc_1_itm_32_1;
  wire alu_loop_op_13_else_if_acc_itm_32_1;
  wire alu_loop_op_13_else_else_if_acc_itm_32_1;
  wire alu_loop_op_12_else_if_acc_1_itm_32_1;
  wire alu_loop_op_12_else_else_if_acc_1_itm_32_1;
  wire alu_loop_op_11_else_if_acc_itm_32_1;
  wire alu_loop_op_11_else_else_if_acc_itm_32_1;
  wire alu_loop_op_10_else_if_acc_1_itm_32_1;
  wire alu_loop_op_10_else_else_if_acc_1_itm_32_1;
  wire alu_loop_op_9_else_if_acc_itm_32_1;
  wire alu_loop_op_9_else_else_if_acc_itm_32_1;
  wire alu_loop_op_8_else_if_acc_1_itm_32_1;
  wire alu_loop_op_8_else_else_if_acc_1_itm_32_1;
  wire alu_loop_op_7_else_if_acc_itm_32_1;
  wire alu_loop_op_7_else_else_if_acc_itm_32_1;
  wire alu_loop_op_6_else_if_acc_1_itm_32_1;
  wire alu_loop_op_6_else_else_if_acc_1_itm_32_1;
  wire alu_loop_op_5_else_if_acc_itm_32_1;
  wire alu_loop_op_5_else_else_if_acc_itm_32_1;
  wire alu_loop_op_4_else_if_acc_1_itm_32_1;
  wire alu_loop_op_4_else_else_if_acc_1_itm_32_1;
  wire alu_loop_op_3_else_if_acc_itm_32_1;
  wire alu_loop_op_3_else_else_if_acc_itm_32_1;
  wire alu_loop_op_2_else_if_acc_1_itm_32_1;
  wire alu_loop_op_2_else_else_if_acc_1_itm_32_1;
  wire alu_loop_op_1_else_if_acc_itm_32_1;
  wire alu_loop_op_1_else_else_if_acc_itm_32_1;
  wire[0:0] iExpoWidth_oExpoWidth_prb;
  wire[0:0] iMantWidth_oMantWidth_prb;
  wire[0:0] iMantWidth_oMantWidth_prb_1;
  wire[0:0] iExpoWidth_oExpoWidth_prb_1;
  wire[0:0] iExpoWidth_oExpoWidth_prb_2;
  wire[0:0] iMantWidth_oMantWidth_prb_2;
  wire[0:0] iMantWidth_oMantWidth_prb_3;
  wire[0:0] iExpoWidth_oExpoWidth_prb_3;
  wire[0:0] iExpoWidth_oExpoWidth_prb_4;
  wire[0:0] iMantWidth_oMantWidth_prb_4;
  wire[0:0] iMantWidth_oMantWidth_prb_5;
  wire[0:0] iExpoWidth_oExpoWidth_prb_5;
  wire[0:0] iExpoWidth_oExpoWidth_prb_6;
  wire[0:0] iMantWidth_oMantWidth_prb_6;
  wire[0:0] iMantWidth_oMantWidth_prb_7;
  wire[0:0] iExpoWidth_oExpoWidth_prb_7;
  wire[0:0] iExpoWidth_oExpoWidth_prb_8;
  wire[0:0] iMantWidth_oMantWidth_prb_8;
  wire[0:0] iMantWidth_oMantWidth_prb_9;
  wire[0:0] iExpoWidth_oExpoWidth_prb_9;
  wire[0:0] iExpoWidth_oExpoWidth_prb_10;
  wire[0:0] iMantWidth_oMantWidth_prb_10;
  wire[0:0] iMantWidth_oMantWidth_prb_11;
  wire[0:0] iExpoWidth_oExpoWidth_prb_11;
  wire[0:0] iExpoWidth_oExpoWidth_prb_12;
  wire[0:0] iMantWidth_oMantWidth_prb_12;
  wire[0:0] iMantWidth_oMantWidth_prb_13;
  wire[0:0] iExpoWidth_oExpoWidth_prb_13;
  wire[0:0] iExpoWidth_oExpoWidth_prb_14;
  wire[0:0] iMantWidth_oMantWidth_prb_14;
  wire[0:0] iMantWidth_oMantWidth_prb_15;
  wire[0:0] iExpoWidth_oExpoWidth_prb_15;
  wire[0:0] iExpoWidth_oExpoWidth_prb_16;
  wire[0:0] iMantWidth_oMantWidth_prb_16;
  wire[0:0] iMantWidth_oMantWidth_prb_17;
  wire[0:0] iExpoWidth_oExpoWidth_prb_17;
  wire[0:0] iExpoWidth_oExpoWidth_prb_18;
  wire[0:0] iMantWidth_oMantWidth_prb_18;
  wire[0:0] iMantWidth_oMantWidth_prb_19;
  wire[0:0] iExpoWidth_oExpoWidth_prb_19;
  wire[0:0] iExpoWidth_oExpoWidth_prb_20;
  wire[0:0] iMantWidth_oMantWidth_prb_20;
  wire[0:0] iMantWidth_oMantWidth_prb_21;
  wire[0:0] iExpoWidth_oExpoWidth_prb_21;
  wire[0:0] iExpoWidth_oExpoWidth_prb_22;
  wire[0:0] iMantWidth_oMantWidth_prb_22;
  wire[0:0] iMantWidth_oMantWidth_prb_23;
  wire[0:0] iExpoWidth_oExpoWidth_prb_23;
  wire[0:0] iExpoWidth_oExpoWidth_prb_24;
  wire[0:0] iMantWidth_oMantWidth_prb_24;
  wire[0:0] iMantWidth_oMantWidth_prb_25;
  wire[0:0] iExpoWidth_oExpoWidth_prb_25;
  wire[0:0] iExpoWidth_oExpoWidth_prb_26;
  wire[0:0] iMantWidth_oMantWidth_prb_26;
  wire[0:0] iMantWidth_oMantWidth_prb_27;
  wire[0:0] iExpoWidth_oExpoWidth_prb_27;
  wire[0:0] iExpoWidth_oExpoWidth_prb_28;
  wire[0:0] iMantWidth_oMantWidth_prb_28;
  wire[0:0] iMantWidth_oMantWidth_prb_29;
  wire[0:0] iExpoWidth_oExpoWidth_prb_29;
  wire[0:0] iExpoWidth_oExpoWidth_prb_30;
  wire[0:0] iMantWidth_oMantWidth_prb_30;
  wire[0:0] iMantWidth_oMantWidth_prb_31;
  wire[0:0] iExpoWidth_oExpoWidth_prb_31;
  wire[21:0] FpAlu_8U_23U_and_3_nl;
  wire[21:0] FpAlu_8U_23U_mux1h_1039_nl;
  wire[0:0] FpAlu_8U_23U_not_80_nl;
  wire[3:0] FpAlu_8U_23U_and_2_nl;
  wire[3:0] FpAlu_8U_23U_mux1h_1040_nl;
  wire[0:0] FpAlu_8U_23U_and_610_nl;
  wire[0:0] FpAlu_8U_23U_and_611_nl;
  wire[0:0] FpAlu_8U_23U_and_612_nl;
  wire[0:0] FpAlu_8U_23U_not_114_nl;
  wire[0:0] and_4128_nl;
  wire[0:0] mux_1569_nl;
  wire[0:0] or_5091_nl;
  wire[0:0] nand_nl;
  wire[3:0] FpAlu_8U_23U_FpAlu_8U_23U_nor_16_nl;
  wire[3:0] FpAlu_8U_23U_nor_16_nl;
  wire[3:0] FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_15_nl;
  wire[0:0] and_4125_nl;
  wire[21:0] FpAlu_8U_23U_and_7_nl;
  wire[21:0] FpAlu_8U_23U_mux1h_1036_nl;
  wire[0:0] FpAlu_8U_23U_not_82_nl;
  wire[3:0] FpAlu_8U_23U_and_6_nl;
  wire[3:0] FpAlu_8U_23U_mux1h_1037_nl;
  wire[0:0] FpAlu_8U_23U_and_615_nl;
  wire[0:0] FpAlu_8U_23U_and_616_nl;
  wire[0:0] FpAlu_8U_23U_and_617_nl;
  wire[0:0] FpAlu_8U_23U_not_115_nl;
  wire[0:0] and_4122_nl;
  wire[0:0] mux_1572_nl;
  wire[0:0] or_5097_nl;
  wire[0:0] nand_429_nl;
  wire[3:0] FpAlu_8U_23U_FpAlu_8U_23U_nor_15_nl;
  wire[3:0] FpAlu_8U_23U_nor_15_nl;
  wire[3:0] FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_14_nl;
  wire[0:0] and_4119_nl;
  wire[21:0] FpAlu_8U_23U_and_11_nl;
  wire[21:0] FpAlu_8U_23U_mux1h_1033_nl;
  wire[0:0] FpAlu_8U_23U_not_84_nl;
  wire[3:0] FpAlu_8U_23U_and_10_nl;
  wire[3:0] FpAlu_8U_23U_mux1h_1034_nl;
  wire[0:0] FpAlu_8U_23U_and_620_nl;
  wire[0:0] FpAlu_8U_23U_and_621_nl;
  wire[0:0] FpAlu_8U_23U_and_622_nl;
  wire[0:0] FpAlu_8U_23U_not_116_nl;
  wire[0:0] and_4116_nl;
  wire[0:0] mux_1575_nl;
  wire[0:0] or_5103_nl;
  wire[0:0] nand_430_nl;
  wire[3:0] FpAlu_8U_23U_FpAlu_8U_23U_nor_14_nl;
  wire[3:0] FpAlu_8U_23U_nor_14_nl;
  wire[3:0] FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_13_nl;
  wire[0:0] and_4113_nl;
  wire[21:0] FpAlu_8U_23U_and_15_nl;
  wire[21:0] FpAlu_8U_23U_mux1h_1030_nl;
  wire[0:0] FpAlu_8U_23U_not_86_nl;
  wire[3:0] FpAlu_8U_23U_and_14_nl;
  wire[3:0] FpAlu_8U_23U_mux1h_1031_nl;
  wire[0:0] FpAlu_8U_23U_and_625_nl;
  wire[0:0] FpAlu_8U_23U_and_626_nl;
  wire[0:0] FpAlu_8U_23U_and_627_nl;
  wire[0:0] FpAlu_8U_23U_not_117_nl;
  wire[0:0] and_4110_nl;
  wire[0:0] mux_1578_nl;
  wire[0:0] or_5109_nl;
  wire[0:0] nand_431_nl;
  wire[3:0] FpAlu_8U_23U_FpAlu_8U_23U_nor_13_nl;
  wire[3:0] FpAlu_8U_23U_nor_13_nl;
  wire[3:0] FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_12_nl;
  wire[0:0] and_4107_nl;
  wire[21:0] FpAlu_8U_23U_and_19_nl;
  wire[21:0] FpAlu_8U_23U_mux1h_1027_nl;
  wire[0:0] FpAlu_8U_23U_not_88_nl;
  wire[3:0] FpAlu_8U_23U_and_18_nl;
  wire[3:0] FpAlu_8U_23U_mux1h_1028_nl;
  wire[0:0] FpAlu_8U_23U_and_630_nl;
  wire[0:0] FpAlu_8U_23U_and_631_nl;
  wire[0:0] FpAlu_8U_23U_and_632_nl;
  wire[0:0] FpAlu_8U_23U_not_118_nl;
  wire[0:0] and_4104_nl;
  wire[0:0] mux_1581_nl;
  wire[0:0] or_5115_nl;
  wire[0:0] nand_432_nl;
  wire[3:0] FpAlu_8U_23U_FpAlu_8U_23U_nor_12_nl;
  wire[3:0] FpAlu_8U_23U_nor_12_nl;
  wire[3:0] FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_11_nl;
  wire[0:0] and_4101_nl;
  wire[21:0] FpAlu_8U_23U_and_23_nl;
  wire[21:0] FpAlu_8U_23U_mux1h_292_nl;
  wire[0:0] FpAlu_8U_23U_not_90_nl;
  wire[3:0] FpAlu_8U_23U_and_22_nl;
  wire[3:0] FpAlu_8U_23U_mux1h_1025_nl;
  wire[0:0] FpAlu_8U_23U_and_635_nl;
  wire[0:0] FpAlu_8U_23U_and_636_nl;
  wire[0:0] FpAlu_8U_23U_and_637_nl;
  wire[0:0] FpAlu_8U_23U_not_119_nl;
  wire[0:0] and_4098_nl;
  wire[0:0] mux_1584_nl;
  wire[0:0] or_5121_nl;
  wire[0:0] nand_433_nl;
  wire[3:0] FpAlu_8U_23U_FpAlu_8U_23U_nor_11_nl;
  wire[3:0] FpAlu_8U_23U_nor_11_nl;
  wire[3:0] FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_10_nl;
  wire[0:0] and_4095_nl;
  wire[21:0] FpAlu_8U_23U_and_27_nl;
  wire[21:0] FpAlu_8U_23U_mux1h_344_nl;
  wire[0:0] FpAlu_8U_23U_not_92_nl;
  wire[3:0] FpAlu_8U_23U_and_26_nl;
  wire[3:0] FpAlu_8U_23U_mux1h_1023_nl;
  wire[0:0] FpAlu_8U_23U_and_640_nl;
  wire[0:0] FpAlu_8U_23U_and_641_nl;
  wire[0:0] FpAlu_8U_23U_and_642_nl;
  wire[0:0] FpAlu_8U_23U_not_120_nl;
  wire[0:0] and_4092_nl;
  wire[0:0] mux_1587_nl;
  wire[0:0] or_5127_nl;
  wire[0:0] nand_434_nl;
  wire[3:0] FpAlu_8U_23U_FpAlu_8U_23U_nor_10_nl;
  wire[3:0] FpAlu_8U_23U_nor_10_nl;
  wire[3:0] FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_9_nl;
  wire[0:0] and_4089_nl;
  wire[21:0] FpAlu_8U_23U_and_31_nl;
  wire[21:0] FpAlu_8U_23U_mux1h_396_nl;
  wire[0:0] FpAlu_8U_23U_not_94_nl;
  wire[3:0] FpAlu_8U_23U_and_30_nl;
  wire[3:0] FpAlu_8U_23U_mux1h_1021_nl;
  wire[0:0] FpAlu_8U_23U_and_645_nl;
  wire[0:0] FpAlu_8U_23U_and_646_nl;
  wire[0:0] FpAlu_8U_23U_and_647_nl;
  wire[0:0] FpAlu_8U_23U_not_121_nl;
  wire[0:0] and_4086_nl;
  wire[0:0] mux_1590_nl;
  wire[0:0] or_5133_nl;
  wire[0:0] nand_435_nl;
  wire[3:0] FpAlu_8U_23U_FpAlu_8U_23U_nor_9_nl;
  wire[3:0] FpAlu_8U_23U_nor_9_nl;
  wire[3:0] FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_8_nl;
  wire[0:0] and_4083_nl;
  wire[21:0] FpAlu_8U_23U_and_35_nl;
  wire[21:0] FpAlu_8U_23U_mux1h_448_nl;
  wire[0:0] FpAlu_8U_23U_not_96_nl;
  wire[3:0] FpAlu_8U_23U_and_34_nl;
  wire[3:0] FpAlu_8U_23U_mux1h_1019_nl;
  wire[0:0] FpAlu_8U_23U_and_650_nl;
  wire[0:0] FpAlu_8U_23U_and_651_nl;
  wire[0:0] FpAlu_8U_23U_and_652_nl;
  wire[0:0] FpAlu_8U_23U_not_122_nl;
  wire[0:0] and_4080_nl;
  wire[0:0] mux_1593_nl;
  wire[0:0] or_5139_nl;
  wire[0:0] nand_436_nl;
  wire[3:0] FpAlu_8U_23U_FpAlu_8U_23U_nor_8_nl;
  wire[3:0] FpAlu_8U_23U_nor_8_nl;
  wire[3:0] FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_7_nl;
  wire[0:0] and_4077_nl;
  wire[21:0] FpAlu_8U_23U_and_39_nl;
  wire[21:0] FpAlu_8U_23U_mux1h_500_nl;
  wire[0:0] FpAlu_8U_23U_not_98_nl;
  wire[3:0] FpAlu_8U_23U_and_38_nl;
  wire[3:0] FpAlu_8U_23U_mux1h_1017_nl;
  wire[0:0] FpAlu_8U_23U_and_655_nl;
  wire[0:0] FpAlu_8U_23U_and_656_nl;
  wire[0:0] FpAlu_8U_23U_and_657_nl;
  wire[0:0] FpAlu_8U_23U_not_123_nl;
  wire[0:0] and_4074_nl;
  wire[0:0] mux_1596_nl;
  wire[0:0] or_5145_nl;
  wire[0:0] nand_437_nl;
  wire[3:0] FpAlu_8U_23U_FpAlu_8U_23U_nor_7_nl;
  wire[3:0] FpAlu_8U_23U_nor_7_nl;
  wire[3:0] FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_6_nl;
  wire[0:0] and_4071_nl;
  wire[21:0] FpAlu_8U_23U_and_43_nl;
  wire[21:0] FpAlu_8U_23U_mux1h_552_nl;
  wire[0:0] FpAlu_8U_23U_not_100_nl;
  wire[3:0] FpAlu_8U_23U_and_42_nl;
  wire[3:0] FpAlu_8U_23U_mux1h_1015_nl;
  wire[0:0] FpAlu_8U_23U_and_660_nl;
  wire[0:0] FpAlu_8U_23U_and_661_nl;
  wire[0:0] FpAlu_8U_23U_and_662_nl;
  wire[0:0] FpAlu_8U_23U_not_124_nl;
  wire[0:0] and_4068_nl;
  wire[0:0] mux_1599_nl;
  wire[0:0] or_5151_nl;
  wire[0:0] nand_438_nl;
  wire[3:0] FpAlu_8U_23U_FpAlu_8U_23U_nor_6_nl;
  wire[3:0] FpAlu_8U_23U_nor_6_nl;
  wire[3:0] FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_5_nl;
  wire[0:0] and_4065_nl;
  wire[21:0] FpAlu_8U_23U_and_47_nl;
  wire[21:0] FpAlu_8U_23U_mux1h_604_nl;
  wire[0:0] FpAlu_8U_23U_not_102_nl;
  wire[3:0] FpAlu_8U_23U_and_46_nl;
  wire[3:0] FpAlu_8U_23U_mux1h_1013_nl;
  wire[0:0] FpAlu_8U_23U_and_665_nl;
  wire[0:0] FpAlu_8U_23U_and_666_nl;
  wire[0:0] FpAlu_8U_23U_and_667_nl;
  wire[0:0] FpAlu_8U_23U_not_125_nl;
  wire[0:0] and_4062_nl;
  wire[0:0] mux_1602_nl;
  wire[0:0] or_5157_nl;
  wire[0:0] nand_439_nl;
  wire[3:0] FpAlu_8U_23U_FpAlu_8U_23U_nor_5_nl;
  wire[3:0] FpAlu_8U_23U_nor_5_nl;
  wire[3:0] FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_4_nl;
  wire[0:0] and_4059_nl;
  wire[21:0] FpAlu_8U_23U_and_51_nl;
  wire[21:0] FpAlu_8U_23U_mux1h_656_nl;
  wire[0:0] FpAlu_8U_23U_not_104_nl;
  wire[3:0] FpAlu_8U_23U_and_50_nl;
  wire[3:0] FpAlu_8U_23U_mux1h_1011_nl;
  wire[0:0] FpAlu_8U_23U_and_670_nl;
  wire[0:0] FpAlu_8U_23U_and_671_nl;
  wire[0:0] FpAlu_8U_23U_and_672_nl;
  wire[0:0] FpAlu_8U_23U_not_126_nl;
  wire[0:0] and_4056_nl;
  wire[0:0] mux_1605_nl;
  wire[0:0] or_5163_nl;
  wire[0:0] nand_440_nl;
  wire[3:0] FpAlu_8U_23U_FpAlu_8U_23U_nor_4_nl;
  wire[3:0] FpAlu_8U_23U_nor_4_nl;
  wire[3:0] FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_3_nl;
  wire[0:0] and_4053_nl;
  wire[21:0] FpAlu_8U_23U_and_55_nl;
  wire[21:0] FpAlu_8U_23U_mux1h_708_nl;
  wire[0:0] FpAlu_8U_23U_not_106_nl;
  wire[3:0] FpAlu_8U_23U_and_54_nl;
  wire[3:0] FpAlu_8U_23U_mux1h_1009_nl;
  wire[0:0] FpAlu_8U_23U_and_675_nl;
  wire[0:0] FpAlu_8U_23U_and_676_nl;
  wire[0:0] FpAlu_8U_23U_and_677_nl;
  wire[0:0] FpAlu_8U_23U_not_127_nl;
  wire[0:0] and_4050_nl;
  wire[0:0] mux_1608_nl;
  wire[0:0] or_5169_nl;
  wire[0:0] nand_441_nl;
  wire[3:0] FpAlu_8U_23U_FpAlu_8U_23U_nor_3_nl;
  wire[3:0] FpAlu_8U_23U_nor_3_nl;
  wire[3:0] FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_2_nl;
  wire[0:0] and_4047_nl;
  wire[21:0] FpAlu_8U_23U_and_59_nl;
  wire[21:0] FpAlu_8U_23U_mux1h_760_nl;
  wire[0:0] FpAlu_8U_23U_not_108_nl;
  wire[3:0] FpAlu_8U_23U_and_58_nl;
  wire[3:0] FpAlu_8U_23U_mux1h_1007_nl;
  wire[0:0] FpAlu_8U_23U_and_680_nl;
  wire[0:0] FpAlu_8U_23U_and_681_nl;
  wire[0:0] FpAlu_8U_23U_and_682_nl;
  wire[0:0] FpAlu_8U_23U_not_128_nl;
  wire[0:0] and_4044_nl;
  wire[0:0] mux_1611_nl;
  wire[0:0] or_5175_nl;
  wire[0:0] nand_442_nl;
  wire[3:0] FpAlu_8U_23U_FpAlu_8U_23U_nor_2_nl;
  wire[3:0] FpAlu_8U_23U_nor_2_nl;
  wire[3:0] FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_1_nl;
  wire[0:0] and_4041_nl;
  wire[21:0] FpAlu_8U_23U_and_63_nl;
  wire[21:0] FpAlu_8U_23U_mux1h_1004_nl;
  wire[0:0] FpAlu_8U_23U_not_110_nl;
  wire[3:0] FpAlu_8U_23U_and_62_nl;
  wire[3:0] FpAlu_8U_23U_mux1h_1005_nl;
  wire[0:0] FpAlu_8U_23U_and_685_nl;
  wire[0:0] FpAlu_8U_23U_and_686_nl;
  wire[0:0] FpAlu_8U_23U_and_687_nl;
  wire[0:0] FpAlu_8U_23U_not_129_nl;
  wire[0:0] and_4038_nl;
  wire[0:0] mux_1614_nl;
  wire[0:0] or_5181_nl;
  wire[0:0] nand_443_nl;
  wire[3:0] FpAlu_8U_23U_FpAlu_8U_23U_nor_1_nl;
  wire[3:0] FpAlu_8U_23U_nor_1_nl;
  wire[3:0] FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_nl;
  wire[0:0] and_4035_nl;
  wire[0:0] and_492_nl;
  wire[0:0] mux_15_nl;
  wire[0:0] nor_2055_nl;
  wire[0:0] mux_18_nl;
  wire[0:0] nor_2052_nl;
  wire[0:0] mux_17_nl;
  wire[0:0] or_35_nl;
  wire[0:0] nor_2053_nl;
  wire[0:0] and_509_nl;
  wire[0:0] and_522_nl;
  wire[0:0] and_535_nl;
  wire[0:0] and_548_nl;
  wire[0:0] and_561_nl;
  wire[0:0] and_574_nl;
  wire[0:0] and_587_nl;
  wire[0:0] and_600_nl;
  wire[0:0] and_613_nl;
  wire[0:0] and_626_nl;
  wire[0:0] and_639_nl;
  wire[0:0] and_652_nl;
  wire[0:0] and_665_nl;
  wire[0:0] and_678_nl;
  wire[0:0] and_691_nl;
  wire[0:0] mux_159_nl;
  wire[0:0] mux_158_nl;
  wire[0:0] mux_165_nl;
  wire[0:0] mux_164_nl;
  wire[0:0] mux_172_nl;
  wire[0:0] mux_171_nl;
  wire[0:0] mux_170_nl;
  wire[0:0] or_359_nl;
  wire[0:0] or_361_nl;
  wire[0:0] nor_1931_nl;
  wire[0:0] nor_1929_nl;
  wire[0:0] nor_1867_nl;
  wire[0:0] mux_286_nl;
  wire[0:0] nor_1863_nl;
  wire[0:0] mux_349_nl;
  wire[0:0] nor_1817_nl;
  wire[0:0] mux_348_nl;
  wire[0:0] mux_351_nl;
  wire[0:0] nor_1816_nl;
  wire[0:0] mux_352_nl;
  wire[0:0] nor_1814_nl;
  wire[0:0] mux_386_nl;
  wire[0:0] mux_384_nl;
  wire[0:0] mux_383_nl;
  wire[0:0] nor_1745_nl;
  wire[0:0] nor_1750_nl;
  wire[0:0] mux_385_nl;
  wire[0:0] nor_1751_nl;
  wire[0:0] nor_1752_nl;
  wire[0:0] mux_388_nl;
  wire[0:0] mux_387_nl;
  wire[0:0] and_3766_nl;
  wire[0:0] nor_1744_nl;
  wire[0:0] mux_390_nl;
  wire[0:0] mux_389_nl;
  wire[0:0] nor_1739_nl;
  wire[0:0] nor_1740_nl;
  wire[0:0] nor_1741_nl;
  wire[0:0] mux_395_nl;
  wire[0:0] mux_394_nl;
  wire[0:0] nor_1735_nl;
  wire[0:0] nor_1736_nl;
  wire[0:0] nor_1737_nl;
  wire[0:0] mux_396_nl;
  wire[0:0] nor_1733_nl;
  wire[0:0] nor_1734_nl;
  wire[0:0] mux_397_nl;
  wire[0:0] nor_1731_nl;
  wire[0:0] nor_1732_nl;
  wire[0:0] mux_398_nl;
  wire[0:0] mux_403_nl;
  wire[0:0] mux_402_nl;
  wire[0:0] mux_401_nl;
  wire[0:0] nor_338_nl;
  wire[0:0] mux_404_nl;
  wire[0:0] nor_1726_nl;
  wire[0:0] nor_1729_nl;
  wire[0:0] mux_409_nl;
  wire[0:0] mux_406_nl;
  wire[0:0] mux_405_nl;
  wire[0:0] nor_1717_nl;
  wire[0:0] mux_408_nl;
  wire[0:0] mux_407_nl;
  wire[0:0] nor_1722_nl;
  wire[0:0] mux_411_nl;
  wire[0:0] mux_410_nl;
  wire[0:0] and_3763_nl;
  wire[0:0] nor_1716_nl;
  wire[0:0] mux_413_nl;
  wire[0:0] mux_412_nl;
  wire[0:0] nor_1711_nl;
  wire[0:0] nor_1712_nl;
  wire[0:0] nor_1713_nl;
  wire[0:0] mux_417_nl;
  wire[0:0] mux_416_nl;
  wire[0:0] nor_1708_nl;
  wire[0:0] nor_1709_nl;
  wire[0:0] nor_1710_nl;
  wire[0:0] mux_418_nl;
  wire[0:0] nor_1706_nl;
  wire[0:0] nor_1707_nl;
  wire[0:0] mux_419_nl;
  wire[0:0] nor_1704_nl;
  wire[0:0] nor_1705_nl;
  wire[0:0] mux_425_nl;
  wire[0:0] nor_1699_nl;
  wire[0:0] nor_1702_nl;
  wire[0:0] mux_430_nl;
  wire[0:0] mux_427_nl;
  wire[0:0] mux_426_nl;
  wire[0:0] nor_1690_nl;
  wire[0:0] mux_429_nl;
  wire[0:0] mux_428_nl;
  wire[0:0] nor_1695_nl;
  wire[0:0] mux_432_nl;
  wire[0:0] mux_431_nl;
  wire[0:0] and_3760_nl;
  wire[0:0] nor_1689_nl;
  wire[0:0] mux_434_nl;
  wire[0:0] mux_433_nl;
  wire[0:0] nor_1684_nl;
  wire[0:0] nor_1685_nl;
  wire[0:0] nor_1686_nl;
  wire[0:0] mux_438_nl;
  wire[0:0] mux_437_nl;
  wire[0:0] nor_1681_nl;
  wire[0:0] nor_1682_nl;
  wire[0:0] nor_1683_nl;
  wire[0:0] mux_439_nl;
  wire[0:0] nor_1679_nl;
  wire[0:0] nor_1680_nl;
  wire[0:0] mux_440_nl;
  wire[0:0] nor_1677_nl;
  wire[0:0] nor_1678_nl;
  wire[0:0] mux_446_nl;
  wire[0:0] nor_1672_nl;
  wire[0:0] nor_1675_nl;
  wire[0:0] mux_451_nl;
  wire[0:0] mux_448_nl;
  wire[0:0] mux_447_nl;
  wire[0:0] nor_1663_nl;
  wire[0:0] mux_450_nl;
  wire[0:0] mux_449_nl;
  wire[0:0] nor_1668_nl;
  wire[0:0] mux_453_nl;
  wire[0:0] mux_452_nl;
  wire[0:0] and_3757_nl;
  wire[0:0] nor_1662_nl;
  wire[0:0] mux_455_nl;
  wire[0:0] mux_454_nl;
  wire[0:0] nor_1657_nl;
  wire[0:0] nor_1658_nl;
  wire[0:0] nor_1659_nl;
  wire[0:0] mux_459_nl;
  wire[0:0] mux_458_nl;
  wire[0:0] nor_1654_nl;
  wire[0:0] nor_1655_nl;
  wire[0:0] nor_1656_nl;
  wire[0:0] mux_460_nl;
  wire[0:0] nor_1652_nl;
  wire[0:0] nor_1653_nl;
  wire[0:0] mux_461_nl;
  wire[0:0] nor_1650_nl;
  wire[0:0] nor_1651_nl;
  wire[0:0] mux_467_nl;
  wire[0:0] nor_1645_nl;
  wire[0:0] nor_1648_nl;
  wire[0:0] mux_472_nl;
  wire[0:0] mux_469_nl;
  wire[0:0] mux_468_nl;
  wire[0:0] nor_1636_nl;
  wire[0:0] mux_471_nl;
  wire[0:0] mux_470_nl;
  wire[0:0] nor_1641_nl;
  wire[0:0] mux_474_nl;
  wire[0:0] mux_473_nl;
  wire[0:0] and_3754_nl;
  wire[0:0] nor_1635_nl;
  wire[0:0] mux_476_nl;
  wire[0:0] mux_475_nl;
  wire[0:0] nor_1630_nl;
  wire[0:0] nor_1631_nl;
  wire[0:0] nor_1632_nl;
  wire[0:0] mux_480_nl;
  wire[0:0] mux_479_nl;
  wire[0:0] nor_1627_nl;
  wire[0:0] nor_1628_nl;
  wire[0:0] nor_1629_nl;
  wire[0:0] mux_481_nl;
  wire[0:0] nor_1625_nl;
  wire[0:0] nor_1626_nl;
  wire[0:0] mux_482_nl;
  wire[0:0] nor_1623_nl;
  wire[0:0] nor_1624_nl;
  wire[0:0] mux_488_nl;
  wire[0:0] nor_1618_nl;
  wire[0:0] nor_1621_nl;
  wire[0:0] mux_493_nl;
  wire[0:0] mux_490_nl;
  wire[0:0] mux_489_nl;
  wire[0:0] nor_1609_nl;
  wire[0:0] mux_492_nl;
  wire[0:0] mux_491_nl;
  wire[0:0] nor_1614_nl;
  wire[0:0] mux_495_nl;
  wire[0:0] mux_494_nl;
  wire[0:0] and_3751_nl;
  wire[0:0] nor_1608_nl;
  wire[0:0] mux_497_nl;
  wire[0:0] mux_496_nl;
  wire[0:0] nor_1603_nl;
  wire[0:0] nor_1604_nl;
  wire[0:0] nor_1605_nl;
  wire[0:0] mux_501_nl;
  wire[0:0] mux_500_nl;
  wire[0:0] nor_1600_nl;
  wire[0:0] nor_1601_nl;
  wire[0:0] nor_1602_nl;
  wire[0:0] mux_502_nl;
  wire[0:0] nor_1598_nl;
  wire[0:0] nor_1599_nl;
  wire[0:0] mux_503_nl;
  wire[0:0] nor_1596_nl;
  wire[0:0] nor_1597_nl;
  wire[0:0] mux_509_nl;
  wire[0:0] nor_1591_nl;
  wire[0:0] nor_1594_nl;
  wire[0:0] mux_514_nl;
  wire[0:0] mux_511_nl;
  wire[0:0] mux_510_nl;
  wire[0:0] nor_1582_nl;
  wire[0:0] mux_513_nl;
  wire[0:0] mux_512_nl;
  wire[0:0] nor_1587_nl;
  wire[0:0] mux_516_nl;
  wire[0:0] mux_515_nl;
  wire[0:0] and_3747_nl;
  wire[0:0] and_3748_nl;
  wire[0:0] nor_1581_nl;
  wire[0:0] mux_518_nl;
  wire[0:0] mux_517_nl;
  wire[0:0] nor_1577_nl;
  wire[0:0] nor_1578_nl;
  wire[0:0] nor_1579_nl;
  wire[0:0] mux_522_nl;
  wire[0:0] mux_521_nl;
  wire[0:0] nor_1574_nl;
  wire[0:0] nor_1575_nl;
  wire[0:0] nor_1576_nl;
  wire[0:0] mux_523_nl;
  wire[0:0] nor_1572_nl;
  wire[0:0] nor_1573_nl;
  wire[0:0] mux_524_nl;
  wire[0:0] nor_1570_nl;
  wire[0:0] nor_1571_nl;
  wire[0:0] mux_530_nl;
  wire[0:0] nor_1565_nl;
  wire[0:0] nor_1568_nl;
  wire[0:0] mux_535_nl;
  wire[0:0] mux_532_nl;
  wire[0:0] mux_531_nl;
  wire[0:0] nor_1556_nl;
  wire[0:0] mux_534_nl;
  wire[0:0] mux_533_nl;
  wire[0:0] nor_1561_nl;
  wire[0:0] mux_537_nl;
  wire[0:0] mux_536_nl;
  wire[0:0] and_3743_nl;
  wire[0:0] and_3744_nl;
  wire[0:0] nor_1555_nl;
  wire[0:0] mux_539_nl;
  wire[0:0] mux_538_nl;
  wire[0:0] nor_1551_nl;
  wire[0:0] nor_1552_nl;
  wire[0:0] nor_1553_nl;
  wire[0:0] mux_543_nl;
  wire[0:0] mux_542_nl;
  wire[0:0] nor_1548_nl;
  wire[0:0] nor_1549_nl;
  wire[0:0] nor_1550_nl;
  wire[0:0] mux_544_nl;
  wire[0:0] nor_1546_nl;
  wire[0:0] nor_1547_nl;
  wire[0:0] mux_545_nl;
  wire[0:0] nor_1544_nl;
  wire[0:0] nor_1545_nl;
  wire[0:0] mux_551_nl;
  wire[0:0] nor_1539_nl;
  wire[0:0] nor_1542_nl;
  wire[0:0] mux_556_nl;
  wire[0:0] mux_553_nl;
  wire[0:0] mux_552_nl;
  wire[0:0] nor_1530_nl;
  wire[0:0] mux_555_nl;
  wire[0:0] mux_554_nl;
  wire[0:0] nor_1535_nl;
  wire[0:0] mux_558_nl;
  wire[0:0] mux_557_nl;
  wire[0:0] and_3739_nl;
  wire[0:0] and_3740_nl;
  wire[0:0] nor_1529_nl;
  wire[0:0] mux_560_nl;
  wire[0:0] mux_559_nl;
  wire[0:0] nor_1525_nl;
  wire[0:0] nor_1526_nl;
  wire[0:0] nor_1527_nl;
  wire[0:0] mux_564_nl;
  wire[0:0] mux_563_nl;
  wire[0:0] nor_1522_nl;
  wire[0:0] nor_1523_nl;
  wire[0:0] nor_1524_nl;
  wire[0:0] mux_565_nl;
  wire[0:0] nor_1520_nl;
  wire[0:0] nor_1521_nl;
  wire[0:0] mux_566_nl;
  wire[0:0] nor_1518_nl;
  wire[0:0] nor_1519_nl;
  wire[0:0] mux_572_nl;
  wire[0:0] nor_1513_nl;
  wire[0:0] nor_1516_nl;
  wire[0:0] mux_577_nl;
  wire[0:0] mux_574_nl;
  wire[0:0] mux_573_nl;
  wire[0:0] nor_1504_nl;
  wire[0:0] mux_576_nl;
  wire[0:0] mux_575_nl;
  wire[0:0] nor_1509_nl;
  wire[0:0] mux_579_nl;
  wire[0:0] mux_578_nl;
  wire[0:0] and_3735_nl;
  wire[0:0] and_3736_nl;
  wire[0:0] nor_1503_nl;
  wire[0:0] mux_581_nl;
  wire[0:0] mux_580_nl;
  wire[0:0] nor_1499_nl;
  wire[0:0] nor_1500_nl;
  wire[0:0] nor_1501_nl;
  wire[0:0] mux_585_nl;
  wire[0:0] mux_584_nl;
  wire[0:0] nor_1496_nl;
  wire[0:0] nor_1497_nl;
  wire[0:0] nor_1498_nl;
  wire[0:0] mux_586_nl;
  wire[0:0] nor_1494_nl;
  wire[0:0] nor_1495_nl;
  wire[0:0] mux_587_nl;
  wire[0:0] nor_1492_nl;
  wire[0:0] nor_1493_nl;
  wire[0:0] mux_593_nl;
  wire[0:0] nor_1487_nl;
  wire[0:0] nor_1490_nl;
  wire[0:0] mux_598_nl;
  wire[0:0] mux_595_nl;
  wire[0:0] mux_594_nl;
  wire[0:0] nor_1478_nl;
  wire[0:0] mux_597_nl;
  wire[0:0] mux_596_nl;
  wire[0:0] nor_1483_nl;
  wire[0:0] mux_600_nl;
  wire[0:0] mux_599_nl;
  wire[0:0] and_3731_nl;
  wire[0:0] and_3732_nl;
  wire[0:0] nor_1477_nl;
  wire[0:0] mux_602_nl;
  wire[0:0] mux_601_nl;
  wire[0:0] nor_1473_nl;
  wire[0:0] nor_1474_nl;
  wire[0:0] nor_1475_nl;
  wire[0:0] mux_606_nl;
  wire[0:0] mux_605_nl;
  wire[0:0] nor_1470_nl;
  wire[0:0] nor_1471_nl;
  wire[0:0] nor_1472_nl;
  wire[0:0] mux_607_nl;
  wire[0:0] nor_1468_nl;
  wire[0:0] nor_1469_nl;
  wire[0:0] mux_608_nl;
  wire[0:0] nor_1466_nl;
  wire[0:0] nor_1467_nl;
  wire[0:0] mux_614_nl;
  wire[0:0] nor_1461_nl;
  wire[0:0] nor_1464_nl;
  wire[0:0] mux_619_nl;
  wire[0:0] mux_616_nl;
  wire[0:0] mux_615_nl;
  wire[0:0] nor_1452_nl;
  wire[0:0] mux_618_nl;
  wire[0:0] mux_617_nl;
  wire[0:0] nor_1457_nl;
  wire[0:0] mux_621_nl;
  wire[0:0] mux_620_nl;
  wire[0:0] and_3727_nl;
  wire[0:0] and_3728_nl;
  wire[0:0] nor_1451_nl;
  wire[0:0] mux_623_nl;
  wire[0:0] mux_622_nl;
  wire[0:0] nor_1447_nl;
  wire[0:0] nor_1448_nl;
  wire[0:0] nor_1449_nl;
  wire[0:0] mux_627_nl;
  wire[0:0] mux_626_nl;
  wire[0:0] nor_1444_nl;
  wire[0:0] nor_1445_nl;
  wire[0:0] nor_1446_nl;
  wire[0:0] mux_628_nl;
  wire[0:0] nor_1442_nl;
  wire[0:0] nor_1443_nl;
  wire[0:0] mux_629_nl;
  wire[0:0] nor_1440_nl;
  wire[0:0] nor_1441_nl;
  wire[0:0] mux_635_nl;
  wire[0:0] nor_1435_nl;
  wire[0:0] nor_1438_nl;
  wire[0:0] mux_640_nl;
  wire[0:0] mux_637_nl;
  wire[0:0] mux_636_nl;
  wire[0:0] nor_1426_nl;
  wire[0:0] mux_639_nl;
  wire[0:0] mux_638_nl;
  wire[0:0] nor_1431_nl;
  wire[0:0] mux_642_nl;
  wire[0:0] mux_641_nl;
  wire[0:0] and_3723_nl;
  wire[0:0] and_3724_nl;
  wire[0:0] nor_1425_nl;
  wire[0:0] mux_644_nl;
  wire[0:0] mux_643_nl;
  wire[0:0] nor_1421_nl;
  wire[0:0] nor_1422_nl;
  wire[0:0] nor_1423_nl;
  wire[0:0] mux_648_nl;
  wire[0:0] mux_647_nl;
  wire[0:0] nor_1418_nl;
  wire[0:0] nor_1419_nl;
  wire[0:0] nor_1420_nl;
  wire[0:0] mux_649_nl;
  wire[0:0] nor_1416_nl;
  wire[0:0] nor_1417_nl;
  wire[0:0] mux_650_nl;
  wire[0:0] nor_1414_nl;
  wire[0:0] nor_1415_nl;
  wire[0:0] mux_656_nl;
  wire[0:0] nor_1409_nl;
  wire[0:0] nor_1412_nl;
  wire[0:0] mux_661_nl;
  wire[0:0] mux_658_nl;
  wire[0:0] mux_657_nl;
  wire[0:0] nor_1400_nl;
  wire[0:0] mux_660_nl;
  wire[0:0] mux_659_nl;
  wire[0:0] nor_1405_nl;
  wire[0:0] mux_663_nl;
  wire[0:0] mux_662_nl;
  wire[0:0] and_3719_nl;
  wire[0:0] and_3720_nl;
  wire[0:0] nor_1399_nl;
  wire[0:0] mux_665_nl;
  wire[0:0] mux_664_nl;
  wire[0:0] nor_1395_nl;
  wire[0:0] nor_1396_nl;
  wire[0:0] nor_1397_nl;
  wire[0:0] mux_669_nl;
  wire[0:0] mux_668_nl;
  wire[0:0] nor_1392_nl;
  wire[0:0] nor_1393_nl;
  wire[0:0] nor_1394_nl;
  wire[0:0] mux_670_nl;
  wire[0:0] nor_1390_nl;
  wire[0:0] nor_1391_nl;
  wire[0:0] mux_671_nl;
  wire[0:0] nor_1388_nl;
  wire[0:0] nor_1389_nl;
  wire[0:0] mux_677_nl;
  wire[0:0] nor_1383_nl;
  wire[0:0] nor_1386_nl;
  wire[0:0] mux_681_nl;
  wire[0:0] mux_679_nl;
  wire[0:0] mux_678_nl;
  wire[0:0] nor_1375_nl;
  wire[0:0] nor_1380_nl;
  wire[0:0] mux_680_nl;
  wire[0:0] nor_1381_nl;
  wire[0:0] nor_1382_nl;
  wire[0:0] mux_683_nl;
  wire[0:0] mux_682_nl;
  wire[0:0] and_3715_nl;
  wire[0:0] and_3716_nl;
  wire[0:0] nor_1374_nl;
  wire[0:0] mux_685_nl;
  wire[0:0] mux_684_nl;
  wire[0:0] nor_1370_nl;
  wire[0:0] nor_1371_nl;
  wire[0:0] nor_1372_nl;
  wire[0:0] mux_689_nl;
  wire[0:0] mux_688_nl;
  wire[0:0] nor_1367_nl;
  wire[0:0] nor_1368_nl;
  wire[0:0] nor_1369_nl;
  wire[0:0] mux_690_nl;
  wire[0:0] nor_1365_nl;
  wire[0:0] nor_1366_nl;
  wire[0:0] mux_691_nl;
  wire[0:0] nor_1363_nl;
  wire[0:0] nor_1364_nl;
  wire[0:0] mux_697_nl;
  wire[0:0] nor_1358_nl;
  wire[0:0] nor_1361_nl;
  wire[0:0] mux_701_nl;
  wire[0:0] mux_699_nl;
  wire[0:0] mux_698_nl;
  wire[0:0] nor_1350_nl;
  wire[0:0] nor_1355_nl;
  wire[0:0] mux_700_nl;
  wire[0:0] nor_1356_nl;
  wire[0:0] nor_1357_nl;
  wire[0:0] mux_703_nl;
  wire[0:0] mux_702_nl;
  wire[0:0] and_3711_nl;
  wire[0:0] and_3712_nl;
  wire[0:0] nor_1349_nl;
  wire[0:0] mux_705_nl;
  wire[0:0] mux_704_nl;
  wire[0:0] nor_1345_nl;
  wire[0:0] nor_1346_nl;
  wire[0:0] nor_1347_nl;
  wire[0:0] mux_709_nl;
  wire[0:0] mux_708_nl;
  wire[0:0] nor_1342_nl;
  wire[0:0] nor_1343_nl;
  wire[0:0] nor_1344_nl;
  wire[0:0] mux_710_nl;
  wire[0:0] nor_1340_nl;
  wire[0:0] nor_1341_nl;
  wire[0:0] mux_711_nl;
  wire[0:0] nor_1338_nl;
  wire[0:0] nor_1339_nl;
  wire[0:0] mux_717_nl;
  wire[0:0] nor_1333_nl;
  wire[0:0] nor_1336_nl;
  wire[0:0] mux_719_nl;
  wire[0:0] or_1811_nl;
  wire[0:0] mux_718_nl;
  wire[0:0] or_1812_nl;
  wire[0:0] mux_729_nl;
  wire[0:0] or_1825_nl;
  wire[0:0] mux_728_nl;
  wire[0:0] mux_347_nl;
  wire[0:0] mux_751_nl;
  wire[0:0] mux_750_nl;
  wire[0:0] or_1861_nl;
  wire[0:0] or_1922_nl;
  wire[0:0] mux_804_nl;
  wire[0:0] or_1927_nl;
  wire[0:0] or_1931_nl;
  wire[0:0] nand_448_nl;
  wire[0:0] or_1937_nl;
  wire[0:0] mux_813_nl;
  wire[0:0] mux_809_nl;
  wire[0:0] mux_808_nl;
  wire[0:0] mux_806_nl;
  wire[0:0] or_1929_nl;
  wire[0:0] mux_812_nl;
  wire[0:0] or_1936_nl;
  wire[0:0] mux_810_nl;
  wire[0:0] or_1934_nl;
  wire[0:0] mux_816_nl;
  wire[0:0] mux_815_nl;
  wire[0:0] nor_1315_nl;
  wire[0:0] mux_814_nl;
  wire[0:0] nor_1316_nl;
  wire[0:0] nor_1318_nl;
  wire[0:0] mux_817_nl;
  wire[0:0] nor_1305_nl;
  wire[0:0] nor_1306_nl;
  wire[0:0] nor_1307_nl;
  wire[0:0] nor_1309_nl;
  wire[0:0] and_4250_nl;
  wire[0:0] mux_825_nl;
  wire[0:0] mux_821_nl;
  wire[0:0] mux_820_nl;
  wire[0:0] nor_1308_nl;
  wire[0:0] mux_824_nl;
  wire[0:0] mux_822_nl;
  wire[0:0] nor_1311_nl;
  wire[0:0] mux_857_nl;
  wire[0:0] mux_853_nl;
  wire[0:0] mux_852_nl;
  wire[0:0] nor_1271_nl;
  wire[0:0] mux_856_nl;
  wire[0:0] nor_1274_nl;
  wire[0:0] mux_854_nl;
  wire[0:0] or_2030_nl;
  wire[0:0] mux_870_nl;
  wire[0:0] mux_866_nl;
  wire[0:0] mux_865_nl;
  wire[0:0] mux_863_nl;
  wire[0:0] or_2051_nl;
  wire[0:0] mux_869_nl;
  wire[0:0] or_2058_nl;
  wire[0:0] mux_867_nl;
  wire[0:0] or_2056_nl;
  wire[0:0] mux_892_nl;
  wire[0:0] mux_888_nl;
  wire[0:0] mux_887_nl;
  wire[0:0] mux_885_nl;
  wire[0:0] nor_1239_nl;
  wire[0:0] nor_1240_nl;
  wire[0:0] mux_886_nl;
  wire[0:0] nor_1241_nl;
  wire[0:0] nor_1243_nl;
  wire[0:0] mux_891_nl;
  wire[0:0] mux_889_nl;
  wire[0:0] nor_1244_nl;
  wire[0:0] mux_908_nl;
  wire[0:0] mux_904_nl;
  wire[0:0] mux_903_nl;
  wire[0:0] mux_901_nl;
  wire[0:0] or_2132_nl;
  wire[0:0] mux_907_nl;
  wire[0:0] or_2137_nl;
  wire[0:0] mux_906_nl;
  wire[0:0] mux_905_nl;
  wire[0:0] or_2138_nl;
  wire[0:0] mux_912_nl;
  wire[0:0] nor_1222_nl;
  wire[0:0] mux_930_nl;
  wire[0:0] and_3670_nl;
  wire[0:0] nor_1172_nl;
  wire[0:0] mux_976_nl;
  wire[0:0] nor_1173_nl;
  wire[0:0] mux_1042_nl;
  wire[0:0] nor_1122_nl;
  wire[0:0] nor_1123_nl;
  wire[0:0] nor_1087_nl;
  wire[0:0] mux_1079_nl;
  wire[0:0] mux_1077_nl;
  wire[0:0] mux_1076_nl;
  wire[0:0] mux_1078_nl;
  wire[0:0] or_2484_nl;
  wire[0:0] nor_1088_nl;
  wire[0:0] nor_1089_nl;
  wire[0:0] mux_1081_nl;
  wire[0:0] or_2487_nl;
  wire[0:0] nor_1090_nl;
  wire[0:0] and_3622_nl;
  wire[0:0] mux_1088_nl;
  wire[0:0] nor_1084_nl;
  wire[0:0] mux_1087_nl;
  wire[0:0] mux_1086_nl;
  wire[0:0] nor_1085_nl;
  wire[0:0] mux_1085_nl;
  wire[0:0] and_4266_nl;
  wire[0:0] mux_1091_nl;
  wire[0:0] mux_1090_nl;
  wire[0:0] IsNaN_8U_23U_3_aelse_or_nl;
  wire[0:0] or_2817_nl;
  wire[0:0] mux_1348_nl;
  wire[0:0] mux_1353_nl;
  wire[0:0] or_2819_nl;
  wire[0:0] mux_1352_nl;
  wire[0:0] mux_1359_nl;
  wire[0:0] mux_1358_nl;
  wire[0:0] nor_931_nl;
  wire[0:0] or_2821_nl;
  wire[0:0] mux_1391_nl;
  wire[0:0] mux_1390_nl;
  wire[0:0] nor_920_nl;
  wire[0:0] mux_1423_nl;
  wire[0:0] mux_1422_nl;
  wire[0:0] nor_2190_nl;
  wire[0:0] nand_444_nl;
  wire[0:0] nand_445_nl;
  wire[0:0] and_1917_nl;
  wire[0:0] or_2856_nl;
  wire[0:0] mux_1458_nl;
  wire[0:0] mux_1457_nl;
  wire[0:0] or_2858_nl;
  wire[0:0] mux_1503_nl;
  wire[0:0] mux_1502_nl;
  wire[0:0] or_2905_nl;
  wire[0:0] or_2903_nl;
  wire[0:0] and_469_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_144_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_2_nl;
  wire[3:0] alu_loop_op_1_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl;
  wire[4:0] nl_alu_loop_op_1_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl;
  wire[0:0] IsZero_5U_23U_aelse_IsZero_5U_23U_or_15_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_146_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_6_nl;
  wire[3:0] alu_loop_op_2_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl;
  wire[4:0] nl_alu_loop_op_2_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl;
  wire[0:0] IsZero_5U_23U_aelse_IsZero_5U_23U_or_14_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_1_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_148_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_10_nl;
  wire[3:0] alu_loop_op_3_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl;
  wire[4:0] nl_alu_loop_op_3_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl;
  wire[0:0] IsZero_5U_23U_aelse_IsZero_5U_23U_or_13_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_2_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_150_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_14_nl;
  wire[3:0] alu_loop_op_4_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl;
  wire[4:0] nl_alu_loop_op_4_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl;
  wire[0:0] IsZero_5U_23U_aelse_IsZero_5U_23U_or_12_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_3_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_152_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_18_nl;
  wire[3:0] alu_loop_op_5_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl;
  wire[4:0] nl_alu_loop_op_5_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl;
  wire[0:0] IsZero_5U_23U_aelse_IsZero_5U_23U_or_11_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_4_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_154_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_22_nl;
  wire[3:0] alu_loop_op_6_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl;
  wire[4:0] nl_alu_loop_op_6_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl;
  wire[0:0] IsZero_5U_23U_aelse_IsZero_5U_23U_or_10_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_5_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_156_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_26_nl;
  wire[3:0] alu_loop_op_7_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl;
  wire[4:0] nl_alu_loop_op_7_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl;
  wire[0:0] IsZero_5U_23U_aelse_IsZero_5U_23U_or_9_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_6_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_158_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_30_nl;
  wire[3:0] alu_loop_op_8_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl;
  wire[4:0] nl_alu_loop_op_8_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl;
  wire[0:0] IsZero_5U_23U_aelse_IsZero_5U_23U_or_8_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_7_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_160_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_34_nl;
  wire[3:0] alu_loop_op_9_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl;
  wire[4:0] nl_alu_loop_op_9_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl;
  wire[0:0] IsZero_5U_23U_aelse_IsZero_5U_23U_or_7_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_8_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_162_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_38_nl;
  wire[3:0] alu_loop_op_10_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl;
  wire[4:0] nl_alu_loop_op_10_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl;
  wire[0:0] IsZero_5U_23U_aelse_IsZero_5U_23U_or_6_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_9_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_164_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_42_nl;
  wire[3:0] alu_loop_op_11_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl;
  wire[4:0] nl_alu_loop_op_11_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl;
  wire[0:0] IsZero_5U_23U_aelse_IsZero_5U_23U_or_5_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_10_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_166_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_46_nl;
  wire[3:0] alu_loop_op_12_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl;
  wire[4:0] nl_alu_loop_op_12_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl;
  wire[0:0] IsZero_5U_23U_aelse_IsZero_5U_23U_or_4_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_11_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_168_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_50_nl;
  wire[3:0] alu_loop_op_13_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl;
  wire[4:0] nl_alu_loop_op_13_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl;
  wire[0:0] IsZero_5U_23U_aelse_IsZero_5U_23U_or_3_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_12_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_170_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_54_nl;
  wire[3:0] alu_loop_op_14_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl;
  wire[4:0] nl_alu_loop_op_14_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl;
  wire[0:0] IsZero_5U_23U_aelse_IsZero_5U_23U_or_2_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_13_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_172_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_58_nl;
  wire[3:0] alu_loop_op_15_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl;
  wire[4:0] nl_alu_loop_op_15_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl;
  wire[0:0] IsZero_5U_23U_aelse_IsZero_5U_23U_or_1_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_14_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_174_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_62_nl;
  wire[3:0] alu_loop_op_16_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl;
  wire[4:0] nl_alu_loop_op_16_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl;
  wire[0:0] IsZero_5U_23U_aelse_IsZero_5U_23U_or_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_15_nl;
  wire[7:0] alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[8:0] nl_alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[7:0] alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_2_nl;
  wire[8:0] nl_alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_2_nl;
  wire[7:0] alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[8:0] nl_alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[7:0] alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_2_nl;
  wire[8:0] nl_alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_2_nl;
  wire[7:0] alu_loop_op_5_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[8:0] nl_alu_loop_op_5_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[7:0] alu_loop_op_6_FpAdd_8U_23U_if_3_if_acc_2_nl;
  wire[8:0] nl_alu_loop_op_6_FpAdd_8U_23U_if_3_if_acc_2_nl;
  wire[7:0] alu_loop_op_7_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[8:0] nl_alu_loop_op_7_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[7:0] alu_loop_op_8_FpAdd_8U_23U_if_3_if_acc_2_nl;
  wire[8:0] nl_alu_loop_op_8_FpAdd_8U_23U_if_3_if_acc_2_nl;
  wire[7:0] alu_loop_op_9_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[8:0] nl_alu_loop_op_9_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[7:0] alu_loop_op_10_FpAdd_8U_23U_if_3_if_acc_2_nl;
  wire[8:0] nl_alu_loop_op_10_FpAdd_8U_23U_if_3_if_acc_2_nl;
  wire[7:0] alu_loop_op_11_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[8:0] nl_alu_loop_op_11_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[7:0] alu_loop_op_12_FpAdd_8U_23U_if_3_if_acc_2_nl;
  wire[8:0] nl_alu_loop_op_12_FpAdd_8U_23U_if_3_if_acc_2_nl;
  wire[7:0] alu_loop_op_13_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[8:0] nl_alu_loop_op_13_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[7:0] alu_loop_op_14_FpAdd_8U_23U_if_3_if_acc_2_nl;
  wire[8:0] nl_alu_loop_op_14_FpAdd_8U_23U_if_3_if_acc_2_nl;
  wire[7:0] alu_loop_op_15_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[8:0] nl_alu_loop_op_15_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[7:0] alu_loop_op_16_FpAdd_8U_23U_if_3_if_acc_2_nl;
  wire[8:0] nl_alu_loop_op_16_FpAdd_8U_23U_if_3_if_acc_2_nl;
  wire[0:0] and_876_nl;
  wire[0:0] and_878_nl;
  wire[0:0] and_891_nl;
  wire[0:0] and_893_nl;
  wire[0:0] and_906_nl;
  wire[0:0] and_908_nl;
  wire[0:0] and_921_nl;
  wire[0:0] and_923_nl;
  wire[0:0] and_925_nl;
  wire[0:0] and_927_nl;
  wire[0:0] and_929_nl;
  wire[0:0] and_931_nl;
  wire[0:0] and_933_nl;
  wire[0:0] and_935_nl;
  wire[0:0] and_948_nl;
  wire[0:0] and_950_nl;
  wire[0:0] and_952_nl;
  wire[0:0] and_954_nl;
  wire[0:0] and_956_nl;
  wire[0:0] and_958_nl;
  wire[0:0] and_960_nl;
  wire[0:0] and_962_nl;
  wire[0:0] and_964_nl;
  wire[0:0] and_966_nl;
  wire[0:0] and_979_nl;
  wire[0:0] and_981_nl;
  wire[0:0] and_994_nl;
  wire[0:0] and_996_nl;
  wire[0:0] and_1009_nl;
  wire[0:0] and_1011_nl;
  wire[0:0] and_1024_nl;
  wire[0:0] and_1026_nl;
  wire[0:0] FpAlu_8U_23U_FpAlu_8U_23U_mux_15_nl;
  wire[0:0] FpAlu_8U_23U_or_800_nl;
  wire[0:0] FpAlu_8U_23U_FpAlu_8U_23U_mux_14_nl;
  wire[0:0] FpAlu_8U_23U_or_802_nl;
  wire[0:0] FpAlu_8U_23U_FpAlu_8U_23U_mux_13_nl;
  wire[0:0] FpAlu_8U_23U_or_804_nl;
  wire[0:0] FpAlu_8U_23U_FpAlu_8U_23U_mux_12_nl;
  wire[0:0] FpAlu_8U_23U_or_806_nl;
  wire[0:0] FpAlu_8U_23U_FpAlu_8U_23U_mux_11_nl;
  wire[0:0] FpAlu_8U_23U_or_808_nl;
  wire[0:0] FpAlu_8U_23U_FpAlu_8U_23U_mux_10_nl;
  wire[0:0] FpAlu_8U_23U_or_810_nl;
  wire[0:0] FpAlu_8U_23U_FpAlu_8U_23U_mux_9_nl;
  wire[0:0] FpAlu_8U_23U_or_812_nl;
  wire[0:0] FpAlu_8U_23U_FpAlu_8U_23U_mux_8_nl;
  wire[0:0] FpAlu_8U_23U_or_814_nl;
  wire[0:0] FpAlu_8U_23U_FpAlu_8U_23U_mux_7_nl;
  wire[0:0] FpAlu_8U_23U_or_816_nl;
  wire[0:0] FpAlu_8U_23U_FpAlu_8U_23U_mux_6_nl;
  wire[0:0] FpAlu_8U_23U_or_818_nl;
  wire[0:0] FpAlu_8U_23U_FpAlu_8U_23U_mux_5_nl;
  wire[0:0] FpAlu_8U_23U_or_820_nl;
  wire[0:0] FpAlu_8U_23U_FpAlu_8U_23U_mux_4_nl;
  wire[0:0] FpAlu_8U_23U_or_822_nl;
  wire[0:0] FpAlu_8U_23U_FpAlu_8U_23U_mux_3_nl;
  wire[0:0] FpAlu_8U_23U_or_824_nl;
  wire[0:0] FpAlu_8U_23U_FpAlu_8U_23U_mux_2_nl;
  wire[0:0] FpAlu_8U_23U_or_826_nl;
  wire[0:0] FpAlu_8U_23U_FpAlu_8U_23U_mux_1_nl;
  wire[0:0] FpAlu_8U_23U_or_828_nl;
  wire[0:0] FpAlu_8U_23U_FpAlu_8U_23U_mux_nl;
  wire[0:0] FpAlu_8U_23U_or_830_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_177_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_179_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_181_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_1_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_65_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_1_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_145_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_184_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_66_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_2_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_147_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_187_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_3_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_67_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_3_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_149_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_190_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_68_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_4_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_151_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_193_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_5_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_69_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_5_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_153_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_196_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_70_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_6_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_155_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_199_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_7_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_71_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_7_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_157_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_202_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_72_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_8_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_159_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_205_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_9_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_73_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_9_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_161_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_208_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_74_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_10_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_163_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_211_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_11_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_75_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_11_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_165_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_214_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_76_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_12_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_167_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_217_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_13_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_77_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_13_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_169_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_220_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_78_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_14_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_171_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_223_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_15_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_79_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_15_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_173_nl;
  wire[29:0] alu_loop_op_1_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl;
  wire[29:0] alu_loop_op_2_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl;
  wire[29:0] alu_loop_op_3_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl;
  wire[29:0] alu_loop_op_4_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl;
  wire[29:0] alu_loop_op_5_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl;
  wire[29:0] alu_loop_op_6_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl;
  wire[29:0] alu_loop_op_7_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl;
  wire[29:0] alu_loop_op_8_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl;
  wire[29:0] alu_loop_op_9_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl;
  wire[29:0] alu_loop_op_10_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl;
  wire[29:0] alu_loop_op_11_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl;
  wire[29:0] alu_loop_op_12_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl;
  wire[29:0] alu_loop_op_13_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl;
  wire[29:0] alu_loop_op_14_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl;
  wire[29:0] alu_loop_op_15_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl;
  wire[29:0] alu_loop_op_16_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_5_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_5_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_7_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_7_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_9_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_9_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_11_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_11_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_12_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_12_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_13_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_13_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_14_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_14_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_15_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_15_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_16_nl;
  wire[22:0] alu_loop_op_1_FpMantRNE_49U_24U_else_acc_nl;
  wire[23:0] nl_alu_loop_op_1_FpMantRNE_49U_24U_else_acc_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_17_nl;
  wire[22:0] alu_loop_op_2_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[23:0] nl_alu_loop_op_2_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_18_nl;
  wire[22:0] alu_loop_op_3_FpMantRNE_49U_24U_else_acc_nl;
  wire[23:0] nl_alu_loop_op_3_FpMantRNE_49U_24U_else_acc_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_19_nl;
  wire[22:0] alu_loop_op_4_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[23:0] nl_alu_loop_op_4_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_20_nl;
  wire[22:0] alu_loop_op_5_FpMantRNE_49U_24U_else_acc_nl;
  wire[23:0] nl_alu_loop_op_5_FpMantRNE_49U_24U_else_acc_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_21_nl;
  wire[22:0] alu_loop_op_6_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[23:0] nl_alu_loop_op_6_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_22_nl;
  wire[22:0] alu_loop_op_7_FpMantRNE_49U_24U_else_acc_nl;
  wire[23:0] nl_alu_loop_op_7_FpMantRNE_49U_24U_else_acc_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_23_nl;
  wire[22:0] alu_loop_op_8_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[23:0] nl_alu_loop_op_8_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_24_nl;
  wire[22:0] alu_loop_op_9_FpMantRNE_49U_24U_else_acc_nl;
  wire[23:0] nl_alu_loop_op_9_FpMantRNE_49U_24U_else_acc_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_25_nl;
  wire[22:0] alu_loop_op_10_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[23:0] nl_alu_loop_op_10_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_26_nl;
  wire[22:0] alu_loop_op_11_FpMantRNE_49U_24U_else_acc_nl;
  wire[23:0] nl_alu_loop_op_11_FpMantRNE_49U_24U_else_acc_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_27_nl;
  wire[22:0] alu_loop_op_12_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[23:0] nl_alu_loop_op_12_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_28_nl;
  wire[22:0] alu_loop_op_13_FpMantRNE_49U_24U_else_acc_nl;
  wire[23:0] nl_alu_loop_op_13_FpMantRNE_49U_24U_else_acc_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_29_nl;
  wire[22:0] alu_loop_op_14_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[23:0] nl_alu_loop_op_14_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_30_nl;
  wire[22:0] alu_loop_op_15_FpMantRNE_49U_24U_else_acc_nl;
  wire[23:0] nl_alu_loop_op_15_FpMantRNE_49U_24U_else_acc_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_31_nl;
  wire[22:0] alu_loop_op_16_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[23:0] nl_alu_loop_op_16_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_1_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_nl;
  wire[7:0] alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[8:0] nl_alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_3_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_1_nl;
  wire[7:0] alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_2_nl;
  wire[8:0] nl_alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_2_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_5_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_2_nl;
  wire[7:0] alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[8:0] nl_alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_7_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_3_nl;
  wire[7:0] alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_2_nl;
  wire[8:0] nl_alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_2_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_9_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_4_nl;
  wire[7:0] alu_loop_op_5_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[8:0] nl_alu_loop_op_5_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_11_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_5_nl;
  wire[7:0] alu_loop_op_6_FpAdd_8U_23U_if_4_if_acc_2_nl;
  wire[8:0] nl_alu_loop_op_6_FpAdd_8U_23U_if_4_if_acc_2_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_13_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_6_nl;
  wire[7:0] alu_loop_op_7_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[8:0] nl_alu_loop_op_7_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_15_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_7_nl;
  wire[7:0] alu_loop_op_8_FpAdd_8U_23U_if_4_if_acc_2_nl;
  wire[8:0] nl_alu_loop_op_8_FpAdd_8U_23U_if_4_if_acc_2_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_17_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_8_nl;
  wire[7:0] alu_loop_op_9_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[8:0] nl_alu_loop_op_9_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_19_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_9_nl;
  wire[7:0] alu_loop_op_10_FpAdd_8U_23U_if_4_if_acc_2_nl;
  wire[8:0] nl_alu_loop_op_10_FpAdd_8U_23U_if_4_if_acc_2_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_21_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_10_nl;
  wire[7:0] alu_loop_op_11_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[8:0] nl_alu_loop_op_11_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_23_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_11_nl;
  wire[7:0] alu_loop_op_12_FpAdd_8U_23U_if_4_if_acc_2_nl;
  wire[8:0] nl_alu_loop_op_12_FpAdd_8U_23U_if_4_if_acc_2_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_25_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_12_nl;
  wire[7:0] alu_loop_op_13_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[8:0] nl_alu_loop_op_13_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_27_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_13_nl;
  wire[7:0] alu_loop_op_14_FpAdd_8U_23U_if_4_if_acc_2_nl;
  wire[8:0] nl_alu_loop_op_14_FpAdd_8U_23U_if_4_if_acc_2_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_29_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_14_nl;
  wire[7:0] alu_loop_op_15_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[8:0] nl_alu_loop_op_15_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_31_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_15_nl;
  wire[7:0] alu_loop_op_16_FpAdd_8U_23U_if_4_if_acc_2_nl;
  wire[8:0] nl_alu_loop_op_16_FpAdd_8U_23U_if_4_if_acc_2_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_111_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_95_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_110_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_94_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_109_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_93_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_108_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_92_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_107_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_91_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_106_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_90_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_105_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_89_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_104_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_88_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_103_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_87_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_102_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_86_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_101_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_85_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_100_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_84_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_99_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_83_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_98_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_82_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_97_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_81_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_96_nl;
  wire[0:0] alu_nan_to_zero_aelse_not_80_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_47_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_46_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_45_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_44_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_43_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_42_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_41_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_40_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_39_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_38_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_37_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_36_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_35_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_34_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_33_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_32_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_158_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_159_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_160_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_161_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_162_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_163_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_164_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_165_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_166_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_167_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_168_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_169_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_170_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_171_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_172_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_173_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_1_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_3_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_5_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_7_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_9_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_11_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_13_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_15_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_17_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_19_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_21_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_23_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_25_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_27_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_29_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_31_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_33_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_35_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_37_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_39_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_41_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_43_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_45_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_47_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_49_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_51_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_53_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_55_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_57_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_59_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_61_nl;
  wire[0:0] FpCmp_8U_23U_true_else_if_mux_63_nl;
  wire[23:0] FpCmp_8U_23U_false_else_else_if_acc_16_nl;
  wire[25:0] nl_FpCmp_8U_23U_false_else_else_if_acc_16_nl;
  wire[8:0] FpCmp_8U_23U_false_else_if_acc_16_nl;
  wire[10:0] nl_FpCmp_8U_23U_false_else_if_acc_16_nl;
  wire[23:0] FpCmp_8U_23U_false_else_else_if_acc_18_nl;
  wire[25:0] nl_FpCmp_8U_23U_false_else_else_if_acc_18_nl;
  wire[8:0] FpCmp_8U_23U_false_else_if_acc_18_nl;
  wire[10:0] nl_FpCmp_8U_23U_false_else_if_acc_18_nl;
  wire[23:0] FpCmp_8U_23U_false_else_else_if_acc_20_nl;
  wire[25:0] nl_FpCmp_8U_23U_false_else_else_if_acc_20_nl;
  wire[8:0] FpCmp_8U_23U_false_else_if_acc_20_nl;
  wire[10:0] nl_FpCmp_8U_23U_false_else_if_acc_20_nl;
  wire[23:0] FpCmp_8U_23U_false_else_else_if_acc_22_nl;
  wire[25:0] nl_FpCmp_8U_23U_false_else_else_if_acc_22_nl;
  wire[8:0] FpCmp_8U_23U_false_else_if_acc_22_nl;
  wire[10:0] nl_FpCmp_8U_23U_false_else_if_acc_22_nl;
  wire[23:0] FpCmp_8U_23U_false_else_else_if_acc_24_nl;
  wire[25:0] nl_FpCmp_8U_23U_false_else_else_if_acc_24_nl;
  wire[8:0] FpCmp_8U_23U_false_else_if_acc_24_nl;
  wire[10:0] nl_FpCmp_8U_23U_false_else_if_acc_24_nl;
  wire[23:0] FpCmp_8U_23U_false_else_else_if_acc_26_nl;
  wire[25:0] nl_FpCmp_8U_23U_false_else_else_if_acc_26_nl;
  wire[8:0] FpCmp_8U_23U_false_else_if_acc_26_nl;
  wire[10:0] nl_FpCmp_8U_23U_false_else_if_acc_26_nl;
  wire[23:0] FpCmp_8U_23U_false_else_else_if_acc_28_nl;
  wire[25:0] nl_FpCmp_8U_23U_false_else_else_if_acc_28_nl;
  wire[8:0] FpCmp_8U_23U_false_else_if_acc_28_nl;
  wire[10:0] nl_FpCmp_8U_23U_false_else_if_acc_28_nl;
  wire[23:0] FpCmp_8U_23U_false_else_else_if_acc_30_nl;
  wire[25:0] nl_FpCmp_8U_23U_false_else_else_if_acc_30_nl;
  wire[8:0] FpCmp_8U_23U_false_else_if_acc_30_nl;
  wire[10:0] nl_FpCmp_8U_23U_false_else_if_acc_30_nl;
  wire[23:0] FpCmp_8U_23U_false_else_else_if_acc_32_nl;
  wire[25:0] nl_FpCmp_8U_23U_false_else_else_if_acc_32_nl;
  wire[8:0] FpCmp_8U_23U_false_else_if_acc_32_nl;
  wire[10:0] nl_FpCmp_8U_23U_false_else_if_acc_32_nl;
  wire[23:0] FpCmp_8U_23U_false_else_else_if_acc_34_nl;
  wire[25:0] nl_FpCmp_8U_23U_false_else_else_if_acc_34_nl;
  wire[8:0] FpCmp_8U_23U_false_else_if_acc_34_nl;
  wire[10:0] nl_FpCmp_8U_23U_false_else_if_acc_34_nl;
  wire[23:0] FpCmp_8U_23U_false_else_else_if_acc_36_nl;
  wire[25:0] nl_FpCmp_8U_23U_false_else_else_if_acc_36_nl;
  wire[8:0] FpCmp_8U_23U_false_else_if_acc_36_nl;
  wire[10:0] nl_FpCmp_8U_23U_false_else_if_acc_36_nl;
  wire[23:0] FpCmp_8U_23U_false_else_else_if_acc_38_nl;
  wire[25:0] nl_FpCmp_8U_23U_false_else_else_if_acc_38_nl;
  wire[8:0] FpCmp_8U_23U_false_else_if_acc_38_nl;
  wire[10:0] nl_FpCmp_8U_23U_false_else_if_acc_38_nl;
  wire[23:0] FpCmp_8U_23U_false_else_else_if_acc_40_nl;
  wire[25:0] nl_FpCmp_8U_23U_false_else_else_if_acc_40_nl;
  wire[8:0] FpCmp_8U_23U_false_else_if_acc_40_nl;
  wire[10:0] nl_FpCmp_8U_23U_false_else_if_acc_40_nl;
  wire[23:0] FpCmp_8U_23U_false_else_else_if_acc_42_nl;
  wire[25:0] nl_FpCmp_8U_23U_false_else_else_if_acc_42_nl;
  wire[8:0] FpCmp_8U_23U_false_else_if_acc_42_nl;
  wire[10:0] nl_FpCmp_8U_23U_false_else_if_acc_42_nl;
  wire[23:0] FpCmp_8U_23U_false_else_else_if_acc_44_nl;
  wire[25:0] nl_FpCmp_8U_23U_false_else_else_if_acc_44_nl;
  wire[8:0] FpCmp_8U_23U_false_else_if_acc_44_nl;
  wire[10:0] nl_FpCmp_8U_23U_false_else_if_acc_44_nl;
  wire[23:0] FpCmp_8U_23U_false_else_else_if_acc_46_nl;
  wire[25:0] nl_FpCmp_8U_23U_false_else_else_if_acc_46_nl;
  wire[8:0] FpCmp_8U_23U_false_else_if_acc_46_nl;
  wire[10:0] nl_FpCmp_8U_23U_false_else_if_acc_46_nl;
  wire[8:0] FpCmp_8U_23U_true_if_acc_16_nl;
  wire[10:0] nl_FpCmp_8U_23U_true_if_acc_16_nl;
  wire[8:0] FpCmp_8U_23U_true_if_acc_18_nl;
  wire[10:0] nl_FpCmp_8U_23U_true_if_acc_18_nl;
  wire[8:0] FpCmp_8U_23U_true_if_acc_20_nl;
  wire[10:0] nl_FpCmp_8U_23U_true_if_acc_20_nl;
  wire[8:0] FpCmp_8U_23U_true_if_acc_22_nl;
  wire[10:0] nl_FpCmp_8U_23U_true_if_acc_22_nl;
  wire[8:0] FpCmp_8U_23U_true_if_acc_24_nl;
  wire[10:0] nl_FpCmp_8U_23U_true_if_acc_24_nl;
  wire[8:0] FpCmp_8U_23U_true_if_acc_26_nl;
  wire[10:0] nl_FpCmp_8U_23U_true_if_acc_26_nl;
  wire[8:0] FpCmp_8U_23U_true_if_acc_28_nl;
  wire[10:0] nl_FpCmp_8U_23U_true_if_acc_28_nl;
  wire[8:0] FpCmp_8U_23U_true_if_acc_30_nl;
  wire[10:0] nl_FpCmp_8U_23U_true_if_acc_30_nl;
  wire[8:0] FpCmp_8U_23U_true_if_acc_32_nl;
  wire[10:0] nl_FpCmp_8U_23U_true_if_acc_32_nl;
  wire[8:0] FpCmp_8U_23U_true_if_acc_34_nl;
  wire[10:0] nl_FpCmp_8U_23U_true_if_acc_34_nl;
  wire[8:0] FpCmp_8U_23U_true_if_acc_36_nl;
  wire[10:0] nl_FpCmp_8U_23U_true_if_acc_36_nl;
  wire[8:0] FpCmp_8U_23U_true_if_acc_38_nl;
  wire[10:0] nl_FpCmp_8U_23U_true_if_acc_38_nl;
  wire[8:0] FpCmp_8U_23U_true_if_acc_40_nl;
  wire[10:0] nl_FpCmp_8U_23U_true_if_acc_40_nl;
  wire[8:0] FpCmp_8U_23U_true_if_acc_42_nl;
  wire[10:0] nl_FpCmp_8U_23U_true_if_acc_42_nl;
  wire[8:0] FpCmp_8U_23U_true_if_acc_44_nl;
  wire[10:0] nl_FpCmp_8U_23U_true_if_acc_44_nl;
  wire[8:0] FpCmp_8U_23U_true_if_acc_46_nl;
  wire[10:0] nl_FpCmp_8U_23U_true_if_acc_46_nl;
  wire[8:0] alu_loop_op_1_FpNormalize_8U_49U_acc_nl;
  wire[10:0] nl_alu_loop_op_1_FpNormalize_8U_49U_acc_nl;
  wire[8:0] alu_loop_op_2_FpNormalize_8U_49U_acc_1_nl;
  wire[10:0] nl_alu_loop_op_2_FpNormalize_8U_49U_acc_1_nl;
  wire[8:0] alu_loop_op_3_FpNormalize_8U_49U_acc_nl;
  wire[10:0] nl_alu_loop_op_3_FpNormalize_8U_49U_acc_nl;
  wire[8:0] alu_loop_op_4_FpNormalize_8U_49U_acc_1_nl;
  wire[10:0] nl_alu_loop_op_4_FpNormalize_8U_49U_acc_1_nl;
  wire[8:0] alu_loop_op_5_FpNormalize_8U_49U_acc_nl;
  wire[10:0] nl_alu_loop_op_5_FpNormalize_8U_49U_acc_nl;
  wire[8:0] alu_loop_op_6_FpNormalize_8U_49U_acc_1_nl;
  wire[10:0] nl_alu_loop_op_6_FpNormalize_8U_49U_acc_1_nl;
  wire[8:0] alu_loop_op_7_FpNormalize_8U_49U_acc_nl;
  wire[10:0] nl_alu_loop_op_7_FpNormalize_8U_49U_acc_nl;
  wire[8:0] alu_loop_op_8_FpNormalize_8U_49U_acc_1_nl;
  wire[10:0] nl_alu_loop_op_8_FpNormalize_8U_49U_acc_1_nl;
  wire[8:0] alu_loop_op_9_FpNormalize_8U_49U_acc_nl;
  wire[10:0] nl_alu_loop_op_9_FpNormalize_8U_49U_acc_nl;
  wire[8:0] alu_loop_op_10_FpNormalize_8U_49U_acc_1_nl;
  wire[10:0] nl_alu_loop_op_10_FpNormalize_8U_49U_acc_1_nl;
  wire[8:0] alu_loop_op_11_FpNormalize_8U_49U_acc_nl;
  wire[10:0] nl_alu_loop_op_11_FpNormalize_8U_49U_acc_nl;
  wire[8:0] alu_loop_op_12_FpNormalize_8U_49U_acc_1_nl;
  wire[10:0] nl_alu_loop_op_12_FpNormalize_8U_49U_acc_1_nl;
  wire[8:0] alu_loop_op_13_FpNormalize_8U_49U_acc_nl;
  wire[10:0] nl_alu_loop_op_13_FpNormalize_8U_49U_acc_nl;
  wire[8:0] alu_loop_op_14_FpNormalize_8U_49U_acc_1_nl;
  wire[10:0] nl_alu_loop_op_14_FpNormalize_8U_49U_acc_1_nl;
  wire[8:0] alu_loop_op_15_FpNormalize_8U_49U_acc_nl;
  wire[10:0] nl_alu_loop_op_15_FpNormalize_8U_49U_acc_nl;
  wire[8:0] alu_loop_op_16_FpNormalize_8U_49U_acc_1_nl;
  wire[10:0] nl_alu_loop_op_16_FpNormalize_8U_49U_acc_1_nl;
  wire[32:0] alu_loop_op_16_else_if_acc_1_nl;
  wire[33:0] nl_alu_loop_op_16_else_if_acc_1_nl;
  wire[32:0] alu_loop_op_16_else_else_if_acc_1_nl;
  wire[34:0] nl_alu_loop_op_16_else_else_if_acc_1_nl;
  wire[32:0] alu_loop_op_15_else_if_acc_nl;
  wire[33:0] nl_alu_loop_op_15_else_if_acc_nl;
  wire[32:0] alu_loop_op_15_else_else_if_acc_nl;
  wire[34:0] nl_alu_loop_op_15_else_else_if_acc_nl;
  wire[32:0] alu_loop_op_14_else_if_acc_1_nl;
  wire[33:0] nl_alu_loop_op_14_else_if_acc_1_nl;
  wire[32:0] alu_loop_op_14_else_else_if_acc_1_nl;
  wire[34:0] nl_alu_loop_op_14_else_else_if_acc_1_nl;
  wire[32:0] alu_loop_op_13_else_if_acc_nl;
  wire[33:0] nl_alu_loop_op_13_else_if_acc_nl;
  wire[32:0] alu_loop_op_13_else_else_if_acc_nl;
  wire[34:0] nl_alu_loop_op_13_else_else_if_acc_nl;
  wire[32:0] alu_loop_op_12_else_if_acc_1_nl;
  wire[33:0] nl_alu_loop_op_12_else_if_acc_1_nl;
  wire[32:0] alu_loop_op_12_else_else_if_acc_1_nl;
  wire[34:0] nl_alu_loop_op_12_else_else_if_acc_1_nl;
  wire[32:0] alu_loop_op_11_else_if_acc_nl;
  wire[33:0] nl_alu_loop_op_11_else_if_acc_nl;
  wire[32:0] alu_loop_op_11_else_else_if_acc_nl;
  wire[34:0] nl_alu_loop_op_11_else_else_if_acc_nl;
  wire[32:0] alu_loop_op_10_else_if_acc_1_nl;
  wire[33:0] nl_alu_loop_op_10_else_if_acc_1_nl;
  wire[32:0] alu_loop_op_10_else_else_if_acc_1_nl;
  wire[34:0] nl_alu_loop_op_10_else_else_if_acc_1_nl;
  wire[32:0] alu_loop_op_9_else_if_acc_nl;
  wire[33:0] nl_alu_loop_op_9_else_if_acc_nl;
  wire[32:0] alu_loop_op_9_else_else_if_acc_nl;
  wire[34:0] nl_alu_loop_op_9_else_else_if_acc_nl;
  wire[32:0] alu_loop_op_8_else_if_acc_1_nl;
  wire[33:0] nl_alu_loop_op_8_else_if_acc_1_nl;
  wire[32:0] alu_loop_op_8_else_else_if_acc_1_nl;
  wire[34:0] nl_alu_loop_op_8_else_else_if_acc_1_nl;
  wire[32:0] alu_loop_op_7_else_if_acc_nl;
  wire[33:0] nl_alu_loop_op_7_else_if_acc_nl;
  wire[32:0] alu_loop_op_7_else_else_if_acc_nl;
  wire[34:0] nl_alu_loop_op_7_else_else_if_acc_nl;
  wire[32:0] alu_loop_op_6_else_if_acc_1_nl;
  wire[33:0] nl_alu_loop_op_6_else_if_acc_1_nl;
  wire[32:0] alu_loop_op_6_else_else_if_acc_1_nl;
  wire[34:0] nl_alu_loop_op_6_else_else_if_acc_1_nl;
  wire[32:0] alu_loop_op_5_else_if_acc_nl;
  wire[33:0] nl_alu_loop_op_5_else_if_acc_nl;
  wire[32:0] alu_loop_op_5_else_else_if_acc_nl;
  wire[34:0] nl_alu_loop_op_5_else_else_if_acc_nl;
  wire[32:0] alu_loop_op_4_else_if_acc_1_nl;
  wire[33:0] nl_alu_loop_op_4_else_if_acc_1_nl;
  wire[32:0] alu_loop_op_4_else_else_if_acc_1_nl;
  wire[34:0] nl_alu_loop_op_4_else_else_if_acc_1_nl;
  wire[32:0] alu_loop_op_3_else_if_acc_nl;
  wire[33:0] nl_alu_loop_op_3_else_if_acc_nl;
  wire[32:0] alu_loop_op_3_else_else_if_acc_nl;
  wire[34:0] nl_alu_loop_op_3_else_else_if_acc_nl;
  wire[32:0] alu_loop_op_2_else_if_acc_1_nl;
  wire[33:0] nl_alu_loop_op_2_else_if_acc_1_nl;
  wire[32:0] alu_loop_op_2_else_else_if_acc_1_nl;
  wire[34:0] nl_alu_loop_op_2_else_else_if_acc_1_nl;
  wire[32:0] alu_loop_op_1_else_if_acc_nl;
  wire[33:0] nl_alu_loop_op_1_else_if_acc_nl;
  wire[32:0] alu_loop_op_1_else_else_if_acc_nl;
  wire[34:0] nl_alu_loop_op_1_else_else_if_acc_nl;
  wire[0:0] nor_2056_nl;
  wire[0:0] nor_2057_nl;
  wire[0:0] or_32_nl;
  wire[0:0] or_341_nl;
  wire[0:0] nor_1962_nl;
  wire[0:0] mux_392_nl;
  wire[0:0] or_902_nl;
  wire[0:0] or_904_nl;
  wire[0:0] and_224_nl;
  wire[0:0] and_225_nl;
  wire[0:0] mux_414_nl;
  wire[0:0] mux_784_nl;
  wire[0:0] or_1868_nl;
  wire[0:0] nor_1329_nl;
  wire[0:0] or_1872_nl;
  wire[0:0] nor_1327_nl;
  wire[0:0] mux_787_nl;
  wire[0:0] or_1876_nl;
  wire[0:0] and_284_nl;
  wire[0:0] or_1879_nl;
  wire[0:0] and_285_nl;
  wire[0:0] or_1882_nl;
  wire[0:0] and_286_nl;
  wire[0:0] mux_791_nl;
  wire[0:0] or_1884_nl;
  wire[0:0] and_3691_nl;
  wire[0:0] or_1886_nl;
  wire[0:0] nor_1326_nl;
  wire[0:0] or_1890_nl;
  wire[0:0] nor_1325_nl;
  wire[0:0] or_1894_nl;
  wire[0:0] nor_1324_nl;
  wire[0:0] or_1899_nl;
  wire[0:0] and_287_nl;
  wire[0:0] or_1901_nl;
  wire[0:0] nor_1323_nl;
  wire[0:0] or_1905_nl;
  wire[0:0] nor_1322_nl;
  wire[0:0] or_1909_nl;
  wire[0:0] nor_1321_nl;
  wire[0:0] or_1913_nl;
  wire[0:0] nor_1320_nl;
  wire[0:0] mux_801_nl;
  wire[0:0] or_1915_nl;
  wire[0:0] and_3690_nl;
  wire[0:0] or_1917_nl;
  wire[0:0] nor_1319_nl;
  wire[0:0] mux_829_nl;
  wire[0:0] or_2494_nl;
  wire[0:0] and_3623_nl;
  wire[0:0] mux_1424_nl;
  wire[0:0] or_2855_nl;
  wire[0:0] and_3551_nl;
  wire[0:0] mux_1522_nl;
  wire[0:0] nor_913_nl;
  wire[0:0] and_3550_nl;
  wire[0:0] mux_1523_nl;
  wire[0:0] nor_911_nl;
  wire[0:0] nor_912_nl;
  wire[0:0] mux_1524_nl;
  wire[0:0] nor_910_nl;
  wire[0:0] and_3549_nl;
  wire[0:0] mux_1525_nl;
  wire[0:0] nor_908_nl;
  wire[0:0] nor_909_nl;
  wire[0:0] mux_1526_nl;
  wire[0:0] nor_907_nl;
  wire[0:0] and_3548_nl;
  wire[0:0] mux_1527_nl;
  wire[0:0] nor_905_nl;
  wire[0:0] nor_906_nl;
  wire[0:0] mux_1528_nl;
  wire[0:0] nor_904_nl;
  wire[0:0] and_3547_nl;
  wire[0:0] mux_1529_nl;
  wire[0:0] nor_902_nl;
  wire[0:0] nor_903_nl;
  wire[0:0] mux_1530_nl;
  wire[0:0] nor_901_nl;
  wire[0:0] and_3546_nl;
  wire[0:0] mux_1531_nl;
  wire[0:0] nor_899_nl;
  wire[0:0] nor_900_nl;
  wire[0:0] mux_1532_nl;
  wire[0:0] nor_898_nl;
  wire[0:0] and_3545_nl;
  wire[0:0] mux_1533_nl;
  wire[0:0] nor_896_nl;
  wire[0:0] nor_897_nl;
  wire[0:0] mux_1534_nl;
  wire[0:0] nor_895_nl;
  wire[0:0] and_3544_nl;
  wire[0:0] mux_1535_nl;
  wire[0:0] nor_893_nl;
  wire[0:0] nor_894_nl;
  wire[0:0] mux_1536_nl;
  wire[0:0] nor_892_nl;
  wire[0:0] and_3543_nl;
  wire[0:0] mux_1537_nl;
  wire[0:0] nor_890_nl;
  wire[0:0] nor_891_nl;
  wire[0:0] mux_1538_nl;
  wire[0:0] nor_889_nl;
  wire[0:0] and_3542_nl;
  wire[0:0] mux_1539_nl;
  wire[0:0] nor_887_nl;
  wire[0:0] nor_888_nl;
  wire[0:0] mux_1540_nl;
  wire[0:0] nor_886_nl;
  wire[0:0] and_3541_nl;
  wire[0:0] mux_1541_nl;
  wire[0:0] nor_884_nl;
  wire[0:0] nor_885_nl;
  wire[0:0] mux_1542_nl;
  wire[0:0] nor_883_nl;
  wire[0:0] and_3540_nl;
  wire[0:0] mux_1543_nl;
  wire[0:0] nor_881_nl;
  wire[0:0] nor_882_nl;
  wire[0:0] mux_1544_nl;
  wire[0:0] nor_880_nl;
  wire[0:0] and_3539_nl;
  wire[0:0] mux_1545_nl;
  wire[0:0] nor_878_nl;
  wire[0:0] nor_879_nl;
  wire[0:0] mux_1546_nl;
  wire[0:0] nor_877_nl;
  wire[0:0] mux_1547_nl;
  wire[0:0] nor_875_nl;
  wire[0:0] nor_876_nl;
  wire[8:0] acc_nl;
  wire[9:0] nl_acc_nl;
  wire[0:0] FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_16_nl;
  wire[5:0] FpAdd_8U_23U_if_3_if_mux_64_nl;
  wire[8:0] acc_1_nl;
  wire[9:0] nl_acc_1_nl;
  wire[0:0] FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_17_nl;
  wire[5:0] FpAdd_8U_23U_if_3_if_mux_65_nl;
  wire[8:0] acc_2_nl;
  wire[9:0] nl_acc_2_nl;
  wire[0:0] FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_18_nl;
  wire[5:0] FpAdd_8U_23U_if_3_if_mux_66_nl;
  wire[8:0] acc_3_nl;
  wire[9:0] nl_acc_3_nl;
  wire[0:0] FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_19_nl;
  wire[5:0] FpAdd_8U_23U_if_3_if_mux_67_nl;
  wire[8:0] acc_4_nl;
  wire[9:0] nl_acc_4_nl;
  wire[0:0] FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_20_nl;
  wire[5:0] FpAdd_8U_23U_if_3_if_mux_68_nl;
  wire[8:0] acc_5_nl;
  wire[9:0] nl_acc_5_nl;
  wire[0:0] FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_21_nl;
  wire[5:0] FpAdd_8U_23U_if_3_if_mux_69_nl;
  wire[8:0] acc_6_nl;
  wire[9:0] nl_acc_6_nl;
  wire[0:0] FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_22_nl;
  wire[5:0] FpAdd_8U_23U_if_3_if_mux_70_nl;
  wire[8:0] acc_7_nl;
  wire[9:0] nl_acc_7_nl;
  wire[0:0] FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_23_nl;
  wire[5:0] FpAdd_8U_23U_if_3_if_mux_71_nl;
  wire[8:0] acc_8_nl;
  wire[9:0] nl_acc_8_nl;
  wire[0:0] FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_24_nl;
  wire[5:0] FpAdd_8U_23U_if_3_if_mux_72_nl;
  wire[8:0] acc_9_nl;
  wire[9:0] nl_acc_9_nl;
  wire[0:0] FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_25_nl;
  wire[5:0] FpAdd_8U_23U_if_3_if_mux_73_nl;
  wire[8:0] acc_10_nl;
  wire[9:0] nl_acc_10_nl;
  wire[0:0] FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_26_nl;
  wire[5:0] FpAdd_8U_23U_if_3_if_mux_74_nl;
  wire[8:0] acc_11_nl;
  wire[9:0] nl_acc_11_nl;
  wire[0:0] FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_27_nl;
  wire[5:0] FpAdd_8U_23U_if_3_if_mux_75_nl;
  wire[8:0] acc_12_nl;
  wire[9:0] nl_acc_12_nl;
  wire[0:0] FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_28_nl;
  wire[5:0] FpAdd_8U_23U_if_3_if_mux_76_nl;
  wire[8:0] acc_13_nl;
  wire[9:0] nl_acc_13_nl;
  wire[0:0] FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_29_nl;
  wire[5:0] FpAdd_8U_23U_if_3_if_mux_77_nl;
  wire[8:0] acc_14_nl;
  wire[9:0] nl_acc_14_nl;
  wire[0:0] FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_30_nl;
  wire[5:0] FpAdd_8U_23U_if_3_if_mux_78_nl;
  wire[8:0] acc_15_nl;
  wire[9:0] nl_acc_15_nl;
  wire[0:0] FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_31_nl;
  wire[5:0] FpAdd_8U_23U_if_3_if_mux_79_nl;
  wire[8:0] acc_16_nl;
  wire[9:0] nl_acc_16_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_32_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_33_nl;
  wire[8:0] acc_17_nl;
  wire[9:0] nl_acc_17_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_34_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_35_nl;
  wire[8:0] acc_18_nl;
  wire[9:0] nl_acc_18_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_36_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_37_nl;
  wire[8:0] acc_19_nl;
  wire[9:0] nl_acc_19_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_38_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_39_nl;
  wire[8:0] acc_20_nl;
  wire[9:0] nl_acc_20_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_40_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_41_nl;
  wire[8:0] acc_21_nl;
  wire[9:0] nl_acc_21_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_42_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_43_nl;
  wire[8:0] acc_22_nl;
  wire[9:0] nl_acc_22_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_44_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_45_nl;
  wire[8:0] acc_23_nl;
  wire[9:0] nl_acc_23_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_46_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_47_nl;
  wire[8:0] acc_24_nl;
  wire[9:0] nl_acc_24_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_48_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_49_nl;
  wire[8:0] acc_25_nl;
  wire[9:0] nl_acc_25_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_50_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_51_nl;
  wire[8:0] acc_26_nl;
  wire[9:0] nl_acc_26_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_52_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_53_nl;
  wire[8:0] acc_27_nl;
  wire[9:0] nl_acc_27_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_54_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_55_nl;
  wire[8:0] acc_28_nl;
  wire[9:0] nl_acc_28_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_56_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_57_nl;
  wire[8:0] acc_29_nl;
  wire[9:0] nl_acc_29_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_58_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_59_nl;
  wire[8:0] acc_30_nl;
  wire[9:0] nl_acc_30_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_60_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_61_nl;
  wire[8:0] acc_31_nl;
  wire[9:0] nl_acc_31_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_62_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_63_nl;
// Interconnect Declarations for Component Instantiations
  wire [23:0] nl_alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  assign nl_alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = {alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp_2};
  wire [8:0] nl_alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  assign nl_alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = {alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_itm_2
      , (~ alu_loop_op_1_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2)};
  wire [23:0] nl_alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  assign nl_alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = {alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5
      , (AluIn_data_sva_502[22:0])};
  wire [8:0] nl_alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  assign nl_alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = {alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_itm_2
      , (~ alu_loop_op_1_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2)};
  wire [23:0] nl_alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a;
  assign nl_alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a = {IsNaN_8U_23U_3_land_2_lpi_1_dfm_7
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp_2};
  wire [8:0] nl_alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s;
  assign nl_alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s = {alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_1_itm_2
      , (~ alu_loop_op_2_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2)};
  wire [23:0] nl_alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a;
  assign nl_alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a = {alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5
      , (AluIn_data_sva_502[54:32])};
  wire [8:0] nl_alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s;
  assign nl_alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s = {alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_1_itm_2
      , (~ alu_loop_op_2_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2)};
  wire [23:0] nl_alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  assign nl_alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = {alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp_2};
  wire [8:0] nl_alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  assign nl_alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = {alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_itm_2
      , (~ alu_loop_op_3_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2)};
  wire [23:0] nl_alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  assign nl_alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = {alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5
      , (AluIn_data_sva_502[86:64])};
  wire [8:0] nl_alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  assign nl_alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = {alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_itm_2
      , (~ alu_loop_op_3_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2)};
  wire [23:0] nl_alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a;
  assign nl_alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a = {IsNaN_8U_23U_3_land_4_lpi_1_dfm_7
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp_2};
  wire [8:0] nl_alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s;
  assign nl_alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s = {alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_1_itm_2
      , (~ alu_loop_op_4_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2)};
  wire [23:0] nl_alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a;
  assign nl_alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a = {alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5
      , (AluIn_data_sva_502[118:96])};
  wire [8:0] nl_alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s;
  assign nl_alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s = {alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_1_itm_2
      , (~ alu_loop_op_4_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2)};
  wire [23:0] nl_alu_loop_op_5_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  assign nl_alu_loop_op_5_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = {IsNaN_8U_23U_3_land_5_lpi_1_dfm_7
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp_2};
  wire [8:0] nl_alu_loop_op_5_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  assign nl_alu_loop_op_5_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = {alu_loop_op_5_FpAdd_8U_23U_b_left_shift_acc_itm_2
      , (~ alu_loop_op_5_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2)};
  wire [23:0] nl_alu_loop_op_5_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  assign nl_alu_loop_op_5_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = {alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5
      , (AluIn_data_sva_502[150:128])};
  wire [8:0] nl_alu_loop_op_5_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  assign nl_alu_loop_op_5_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = {alu_loop_op_5_FpAdd_8U_23U_a_left_shift_acc_itm_2
      , (~ alu_loop_op_5_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2)};
  wire [23:0] nl_alu_loop_op_6_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a;
  assign nl_alu_loop_op_6_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a = {IsNaN_8U_23U_3_land_6_lpi_1_dfm_7
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp_2};
  wire [8:0] nl_alu_loop_op_6_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s;
  assign nl_alu_loop_op_6_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s = {alu_loop_op_6_FpAdd_8U_23U_b_left_shift_acc_1_itm_2
      , (~ alu_loop_op_6_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2)};
  wire [23:0] nl_alu_loop_op_6_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a;
  assign nl_alu_loop_op_6_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a = {alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5
      , (AluIn_data_sva_502[182:160])};
  wire [8:0] nl_alu_loop_op_6_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s;
  assign nl_alu_loop_op_6_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s = {alu_loop_op_6_FpAdd_8U_23U_a_left_shift_acc_1_itm_2
      , (~ alu_loop_op_6_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2)};
  wire [23:0] nl_alu_loop_op_7_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  assign nl_alu_loop_op_7_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = {alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp_2};
  wire [8:0] nl_alu_loop_op_7_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  assign nl_alu_loop_op_7_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = {alu_loop_op_7_FpAdd_8U_23U_b_left_shift_acc_itm_2
      , (~ alu_loop_op_7_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2)};
  wire [23:0] nl_alu_loop_op_7_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  assign nl_alu_loop_op_7_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = {alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5
      , (AluIn_data_sva_502[214:192])};
  wire [8:0] nl_alu_loop_op_7_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  assign nl_alu_loop_op_7_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = {alu_loop_op_7_FpAdd_8U_23U_a_left_shift_acc_itm_2
      , (~ alu_loop_op_7_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2)};
  wire [23:0] nl_alu_loop_op_8_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a;
  assign nl_alu_loop_op_8_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a = {alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp_2};
  wire [8:0] nl_alu_loop_op_8_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s;
  assign nl_alu_loop_op_8_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s = {alu_loop_op_8_FpAdd_8U_23U_b_left_shift_acc_1_itm_2
      , (~ alu_loop_op_8_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2)};
  wire [23:0] nl_alu_loop_op_8_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a;
  assign nl_alu_loop_op_8_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a = {alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5
      , (AluIn_data_sva_502[246:224])};
  wire [8:0] nl_alu_loop_op_8_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s;
  assign nl_alu_loop_op_8_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s = {alu_loop_op_8_FpAdd_8U_23U_a_left_shift_acc_1_itm_2
      , (~ alu_loop_op_8_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2)};
  wire [23:0] nl_alu_loop_op_9_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  assign nl_alu_loop_op_9_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = {IsNaN_8U_23U_3_land_9_lpi_1_dfm_7
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp_2};
  wire [8:0] nl_alu_loop_op_9_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  assign nl_alu_loop_op_9_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = {alu_loop_op_9_FpAdd_8U_23U_b_left_shift_acc_itm_2
      , (~ alu_loop_op_9_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2)};
  wire [23:0] nl_alu_loop_op_9_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  assign nl_alu_loop_op_9_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = {alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5
      , (AluIn_data_sva_502[278:256])};
  wire [8:0] nl_alu_loop_op_9_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  assign nl_alu_loop_op_9_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = {alu_loop_op_9_FpAdd_8U_23U_a_left_shift_acc_itm_2
      , (~ alu_loop_op_9_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2)};
  wire [23:0] nl_alu_loop_op_10_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a;
  assign nl_alu_loop_op_10_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a = {IsNaN_8U_23U_3_land_10_lpi_1_dfm_7
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp_2};
  wire [8:0] nl_alu_loop_op_10_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s;
  assign nl_alu_loop_op_10_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s = {alu_loop_op_10_FpAdd_8U_23U_b_left_shift_acc_1_itm_2
      , (~ alu_loop_op_10_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2)};
  wire [23:0] nl_alu_loop_op_10_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a;
  assign nl_alu_loop_op_10_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a = {alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5
      , (AluIn_data_sva_502[310:288])};
  wire [8:0] nl_alu_loop_op_10_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s;
  assign nl_alu_loop_op_10_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s = {alu_loop_op_10_FpAdd_8U_23U_a_left_shift_acc_1_itm_2
      , (~ alu_loop_op_10_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2)};
  wire [23:0] nl_alu_loop_op_11_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  assign nl_alu_loop_op_11_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = {IsNaN_8U_23U_3_land_11_lpi_1_dfm_7
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp_2};
  wire [8:0] nl_alu_loop_op_11_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  assign nl_alu_loop_op_11_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = {alu_loop_op_11_FpAdd_8U_23U_b_left_shift_acc_itm_2
      , (~ alu_loop_op_11_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2)};
  wire [23:0] nl_alu_loop_op_11_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  assign nl_alu_loop_op_11_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = {alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5
      , (AluIn_data_sva_502[342:320])};
  wire [8:0] nl_alu_loop_op_11_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  assign nl_alu_loop_op_11_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = {alu_loop_op_11_FpAdd_8U_23U_a_left_shift_acc_itm_2
      , (~ alu_loop_op_11_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2)};
  wire [23:0] nl_alu_loop_op_12_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a;
  assign nl_alu_loop_op_12_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a = {IsNaN_8U_23U_3_land_12_lpi_1_dfm_7
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp_2};
  wire [8:0] nl_alu_loop_op_12_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s;
  assign nl_alu_loop_op_12_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s = {alu_loop_op_12_FpAdd_8U_23U_b_left_shift_acc_1_itm_2
      , (~ alu_loop_op_12_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2)};
  wire [23:0] nl_alu_loop_op_12_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a;
  assign nl_alu_loop_op_12_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a = {alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5
      , (AluIn_data_sva_502[374:352])};
  wire [8:0] nl_alu_loop_op_12_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s;
  assign nl_alu_loop_op_12_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s = {alu_loop_op_12_FpAdd_8U_23U_a_left_shift_acc_1_itm_2
      , (~ alu_loop_op_12_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2)};
  wire [23:0] nl_alu_loop_op_13_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  assign nl_alu_loop_op_13_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = {IsNaN_8U_23U_3_land_13_lpi_1_dfm_7
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp_2};
  wire [8:0] nl_alu_loop_op_13_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  assign nl_alu_loop_op_13_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = {alu_loop_op_13_FpAdd_8U_23U_b_left_shift_acc_itm_2
      , (~ alu_loop_op_13_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2)};
  wire [23:0] nl_alu_loop_op_13_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  assign nl_alu_loop_op_13_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = {alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5
      , (AluIn_data_sva_502[406:384])};
  wire [8:0] nl_alu_loop_op_13_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  assign nl_alu_loop_op_13_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = {alu_loop_op_13_FpAdd_8U_23U_a_left_shift_acc_itm_2
      , (~ alu_loop_op_13_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2)};
  wire [23:0] nl_alu_loop_op_14_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a;
  assign nl_alu_loop_op_14_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a = {IsNaN_8U_23U_3_land_14_lpi_1_dfm_7
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp_2};
  wire [8:0] nl_alu_loop_op_14_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s;
  assign nl_alu_loop_op_14_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s = {alu_loop_op_14_FpAdd_8U_23U_b_left_shift_acc_1_itm_2
      , (~ alu_loop_op_14_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2)};
  wire [23:0] nl_alu_loop_op_14_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a;
  assign nl_alu_loop_op_14_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a = {alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5
      , (AluIn_data_sva_502[438:416])};
  wire [8:0] nl_alu_loop_op_14_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s;
  assign nl_alu_loop_op_14_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s = {alu_loop_op_14_FpAdd_8U_23U_a_left_shift_acc_1_itm_2
      , (~ alu_loop_op_14_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2)};
  wire [23:0] nl_alu_loop_op_15_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  assign nl_alu_loop_op_15_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = {alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp_2};
  wire [8:0] nl_alu_loop_op_15_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  assign nl_alu_loop_op_15_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = {alu_loop_op_15_FpAdd_8U_23U_b_left_shift_acc_itm_2
      , (~ alu_loop_op_15_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2)};
  wire [23:0] nl_alu_loop_op_15_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  assign nl_alu_loop_op_15_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = {alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5
      , (AluIn_data_sva_502[470:448])};
  wire [8:0] nl_alu_loop_op_15_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  assign nl_alu_loop_op_15_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = {alu_loop_op_15_FpAdd_8U_23U_a_left_shift_acc_itm_2
      , (~ alu_loop_op_15_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2)};
  wire [23:0] nl_alu_loop_op_16_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a;
  assign nl_alu_loop_op_16_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a = {alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp_2};
  wire [8:0] nl_alu_loop_op_16_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s;
  assign nl_alu_loop_op_16_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s = {alu_loop_op_16_FpAdd_8U_23U_b_left_shift_acc_1_itm_2
      , (~ alu_loop_op_16_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2)};
  wire [23:0] nl_alu_loop_op_16_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a;
  assign nl_alu_loop_op_16_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a = {alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5
      , (AluIn_data_sva_502[502:480])};
  wire [8:0] nl_alu_loop_op_16_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s;
  assign nl_alu_loop_op_16_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s = {alu_loop_op_16_FpAdd_8U_23U_a_left_shift_acc_1_itm_2
      , (~ alu_loop_op_16_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2)};
  wire [48:0] nl_alu_loop_op_1_FpNormalize_8U_49U_else_lshift_rg_a;
  assign nl_alu_loop_op_1_FpNormalize_8U_49U_else_lshift_rg_a = FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_2_FpNormalize_8U_49U_else_lshift_1_rg_a;
  assign nl_alu_loop_op_2_FpNormalize_8U_49U_else_lshift_1_rg_a = FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_3_FpNormalize_8U_49U_else_lshift_rg_a;
  assign nl_alu_loop_op_3_FpNormalize_8U_49U_else_lshift_rg_a = FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_4_FpNormalize_8U_49U_else_lshift_1_rg_a;
  assign nl_alu_loop_op_4_FpNormalize_8U_49U_else_lshift_1_rg_a = FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_5_FpNormalize_8U_49U_else_lshift_rg_a;
  assign nl_alu_loop_op_5_FpNormalize_8U_49U_else_lshift_rg_a = FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_6_FpNormalize_8U_49U_else_lshift_1_rg_a;
  assign nl_alu_loop_op_6_FpNormalize_8U_49U_else_lshift_1_rg_a = FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_7_FpNormalize_8U_49U_else_lshift_rg_a;
  assign nl_alu_loop_op_7_FpNormalize_8U_49U_else_lshift_rg_a = FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_8_FpNormalize_8U_49U_else_lshift_1_rg_a;
  assign nl_alu_loop_op_8_FpNormalize_8U_49U_else_lshift_1_rg_a = FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_9_FpNormalize_8U_49U_else_lshift_rg_a;
  assign nl_alu_loop_op_9_FpNormalize_8U_49U_else_lshift_rg_a = FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_10_FpNormalize_8U_49U_else_lshift_1_rg_a;
  assign nl_alu_loop_op_10_FpNormalize_8U_49U_else_lshift_1_rg_a = FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_11_FpNormalize_8U_49U_else_lshift_rg_a;
  assign nl_alu_loop_op_11_FpNormalize_8U_49U_else_lshift_rg_a = FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_12_FpNormalize_8U_49U_else_lshift_1_rg_a;
  assign nl_alu_loop_op_12_FpNormalize_8U_49U_else_lshift_1_rg_a = FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_13_FpNormalize_8U_49U_else_lshift_rg_a;
  assign nl_alu_loop_op_13_FpNormalize_8U_49U_else_lshift_rg_a = FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_14_FpNormalize_8U_49U_else_lshift_1_rg_a;
  assign nl_alu_loop_op_14_FpNormalize_8U_49U_else_lshift_1_rg_a = FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_15_FpNormalize_8U_49U_else_lshift_rg_a;
  assign nl_alu_loop_op_15_FpNormalize_8U_49U_else_lshift_rg_a = FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_16_FpNormalize_8U_49U_else_lshift_1_rg_a;
  assign nl_alu_loop_op_16_FpNormalize_8U_49U_else_lshift_1_rg_a = FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[48:0];
  wire [22:0] nl_alu_loop_op_1_leading_sign_23_0_rg_mantissa;
  assign nl_alu_loop_op_1_leading_sign_23_0_rg_mantissa = {alu_nan_to_zero_op_mant_1_lpi_1_dfm
      , 13'b0};
  wire [22:0] nl_alu_loop_op_2_leading_sign_23_0_1_rg_mantissa;
  assign nl_alu_loop_op_2_leading_sign_23_0_1_rg_mantissa = {alu_nan_to_zero_op_mant_2_lpi_1_dfm
      , 13'b0};
  wire [22:0] nl_alu_loop_op_3_leading_sign_23_0_rg_mantissa;
  assign nl_alu_loop_op_3_leading_sign_23_0_rg_mantissa = {alu_nan_to_zero_op_mant_3_lpi_1_dfm
      , 13'b0};
  wire [22:0] nl_alu_loop_op_4_leading_sign_23_0_1_rg_mantissa;
  assign nl_alu_loop_op_4_leading_sign_23_0_1_rg_mantissa = {alu_nan_to_zero_op_mant_4_lpi_1_dfm
      , 13'b0};
  wire [22:0] nl_alu_loop_op_5_leading_sign_23_0_rg_mantissa;
  assign nl_alu_loop_op_5_leading_sign_23_0_rg_mantissa = {alu_nan_to_zero_op_mant_5_lpi_1_dfm
      , 13'b0};
  wire [22:0] nl_alu_loop_op_6_leading_sign_23_0_1_rg_mantissa;
  assign nl_alu_loop_op_6_leading_sign_23_0_1_rg_mantissa = {alu_nan_to_zero_op_mant_6_lpi_1_dfm
      , 13'b0};
  wire [22:0] nl_alu_loop_op_7_leading_sign_23_0_rg_mantissa;
  assign nl_alu_loop_op_7_leading_sign_23_0_rg_mantissa = {alu_nan_to_zero_op_mant_7_lpi_1_dfm
      , 13'b0};
  wire [22:0] nl_alu_loop_op_8_leading_sign_23_0_1_rg_mantissa;
  assign nl_alu_loop_op_8_leading_sign_23_0_1_rg_mantissa = {alu_nan_to_zero_op_mant_8_lpi_1_dfm
      , 13'b0};
  wire [22:0] nl_alu_loop_op_9_leading_sign_23_0_rg_mantissa;
  assign nl_alu_loop_op_9_leading_sign_23_0_rg_mantissa = {alu_nan_to_zero_op_mant_9_lpi_1_dfm
      , 13'b0};
  wire [22:0] nl_alu_loop_op_10_leading_sign_23_0_1_rg_mantissa;
  assign nl_alu_loop_op_10_leading_sign_23_0_1_rg_mantissa = {alu_nan_to_zero_op_mant_10_lpi_1_dfm
      , 13'b0};
  wire [22:0] nl_alu_loop_op_11_leading_sign_23_0_rg_mantissa;
  assign nl_alu_loop_op_11_leading_sign_23_0_rg_mantissa = {alu_nan_to_zero_op_mant_11_lpi_1_dfm
      , 13'b0};
  wire [22:0] nl_alu_loop_op_12_leading_sign_23_0_1_rg_mantissa;
  assign nl_alu_loop_op_12_leading_sign_23_0_1_rg_mantissa = {alu_nan_to_zero_op_mant_12_lpi_1_dfm
      , 13'b0};
  wire [22:0] nl_alu_loop_op_13_leading_sign_23_0_rg_mantissa;
  assign nl_alu_loop_op_13_leading_sign_23_0_rg_mantissa = {alu_nan_to_zero_op_mant_13_lpi_1_dfm
      , 13'b0};
  wire [22:0] nl_alu_loop_op_14_leading_sign_23_0_1_rg_mantissa;
  assign nl_alu_loop_op_14_leading_sign_23_0_1_rg_mantissa = {alu_nan_to_zero_op_mant_14_lpi_1_dfm
      , 13'b0};
  wire [22:0] nl_alu_loop_op_15_leading_sign_23_0_rg_mantissa;
  assign nl_alu_loop_op_15_leading_sign_23_0_rg_mantissa = {alu_nan_to_zero_op_mant_15_lpi_1_dfm
      , 13'b0};
  wire [22:0] nl_alu_loop_op_16_leading_sign_23_0_1_rg_mantissa;
  assign nl_alu_loop_op_16_leading_sign_23_0_1_rg_mantissa = {alu_nan_to_zero_op_mant_lpi_1_dfm
      , 13'b0};
  wire [48:0] nl_alu_loop_op_1_leading_sign_49_0_rg_mantissa;
  assign nl_alu_loop_op_1_leading_sign_49_0_rg_mantissa = FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_mx2[48:0];
  wire [48:0] nl_alu_loop_op_2_leading_sign_49_0_1_rg_mantissa;
  assign nl_alu_loop_op_2_leading_sign_49_0_1_rg_mantissa = FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_mx2[48:0];
  wire [48:0] nl_alu_loop_op_3_leading_sign_49_0_rg_mantissa;
  assign nl_alu_loop_op_3_leading_sign_49_0_rg_mantissa = FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_mx2[48:0];
  wire [48:0] nl_alu_loop_op_4_leading_sign_49_0_1_rg_mantissa;
  assign nl_alu_loop_op_4_leading_sign_49_0_1_rg_mantissa = FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_mx2[48:0];
  wire [48:0] nl_alu_loop_op_5_leading_sign_49_0_rg_mantissa;
  assign nl_alu_loop_op_5_leading_sign_49_0_rg_mantissa = FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_mx2[48:0];
  wire [48:0] nl_alu_loop_op_6_leading_sign_49_0_1_rg_mantissa;
  assign nl_alu_loop_op_6_leading_sign_49_0_1_rg_mantissa = FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_mx2[48:0];
  wire [48:0] nl_alu_loop_op_7_leading_sign_49_0_rg_mantissa;
  assign nl_alu_loop_op_7_leading_sign_49_0_rg_mantissa = FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_mx2[48:0];
  wire [48:0] nl_alu_loop_op_8_leading_sign_49_0_1_rg_mantissa;
  assign nl_alu_loop_op_8_leading_sign_49_0_1_rg_mantissa = FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_mx2[48:0];
  wire [48:0] nl_alu_loop_op_9_leading_sign_49_0_rg_mantissa;
  assign nl_alu_loop_op_9_leading_sign_49_0_rg_mantissa = FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_mx2[48:0];
  wire [48:0] nl_alu_loop_op_10_leading_sign_49_0_1_rg_mantissa;
  assign nl_alu_loop_op_10_leading_sign_49_0_1_rg_mantissa = FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_mx2[48:0];
  wire [48:0] nl_alu_loop_op_11_leading_sign_49_0_rg_mantissa;
  assign nl_alu_loop_op_11_leading_sign_49_0_rg_mantissa = FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_mx2[48:0];
  wire [48:0] nl_alu_loop_op_12_leading_sign_49_0_1_rg_mantissa;
  assign nl_alu_loop_op_12_leading_sign_49_0_1_rg_mantissa = FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_mx2[48:0];
  wire [48:0] nl_alu_loop_op_13_leading_sign_49_0_rg_mantissa;
  assign nl_alu_loop_op_13_leading_sign_49_0_rg_mantissa = FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_mx2[48:0];
  wire [48:0] nl_alu_loop_op_14_leading_sign_49_0_1_rg_mantissa;
  assign nl_alu_loop_op_14_leading_sign_49_0_1_rg_mantissa = FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_mx2[48:0];
  wire [48:0] nl_alu_loop_op_15_leading_sign_49_0_rg_mantissa;
  assign nl_alu_loop_op_15_leading_sign_49_0_rg_mantissa = FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_mx2[48:0];
  wire [48:0] nl_alu_loop_op_16_leading_sign_49_0_1_rg_mantissa;
  assign nl_alu_loop_op_16_leading_sign_49_0_1_rg_mantissa = FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_mx2[48:0];
  wire [21:0] nl_alu_loop_op_1_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_alu_loop_op_1_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a = {(alu_nan_to_zero_op_mant_1_lpi_1_dfm[8:0])
      , 13'b0};
  wire [6:0] nl_alu_loop_op_1_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_alu_loop_op_1_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_16)
      + 6'b1;
  wire [21:0] nl_alu_loop_op_2_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a;
  assign nl_alu_loop_op_2_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a =
      {(alu_nan_to_zero_op_mant_2_lpi_1_dfm[8:0]) , 13'b0};
  wire [6:0] nl_alu_loop_op_2_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s;
  assign nl_alu_loop_op_2_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s =
      conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_17)
      + 6'b1;
  wire [21:0] nl_alu_loop_op_3_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_alu_loop_op_3_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a = {(alu_nan_to_zero_op_mant_3_lpi_1_dfm[8:0])
      , 13'b0};
  wire [6:0] nl_alu_loop_op_3_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_alu_loop_op_3_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_18)
      + 6'b1;
  wire [21:0] nl_alu_loop_op_4_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a;
  assign nl_alu_loop_op_4_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a =
      {(alu_nan_to_zero_op_mant_4_lpi_1_dfm[8:0]) , 13'b0};
  wire [6:0] nl_alu_loop_op_4_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s;
  assign nl_alu_loop_op_4_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s =
      conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_19)
      + 6'b1;
  wire [21:0] nl_alu_loop_op_5_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_alu_loop_op_5_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a = {(alu_nan_to_zero_op_mant_5_lpi_1_dfm[8:0])
      , 13'b0};
  wire [6:0] nl_alu_loop_op_5_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_alu_loop_op_5_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_20)
      + 6'b1;
  wire [21:0] nl_alu_loop_op_6_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a;
  assign nl_alu_loop_op_6_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a =
      {(alu_nan_to_zero_op_mant_6_lpi_1_dfm[8:0]) , 13'b0};
  wire [6:0] nl_alu_loop_op_6_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s;
  assign nl_alu_loop_op_6_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s =
      conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_21)
      + 6'b1;
  wire [21:0] nl_alu_loop_op_7_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_alu_loop_op_7_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a = {(alu_nan_to_zero_op_mant_7_lpi_1_dfm[8:0])
      , 13'b0};
  wire [6:0] nl_alu_loop_op_7_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_alu_loop_op_7_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_22)
      + 6'b1;
  wire [21:0] nl_alu_loop_op_8_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a;
  assign nl_alu_loop_op_8_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a =
      {(alu_nan_to_zero_op_mant_8_lpi_1_dfm[8:0]) , 13'b0};
  wire [6:0] nl_alu_loop_op_8_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s;
  assign nl_alu_loop_op_8_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s =
      conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_23)
      + 6'b1;
  wire [21:0] nl_alu_loop_op_9_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_alu_loop_op_9_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a = {(alu_nan_to_zero_op_mant_9_lpi_1_dfm[8:0])
      , 13'b0};
  wire [6:0] nl_alu_loop_op_9_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_alu_loop_op_9_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_24)
      + 6'b1;
  wire [21:0] nl_alu_loop_op_10_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a;
  assign nl_alu_loop_op_10_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a =
      {(alu_nan_to_zero_op_mant_10_lpi_1_dfm[8:0]) , 13'b0};
  wire [6:0] nl_alu_loop_op_10_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s;
  assign nl_alu_loop_op_10_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s =
      conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_25)
      + 6'b1;
  wire [21:0] nl_alu_loop_op_11_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_alu_loop_op_11_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a = {(alu_nan_to_zero_op_mant_11_lpi_1_dfm[8:0])
      , 13'b0};
  wire [6:0] nl_alu_loop_op_11_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_alu_loop_op_11_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_26)
      + 6'b1;
  wire [21:0] nl_alu_loop_op_12_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a;
  assign nl_alu_loop_op_12_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a =
      {(alu_nan_to_zero_op_mant_12_lpi_1_dfm[8:0]) , 13'b0};
  wire [6:0] nl_alu_loop_op_12_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s;
  assign nl_alu_loop_op_12_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s =
      conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_27)
      + 6'b1;
  wire [21:0] nl_alu_loop_op_13_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_alu_loop_op_13_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a = {(alu_nan_to_zero_op_mant_13_lpi_1_dfm[8:0])
      , 13'b0};
  wire [6:0] nl_alu_loop_op_13_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_alu_loop_op_13_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_28)
      + 6'b1;
  wire [21:0] nl_alu_loop_op_14_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a;
  assign nl_alu_loop_op_14_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a =
      {(alu_nan_to_zero_op_mant_14_lpi_1_dfm[8:0]) , 13'b0};
  wire [6:0] nl_alu_loop_op_14_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s;
  assign nl_alu_loop_op_14_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s =
      conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_29)
      + 6'b1;
  wire [21:0] nl_alu_loop_op_15_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_alu_loop_op_15_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a = {(alu_nan_to_zero_op_mant_15_lpi_1_dfm[8:0])
      , 13'b0};
  wire [6:0] nl_alu_loop_op_15_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_alu_loop_op_15_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_30)
      + 6'b1;
  wire [21:0] nl_alu_loop_op_16_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a;
  assign nl_alu_loop_op_16_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a =
      {(alu_nan_to_zero_op_mant_lpi_1_dfm[8:0]) , 13'b0};
  wire [6:0] nl_alu_loop_op_16_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s;
  assign nl_alu_loop_op_16_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s =
      conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_31)
      + 6'b1;
  wire [15:0] nl_alu_loop_op_16_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a;
  assign nl_alu_loop_op_16_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a = {else_AluOp_data_15_15_lpi_1_dfm_mx0
      , else_AluOp_data_15_14_10_lpi_1_dfm_mx0 , else_AluOp_data_15_9_0_lpi_1_dfm_mx0};
  wire [15:0] nl_alu_loop_op_15_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a;
  assign nl_alu_loop_op_15_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a = {else_AluOp_data_14_15_lpi_1_dfm_mx0
      , else_AluOp_data_14_14_10_lpi_1_dfm_mx0 , else_AluOp_data_14_9_0_lpi_1_dfm_mx0};
  wire [15:0] nl_alu_loop_op_14_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a;
  assign nl_alu_loop_op_14_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a = {else_AluOp_data_13_15_lpi_1_dfm_mx0
      , else_AluOp_data_13_14_10_lpi_1_dfm_mx0 , else_AluOp_data_13_9_0_lpi_1_dfm_mx0};
  wire [15:0] nl_alu_loop_op_13_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a;
  assign nl_alu_loop_op_13_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a = {else_AluOp_data_12_15_lpi_1_dfm_mx0
      , else_AluOp_data_12_14_10_lpi_1_dfm_mx0 , else_AluOp_data_12_9_0_lpi_1_dfm_mx0};
  wire [15:0] nl_alu_loop_op_12_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a;
  assign nl_alu_loop_op_12_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a = {else_AluOp_data_11_15_lpi_1_dfm_mx0
      , else_AluOp_data_11_14_10_lpi_1_dfm_mx0 , else_AluOp_data_11_9_0_lpi_1_dfm_mx0};
  wire [15:0] nl_alu_loop_op_11_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a;
  assign nl_alu_loop_op_11_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a = {else_AluOp_data_10_15_lpi_1_dfm_mx0
      , else_AluOp_data_10_14_10_lpi_1_dfm_mx0 , else_AluOp_data_10_9_0_lpi_1_dfm_mx0};
  wire [15:0] nl_alu_loop_op_10_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a;
  assign nl_alu_loop_op_10_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a = {else_AluOp_data_9_15_lpi_1_dfm_mx0
      , else_AluOp_data_9_14_10_lpi_1_dfm_mx0 , else_AluOp_data_9_9_0_lpi_1_dfm_mx0};
  wire [15:0] nl_alu_loop_op_9_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a;
  assign nl_alu_loop_op_9_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a = {else_AluOp_data_8_15_lpi_1_dfm_mx0
      , else_AluOp_data_8_14_10_lpi_1_dfm_mx0 , else_AluOp_data_8_9_0_lpi_1_dfm_mx0};
  wire [15:0] nl_alu_loop_op_8_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a;
  assign nl_alu_loop_op_8_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a = {else_AluOp_data_7_15_lpi_1_dfm_mx0
      , else_AluOp_data_7_14_10_lpi_1_dfm_mx0 , else_AluOp_data_7_9_0_lpi_1_dfm_mx0};
  wire [15:0] nl_alu_loop_op_7_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a;
  assign nl_alu_loop_op_7_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a = {else_AluOp_data_6_15_lpi_1_dfm_mx0
      , else_AluOp_data_6_14_10_lpi_1_dfm_mx0 , else_AluOp_data_6_9_0_lpi_1_dfm_mx0};
  wire [15:0] nl_alu_loop_op_6_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a;
  assign nl_alu_loop_op_6_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a = {else_AluOp_data_5_15_lpi_1_dfm_mx0
      , else_AluOp_data_5_14_10_lpi_1_dfm_mx0 , else_AluOp_data_5_9_0_lpi_1_dfm_mx0};
  wire [15:0] nl_alu_loop_op_5_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a;
  assign nl_alu_loop_op_5_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a = {else_AluOp_data_4_15_lpi_1_dfm_mx0
      , else_AluOp_data_4_14_10_lpi_1_dfm_mx0 , else_AluOp_data_4_9_0_lpi_1_dfm_mx0};
  wire [15:0] nl_alu_loop_op_4_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a;
  assign nl_alu_loop_op_4_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a = {else_AluOp_data_3_15_lpi_1_dfm_mx0
      , else_AluOp_data_3_14_10_lpi_1_dfm_mx0 , else_AluOp_data_3_9_0_lpi_1_dfm_mx0};
  wire [15:0] nl_alu_loop_op_3_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a;
  assign nl_alu_loop_op_3_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a = {else_AluOp_data_2_15_lpi_1_dfm_mx0
      , else_AluOp_data_2_14_10_lpi_1_dfm_mx0 , else_AluOp_data_2_9_0_lpi_1_dfm_mx0};
  wire [15:0] nl_alu_loop_op_2_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a;
  assign nl_alu_loop_op_2_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a = {else_AluOp_data_1_15_lpi_1_dfm_mx0
      , else_AluOp_data_1_14_10_lpi_1_dfm_mx0 , else_AluOp_data_1_9_0_lpi_1_dfm_mx0};
  wire [15:0] nl_alu_loop_op_1_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a;
  assign nl_alu_loop_op_1_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a = {else_AluOp_data_0_15_lpi_1_dfm_mx0
      , else_AluOp_data_0_14_10_lpi_1_dfm_mx0 , else_AluOp_data_0_9_0_lpi_1_dfm_mx0};
  wire [527:0] nl_X_alu_core_chn_alu_out_rsci_inst_chn_alu_out_rsci_d;
  assign nl_X_alu_core_chn_alu_out_rsci_inst_chn_alu_out_rsci_d = {chn_alu_out_rsci_d_527_526
      , chn_alu_out_rsci_d_525_522 , chn_alu_out_rsci_d_521_518 , chn_alu_out_rsci_d_517_496
      , chn_alu_out_rsci_d_495 , chn_alu_out_rsci_d_494_493 , chn_alu_out_rsci_d_492_489
      , chn_alu_out_rsci_d_488_485 , chn_alu_out_rsci_d_484_463 , chn_alu_out_rsci_d_462
      , chn_alu_out_rsci_d_461_460 , chn_alu_out_rsci_d_459_456 , chn_alu_out_rsci_d_455_452
      , chn_alu_out_rsci_d_451_430 , chn_alu_out_rsci_d_429 , chn_alu_out_rsci_d_428_427
      , chn_alu_out_rsci_d_426_423 , chn_alu_out_rsci_d_422_419 , chn_alu_out_rsci_d_418_397
      , chn_alu_out_rsci_d_396 , chn_alu_out_rsci_d_395_394 , chn_alu_out_rsci_d_393_390
      , chn_alu_out_rsci_d_389_386 , chn_alu_out_rsci_d_385_364 , chn_alu_out_rsci_d_363
      , chn_alu_out_rsci_d_362_361 , chn_alu_out_rsci_d_360_357 , chn_alu_out_rsci_d_356_353
      , chn_alu_out_rsci_d_352_331 , chn_alu_out_rsci_d_330 , chn_alu_out_rsci_d_329_328
      , chn_alu_out_rsci_d_327_324 , chn_alu_out_rsci_d_323_320 , chn_alu_out_rsci_d_319_298
      , chn_alu_out_rsci_d_297 , chn_alu_out_rsci_d_296_295 , chn_alu_out_rsci_d_294_291
      , chn_alu_out_rsci_d_290_287 , chn_alu_out_rsci_d_286_265 , chn_alu_out_rsci_d_264
      , chn_alu_out_rsci_d_263_262 , chn_alu_out_rsci_d_261_258 , chn_alu_out_rsci_d_257_254
      , chn_alu_out_rsci_d_253_232 , chn_alu_out_rsci_d_231 , chn_alu_out_rsci_d_230_229
      , chn_alu_out_rsci_d_228_225 , chn_alu_out_rsci_d_224_221 , chn_alu_out_rsci_d_220_199
      , chn_alu_out_rsci_d_198 , chn_alu_out_rsci_d_197_196 , chn_alu_out_rsci_d_195_192
      , chn_alu_out_rsci_d_191_188 , chn_alu_out_rsci_d_187_166 , chn_alu_out_rsci_d_165
      , chn_alu_out_rsci_d_164_163 , chn_alu_out_rsci_d_162_159 , chn_alu_out_rsci_d_158_155
      , chn_alu_out_rsci_d_154_133 , chn_alu_out_rsci_d_132 , chn_alu_out_rsci_d_131_130
      , chn_alu_out_rsci_d_129_126 , chn_alu_out_rsci_d_125_122 , chn_alu_out_rsci_d_121_100
      , chn_alu_out_rsci_d_99 , chn_alu_out_rsci_d_98_97 , chn_alu_out_rsci_d_96_93
      , chn_alu_out_rsci_d_92_89 , chn_alu_out_rsci_d_88_67 , chn_alu_out_rsci_d_66
      , chn_alu_out_rsci_d_65_64 , chn_alu_out_rsci_d_63_60 , chn_alu_out_rsci_d_59_56
      , chn_alu_out_rsci_d_55_34 , chn_alu_out_rsci_d_33 , chn_alu_out_rsci_d_32_31
      , chn_alu_out_rsci_d_30_27 , chn_alu_out_rsci_d_26_23 , chn_alu_out_rsci_d_22_1
      , chn_alu_out_rsci_d_0};
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
      .a(nl_alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_91_mx0w1)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
      .a(nl_alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_1_sva)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg (
      .a(nl_alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a[23:0]),
      .s(nl_alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_85_mx0w1)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg (
      .a(nl_alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a[23:0]),
      .s(nl_alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_2_sva)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
      .a(nl_alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_79_mx0w1)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
      .a(nl_alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_3_sva)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg (
      .a(nl_alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a[23:0]),
      .s(nl_alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_73_mx0w1)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg (
      .a(nl_alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a[23:0]),
      .s(nl_alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_4_sva)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_5_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
      .a(nl_alu_loop_op_5_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_alu_loop_op_5_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_67_mx0w1)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_5_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
      .a(nl_alu_loop_op_5_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_alu_loop_op_5_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_5_sva)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_6_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg (
      .a(nl_alu_loop_op_6_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a[23:0]),
      .s(nl_alu_loop_op_6_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_61_mx0w1)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_6_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg (
      .a(nl_alu_loop_op_6_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a[23:0]),
      .s(nl_alu_loop_op_6_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_6_sva)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_7_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
      .a(nl_alu_loop_op_7_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_alu_loop_op_7_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_55_mx0w1)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_7_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
      .a(nl_alu_loop_op_7_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_alu_loop_op_7_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_7_sva)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_8_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg (
      .a(nl_alu_loop_op_8_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a[23:0]),
      .s(nl_alu_loop_op_8_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_49_mx0w1)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_8_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg (
      .a(nl_alu_loop_op_8_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a[23:0]),
      .s(nl_alu_loop_op_8_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_8_sva)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_9_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
      .a(nl_alu_loop_op_9_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_alu_loop_op_9_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_43_mx0w1)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_9_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
      .a(nl_alu_loop_op_9_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_alu_loop_op_9_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_9_sva)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_10_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg (
      .a(nl_alu_loop_op_10_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a[23:0]),
      .s(nl_alu_loop_op_10_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_37_mx0w1)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_10_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg (
      .a(nl_alu_loop_op_10_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a[23:0]),
      .s(nl_alu_loop_op_10_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_10_sva)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_11_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
      .a(nl_alu_loop_op_11_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_alu_loop_op_11_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_31_mx0w1)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_11_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
      .a(nl_alu_loop_op_11_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_alu_loop_op_11_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_11_sva)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_12_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg (
      .a(nl_alu_loop_op_12_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a[23:0]),
      .s(nl_alu_loop_op_12_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_25_mx0w1)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_12_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg (
      .a(nl_alu_loop_op_12_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a[23:0]),
      .s(nl_alu_loop_op_12_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_12_sva)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_13_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
      .a(nl_alu_loop_op_13_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_alu_loop_op_13_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_19_mx0w1)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_13_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
      .a(nl_alu_loop_op_13_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_alu_loop_op_13_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_13_sva)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_14_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg (
      .a(nl_alu_loop_op_14_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a[23:0]),
      .s(nl_alu_loop_op_14_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_13_mx0w1)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_14_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg (
      .a(nl_alu_loop_op_14_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a[23:0]),
      .s(nl_alu_loop_op_14_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_14_sva)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_15_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
      .a(nl_alu_loop_op_15_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_alu_loop_op_15_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_7_mx0w1)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_15_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
      .a(nl_alu_loop_op_15_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_alu_loop_op_15_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_15_sva)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_16_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg (
      .a(nl_alu_loop_op_16_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a[23:0]),
      .s(nl_alu_loop_op_16_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_1_mx0w1)
    );
  SDP_X_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_16_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg (
      .a(nl_alu_loop_op_16_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a[23:0]),
      .s(nl_alu_loop_op_16_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_sva)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) alu_loop_op_1_FpNormalize_8U_49U_else_lshift_rg (
      .a(nl_alu_loop_op_1_FpNormalize_8U_49U_else_lshift_rg_a[48:0]),
      .s(IntLeadZero_49U_leading_sign_49_0_rtn_1_sva_2),
      .z(alu_loop_op_1_FpNormalize_8U_49U_else_lshift_itm)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) alu_loop_op_2_FpNormalize_8U_49U_else_lshift_1_rg (
      .a(nl_alu_loop_op_2_FpNormalize_8U_49U_else_lshift_1_rg_a[48:0]),
      .s(IntLeadZero_49U_leading_sign_49_0_rtn_2_sva_2),
      .z(alu_loop_op_2_FpNormalize_8U_49U_else_lshift_1_itm)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) alu_loop_op_3_FpNormalize_8U_49U_else_lshift_rg (
      .a(nl_alu_loop_op_3_FpNormalize_8U_49U_else_lshift_rg_a[48:0]),
      .s(IntLeadZero_49U_leading_sign_49_0_rtn_3_sva_2),
      .z(alu_loop_op_3_FpNormalize_8U_49U_else_lshift_itm)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) alu_loop_op_4_FpNormalize_8U_49U_else_lshift_1_rg (
      .a(nl_alu_loop_op_4_FpNormalize_8U_49U_else_lshift_1_rg_a[48:0]),
      .s(IntLeadZero_49U_leading_sign_49_0_rtn_4_sva_2),
      .z(alu_loop_op_4_FpNormalize_8U_49U_else_lshift_1_itm)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) alu_loop_op_5_FpNormalize_8U_49U_else_lshift_rg (
      .a(nl_alu_loop_op_5_FpNormalize_8U_49U_else_lshift_rg_a[48:0]),
      .s(IntLeadZero_49U_leading_sign_49_0_rtn_5_sva_2),
      .z(alu_loop_op_5_FpNormalize_8U_49U_else_lshift_itm)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) alu_loop_op_6_FpNormalize_8U_49U_else_lshift_1_rg (
      .a(nl_alu_loop_op_6_FpNormalize_8U_49U_else_lshift_1_rg_a[48:0]),
      .s(IntLeadZero_49U_leading_sign_49_0_rtn_6_sva_2),
      .z(alu_loop_op_6_FpNormalize_8U_49U_else_lshift_1_itm)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) alu_loop_op_7_FpNormalize_8U_49U_else_lshift_rg (
      .a(nl_alu_loop_op_7_FpNormalize_8U_49U_else_lshift_rg_a[48:0]),
      .s(IntLeadZero_49U_leading_sign_49_0_rtn_7_sva_2),
      .z(alu_loop_op_7_FpNormalize_8U_49U_else_lshift_itm)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) alu_loop_op_8_FpNormalize_8U_49U_else_lshift_1_rg (
      .a(nl_alu_loop_op_8_FpNormalize_8U_49U_else_lshift_1_rg_a[48:0]),
      .s(IntLeadZero_49U_leading_sign_49_0_rtn_8_sva_2),
      .z(alu_loop_op_8_FpNormalize_8U_49U_else_lshift_1_itm)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) alu_loop_op_9_FpNormalize_8U_49U_else_lshift_rg (
      .a(nl_alu_loop_op_9_FpNormalize_8U_49U_else_lshift_rg_a[48:0]),
      .s(IntLeadZero_49U_leading_sign_49_0_rtn_9_sva_2),
      .z(alu_loop_op_9_FpNormalize_8U_49U_else_lshift_itm)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) alu_loop_op_10_FpNormalize_8U_49U_else_lshift_1_rg (
      .a(nl_alu_loop_op_10_FpNormalize_8U_49U_else_lshift_1_rg_a[48:0]),
      .s(IntLeadZero_49U_leading_sign_49_0_rtn_10_sva_2),
      .z(alu_loop_op_10_FpNormalize_8U_49U_else_lshift_1_itm)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) alu_loop_op_11_FpNormalize_8U_49U_else_lshift_rg (
      .a(nl_alu_loop_op_11_FpNormalize_8U_49U_else_lshift_rg_a[48:0]),
      .s(IntLeadZero_49U_leading_sign_49_0_rtn_11_sva_2),
      .z(alu_loop_op_11_FpNormalize_8U_49U_else_lshift_itm)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) alu_loop_op_12_FpNormalize_8U_49U_else_lshift_1_rg (
      .a(nl_alu_loop_op_12_FpNormalize_8U_49U_else_lshift_1_rg_a[48:0]),
      .s(IntLeadZero_49U_leading_sign_49_0_rtn_12_sva_2),
      .z(alu_loop_op_12_FpNormalize_8U_49U_else_lshift_1_itm)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) alu_loop_op_13_FpNormalize_8U_49U_else_lshift_rg (
      .a(nl_alu_loop_op_13_FpNormalize_8U_49U_else_lshift_rg_a[48:0]),
      .s(IntLeadZero_49U_leading_sign_49_0_rtn_13_sva_2),
      .z(alu_loop_op_13_FpNormalize_8U_49U_else_lshift_itm)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) alu_loop_op_14_FpNormalize_8U_49U_else_lshift_1_rg (
      .a(nl_alu_loop_op_14_FpNormalize_8U_49U_else_lshift_1_rg_a[48:0]),
      .s(IntLeadZero_49U_leading_sign_49_0_rtn_14_sva_2),
      .z(alu_loop_op_14_FpNormalize_8U_49U_else_lshift_1_itm)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) alu_loop_op_15_FpNormalize_8U_49U_else_lshift_rg (
      .a(nl_alu_loop_op_15_FpNormalize_8U_49U_else_lshift_rg_a[48:0]),
      .s(IntLeadZero_49U_leading_sign_49_0_rtn_15_sva_2),
      .z(alu_loop_op_15_FpNormalize_8U_49U_else_lshift_itm)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) alu_loop_op_16_FpNormalize_8U_49U_else_lshift_1_rg (
      .a(nl_alu_loop_op_16_FpNormalize_8U_49U_else_lshift_1_rg_a[48:0]),
      .s(IntLeadZero_49U_leading_sign_49_0_rtn_sva_2),
      .z(alu_loop_op_16_FpNormalize_8U_49U_else_lshift_1_itm)
    );
  SDP_X_leading_sign_23_0 alu_loop_op_1_leading_sign_23_0_rg (
      .mantissa(nl_alu_loop_op_1_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_16)
    );
  SDP_X_leading_sign_23_0 alu_loop_op_2_leading_sign_23_0_1_rg (
      .mantissa(nl_alu_loop_op_2_leading_sign_23_0_1_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_17)
    );
  SDP_X_leading_sign_23_0 alu_loop_op_3_leading_sign_23_0_rg (
      .mantissa(nl_alu_loop_op_3_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_18)
    );
  SDP_X_leading_sign_23_0 alu_loop_op_4_leading_sign_23_0_1_rg (
      .mantissa(nl_alu_loop_op_4_leading_sign_23_0_1_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_19)
    );
  SDP_X_leading_sign_23_0 alu_loop_op_5_leading_sign_23_0_rg (
      .mantissa(nl_alu_loop_op_5_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_20)
    );
  SDP_X_leading_sign_23_0 alu_loop_op_6_leading_sign_23_0_1_rg (
      .mantissa(nl_alu_loop_op_6_leading_sign_23_0_1_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_21)
    );
  SDP_X_leading_sign_23_0 alu_loop_op_7_leading_sign_23_0_rg (
      .mantissa(nl_alu_loop_op_7_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_22)
    );
  SDP_X_leading_sign_23_0 alu_loop_op_8_leading_sign_23_0_1_rg (
      .mantissa(nl_alu_loop_op_8_leading_sign_23_0_1_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_23)
    );
  SDP_X_leading_sign_23_0 alu_loop_op_9_leading_sign_23_0_rg (
      .mantissa(nl_alu_loop_op_9_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_24)
    );
  SDP_X_leading_sign_23_0 alu_loop_op_10_leading_sign_23_0_1_rg (
      .mantissa(nl_alu_loop_op_10_leading_sign_23_0_1_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_25)
    );
  SDP_X_leading_sign_23_0 alu_loop_op_11_leading_sign_23_0_rg (
      .mantissa(nl_alu_loop_op_11_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_26)
    );
  SDP_X_leading_sign_23_0 alu_loop_op_12_leading_sign_23_0_1_rg (
      .mantissa(nl_alu_loop_op_12_leading_sign_23_0_1_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_27)
    );
  SDP_X_leading_sign_23_0 alu_loop_op_13_leading_sign_23_0_rg (
      .mantissa(nl_alu_loop_op_13_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_28)
    );
  SDP_X_leading_sign_23_0 alu_loop_op_14_leading_sign_23_0_1_rg (
      .mantissa(nl_alu_loop_op_14_leading_sign_23_0_1_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_29)
    );
  SDP_X_leading_sign_23_0 alu_loop_op_15_leading_sign_23_0_rg (
      .mantissa(nl_alu_loop_op_15_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_30)
    );
  SDP_X_leading_sign_23_0 alu_loop_op_16_leading_sign_23_0_1_rg (
      .mantissa(nl_alu_loop_op_16_leading_sign_23_0_1_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_31)
    );
  SDP_X_leading_sign_49_0 alu_loop_op_1_leading_sign_49_0_rg (
      .mantissa(nl_alu_loop_op_1_leading_sign_49_0_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_16)
    );
  SDP_X_leading_sign_49_0 alu_loop_op_2_leading_sign_49_0_1_rg (
      .mantissa(nl_alu_loop_op_2_leading_sign_49_0_1_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_17)
    );
  SDP_X_leading_sign_49_0 alu_loop_op_3_leading_sign_49_0_rg (
      .mantissa(nl_alu_loop_op_3_leading_sign_49_0_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_18)
    );
  SDP_X_leading_sign_49_0 alu_loop_op_4_leading_sign_49_0_1_rg (
      .mantissa(nl_alu_loop_op_4_leading_sign_49_0_1_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_19)
    );
  SDP_X_leading_sign_49_0 alu_loop_op_5_leading_sign_49_0_rg (
      .mantissa(nl_alu_loop_op_5_leading_sign_49_0_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_20)
    );
  SDP_X_leading_sign_49_0 alu_loop_op_6_leading_sign_49_0_1_rg (
      .mantissa(nl_alu_loop_op_6_leading_sign_49_0_1_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_21)
    );
  SDP_X_leading_sign_49_0 alu_loop_op_7_leading_sign_49_0_rg (
      .mantissa(nl_alu_loop_op_7_leading_sign_49_0_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_22)
    );
  SDP_X_leading_sign_49_0 alu_loop_op_8_leading_sign_49_0_1_rg (
      .mantissa(nl_alu_loop_op_8_leading_sign_49_0_1_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_23)
    );
  SDP_X_leading_sign_49_0 alu_loop_op_9_leading_sign_49_0_rg (
      .mantissa(nl_alu_loop_op_9_leading_sign_49_0_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_24)
    );
  SDP_X_leading_sign_49_0 alu_loop_op_10_leading_sign_49_0_1_rg (
      .mantissa(nl_alu_loop_op_10_leading_sign_49_0_1_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_25)
    );
  SDP_X_leading_sign_49_0 alu_loop_op_11_leading_sign_49_0_rg (
      .mantissa(nl_alu_loop_op_11_leading_sign_49_0_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_26)
    );
  SDP_X_leading_sign_49_0 alu_loop_op_12_leading_sign_49_0_1_rg (
      .mantissa(nl_alu_loop_op_12_leading_sign_49_0_1_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_27)
    );
  SDP_X_leading_sign_49_0 alu_loop_op_13_leading_sign_49_0_rg (
      .mantissa(nl_alu_loop_op_13_leading_sign_49_0_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_28)
    );
  SDP_X_leading_sign_49_0 alu_loop_op_14_leading_sign_49_0_1_rg (
      .mantissa(nl_alu_loop_op_14_leading_sign_49_0_1_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_29)
    );
  SDP_X_leading_sign_49_0 alu_loop_op_15_leading_sign_49_0_rg (
      .mantissa(nl_alu_loop_op_15_leading_sign_49_0_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_30)
    );
  SDP_X_leading_sign_49_0 alu_loop_op_16_leading_sign_49_0_1_rg (
      .mantissa(nl_alu_loop_op_16_leading_sign_49_0_1_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_31)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) alu_loop_op_1_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_alu_loop_op_1_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_alu_loop_op_1_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_sva_2)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) alu_loop_op_2_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg
      (
      .a(nl_alu_loop_op_2_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a[21:0]),
      .s(nl_alu_loop_op_2_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_sva_2)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) alu_loop_op_3_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_alu_loop_op_3_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_alu_loop_op_3_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_sva_2)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) alu_loop_op_4_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg
      (
      .a(nl_alu_loop_op_4_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a[21:0]),
      .s(nl_alu_loop_op_4_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_sva_2)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) alu_loop_op_5_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_alu_loop_op_5_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_alu_loop_op_5_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_sva_2)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) alu_loop_op_6_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg
      (
      .a(nl_alu_loop_op_6_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a[21:0]),
      .s(nl_alu_loop_op_6_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_sva_2)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) alu_loop_op_7_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_alu_loop_op_7_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_alu_loop_op_7_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_sva_2)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) alu_loop_op_8_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg
      (
      .a(nl_alu_loop_op_8_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a[21:0]),
      .s(nl_alu_loop_op_8_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_sva_2)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) alu_loop_op_9_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_alu_loop_op_9_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_alu_loop_op_9_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_sva_2)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) alu_loop_op_10_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg
      (
      .a(nl_alu_loop_op_10_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a[21:0]),
      .s(nl_alu_loop_op_10_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_sva_2)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) alu_loop_op_11_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_alu_loop_op_11_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_alu_loop_op_11_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_sva_2)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) alu_loop_op_12_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg
      (
      .a(nl_alu_loop_op_12_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a[21:0]),
      .s(nl_alu_loop_op_12_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_sva_2)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) alu_loop_op_13_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_alu_loop_op_13_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_alu_loop_op_13_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_sva_2)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) alu_loop_op_14_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg
      (
      .a(nl_alu_loop_op_14_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a[21:0]),
      .s(nl_alu_loop_op_14_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_sva_2)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) alu_loop_op_15_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_alu_loop_op_15_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_alu_loop_op_15_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_sva_2)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) alu_loop_op_16_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg
      (
      .a(nl_alu_loop_op_16_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_a[21:0]),
      .s(nl_alu_loop_op_16_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_1_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_sva_2)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd16),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd79)) alu_loop_op_16_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg
      (
      .a(nl_alu_loop_op_16_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a[15:0]),
      .s(cfg_alu_shift_value_1_sva_1),
      .z(IntShiftLeft_16U_6U_32U_mbits_fixed_sva)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd16),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd79)) alu_loop_op_15_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg
      (
      .a(nl_alu_loop_op_15_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a[15:0]),
      .s(cfg_alu_shift_value_1_sva_1),
      .z(IntShiftLeft_16U_6U_32U_mbits_fixed_15_sva)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd16),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd79)) alu_loop_op_14_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg
      (
      .a(nl_alu_loop_op_14_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a[15:0]),
      .s(cfg_alu_shift_value_1_sva_1),
      .z(IntShiftLeft_16U_6U_32U_mbits_fixed_14_sva)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd16),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd79)) alu_loop_op_13_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg
      (
      .a(nl_alu_loop_op_13_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a[15:0]),
      .s(cfg_alu_shift_value_1_sva_1),
      .z(IntShiftLeft_16U_6U_32U_mbits_fixed_13_sva)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd16),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd79)) alu_loop_op_12_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg
      (
      .a(nl_alu_loop_op_12_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a[15:0]),
      .s(cfg_alu_shift_value_1_sva_1),
      .z(IntShiftLeft_16U_6U_32U_mbits_fixed_12_sva)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd16),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd79)) alu_loop_op_11_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg
      (
      .a(nl_alu_loop_op_11_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a[15:0]),
      .s(cfg_alu_shift_value_1_sva_1),
      .z(IntShiftLeft_16U_6U_32U_mbits_fixed_11_sva)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd16),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd79)) alu_loop_op_10_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg
      (
      .a(nl_alu_loop_op_10_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a[15:0]),
      .s(cfg_alu_shift_value_1_sva_1),
      .z(IntShiftLeft_16U_6U_32U_mbits_fixed_10_sva)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd16),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd79)) alu_loop_op_9_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg
      (
      .a(nl_alu_loop_op_9_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a[15:0]),
      .s(cfg_alu_shift_value_1_sva_1),
      .z(IntShiftLeft_16U_6U_32U_mbits_fixed_9_sva)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd16),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd79)) alu_loop_op_8_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg
      (
      .a(nl_alu_loop_op_8_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a[15:0]),
      .s(cfg_alu_shift_value_1_sva_1),
      .z(IntShiftLeft_16U_6U_32U_mbits_fixed_8_sva)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd16),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd79)) alu_loop_op_7_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg
      (
      .a(nl_alu_loop_op_7_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a[15:0]),
      .s(cfg_alu_shift_value_1_sva_1),
      .z(IntShiftLeft_16U_6U_32U_mbits_fixed_7_sva)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd16),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd79)) alu_loop_op_6_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg
      (
      .a(nl_alu_loop_op_6_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a[15:0]),
      .s(cfg_alu_shift_value_1_sva_1),
      .z(IntShiftLeft_16U_6U_32U_mbits_fixed_6_sva)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd16),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd79)) alu_loop_op_5_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg
      (
      .a(nl_alu_loop_op_5_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a[15:0]),
      .s(cfg_alu_shift_value_1_sva_1),
      .z(IntShiftLeft_16U_6U_32U_mbits_fixed_5_sva)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd16),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd79)) alu_loop_op_4_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg
      (
      .a(nl_alu_loop_op_4_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a[15:0]),
      .s(cfg_alu_shift_value_1_sva_1),
      .z(IntShiftLeft_16U_6U_32U_mbits_fixed_4_sva)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd16),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd79)) alu_loop_op_3_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg
      (
      .a(nl_alu_loop_op_3_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a[15:0]),
      .s(cfg_alu_shift_value_1_sva_1),
      .z(IntShiftLeft_16U_6U_32U_mbits_fixed_3_sva)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd16),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd79)) alu_loop_op_2_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg
      (
      .a(nl_alu_loop_op_2_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_1_rg_a[15:0]),
      .s(cfg_alu_shift_value_1_sva_1),
      .z(IntShiftLeft_16U_6U_32U_mbits_fixed_2_sva)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd16),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd79)) alu_loop_op_1_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg
      (
      .a(nl_alu_loop_op_1_IntShiftLeft_16U_6U_32U_mbits_fixed_lshift_rg_a[15:0]),
      .s(cfg_alu_shift_value_1_sva_1),
      .z(IntShiftLeft_16U_6U_32U_mbits_fixed_1_sva)
    );
  SDP_X_X_alu_core_chn_alu_in_rsci X_alu_core_chn_alu_in_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_in_rsc_z(chn_alu_in_rsc_z),
      .chn_alu_in_rsc_vz(chn_alu_in_rsc_vz),
      .chn_alu_in_rsc_lz(chn_alu_in_rsc_lz),
      .chn_alu_in_rsci_oswt(chn_alu_in_rsci_oswt),
      .core_wen(core_wen),
      .chn_alu_in_rsci_iswt0(chn_alu_in_rsci_iswt0),
      .chn_alu_in_rsci_bawt(chn_alu_in_rsci_bawt),
      .chn_alu_in_rsci_wen_comp(chn_alu_in_rsci_wen_comp),
      .chn_alu_in_rsci_ld_core_psct(chn_alu_in_rsci_ld_core_psct),
      .chn_alu_in_rsci_d_mxwt(chn_alu_in_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  SDP_X_X_alu_core_chn_alu_op_rsci X_alu_core_chn_alu_op_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_op_rsc_z(chn_alu_op_rsc_z),
      .chn_alu_op_rsc_vz(chn_alu_op_rsc_vz),
      .chn_alu_op_rsc_lz(chn_alu_op_rsc_lz),
      .chn_alu_op_rsci_oswt(chn_alu_op_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_alu_op_rsci_iswt0(chn_alu_op_rsci_iswt0),
      .chn_alu_op_rsci_bawt(chn_alu_op_rsci_bawt),
      .chn_alu_op_rsci_wen_comp(chn_alu_op_rsci_wen_comp),
      .chn_alu_op_rsci_ld_core_psct(chn_alu_op_rsci_ld_core_psct),
      .chn_alu_op_rsci_d_mxwt(chn_alu_op_rsci_d_mxwt)
    );
  SDP_X_X_alu_core_chn_alu_out_rsci X_alu_core_chn_alu_out_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_out_rsc_z(chn_alu_out_rsc_z),
      .chn_alu_out_rsc_vz(chn_alu_out_rsc_vz),
      .chn_alu_out_rsc_lz(chn_alu_out_rsc_lz),
      .chn_alu_out_rsci_oswt(chn_alu_out_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_alu_out_rsci_iswt0(chn_alu_out_rsci_iswt0),
      .chn_alu_out_rsci_bawt(chn_alu_out_rsci_bawt),
      .chn_alu_out_rsci_wen_comp(chn_alu_out_rsci_wen_comp),
      .chn_alu_out_rsci_ld_core_psct(reg_chn_alu_out_rsci_ld_core_psct_cse),
      .chn_alu_out_rsci_d(nl_X_alu_core_chn_alu_out_rsci_inst_chn_alu_out_rsci_d[527:0])
    );
  SDP_X_X_alu_core_cfg_alu_op_rsc_triosy_obj X_alu_core_cfg_alu_op_rsc_triosy_obj_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_alu_op_rsc_triosy_lz(cfg_alu_op_rsc_triosy_lz),
      .cfg_alu_op_rsc_triosy_obj_oswt(cfg_alu_op_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_alu_op_rsc_triosy_obj_iswt0(reg_cfg_alu_shift_value_rsc_triosy_obj_ld_core_psct_cse),
      .cfg_alu_op_rsc_triosy_obj_bawt(cfg_alu_op_rsc_triosy_obj_bawt)
    );
  SDP_X_X_alu_core_cfg_alu_bypass_rsc_triosy_obj X_alu_core_cfg_alu_bypass_rsc_triosy_obj_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_alu_bypass_rsc_triosy_lz(cfg_alu_bypass_rsc_triosy_lz),
      .cfg_alu_bypass_rsc_triosy_obj_oswt(cfg_alu_bypass_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_alu_bypass_rsc_triosy_obj_iswt0(reg_cfg_alu_shift_value_rsc_triosy_obj_ld_core_psct_cse),
      .cfg_alu_bypass_rsc_triosy_obj_bawt(cfg_alu_bypass_rsc_triosy_obj_bawt)
    );
  SDP_X_X_alu_core_cfg_alu_algo_rsc_triosy_obj X_alu_core_cfg_alu_algo_rsc_triosy_obj_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_alu_algo_rsc_triosy_lz(cfg_alu_algo_rsc_triosy_lz),
      .cfg_alu_algo_rsc_triosy_obj_oswt(cfg_alu_algo_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_alu_algo_rsc_triosy_obj_iswt0(reg_cfg_alu_shift_value_rsc_triosy_obj_ld_core_psct_cse),
      .cfg_alu_algo_rsc_triosy_obj_bawt(cfg_alu_algo_rsc_triosy_obj_bawt)
    );
  SDP_X_X_alu_core_cfg_alu_src_rsc_triosy_obj X_alu_core_cfg_alu_src_rsc_triosy_obj_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_alu_src_rsc_triosy_lz(cfg_alu_src_rsc_triosy_lz),
      .cfg_alu_src_rsc_triosy_obj_oswt(cfg_alu_src_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_alu_src_rsc_triosy_obj_iswt0(reg_cfg_alu_shift_value_rsc_triosy_obj_ld_core_psct_cse),
      .cfg_alu_src_rsc_triosy_obj_bawt(cfg_alu_src_rsc_triosy_obj_bawt)
    );
  SDP_X_X_alu_core_cfg_alu_shift_value_rsc_triosy_obj X_alu_core_cfg_alu_shift_value_rsc_triosy_obj_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_alu_shift_value_rsc_triosy_lz(cfg_alu_shift_value_rsc_triosy_lz),
      .cfg_alu_shift_value_rsc_triosy_obj_oswt(cfg_alu_shift_value_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_alu_shift_value_rsc_triosy_obj_iswt0(reg_cfg_alu_shift_value_rsc_triosy_obj_ld_core_psct_cse),
      .cfg_alu_shift_value_rsc_triosy_obj_bawt(cfg_alu_shift_value_rsc_triosy_obj_bawt)
    );
  SDP_X_X_alu_core_staller X_alu_core_staller_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .chn_alu_in_rsci_wen_comp(chn_alu_in_rsci_wen_comp),
      .core_wten(core_wten),
      .chn_alu_op_rsci_wen_comp(chn_alu_op_rsci_wen_comp),
      .chn_alu_out_rsci_wen_comp(chn_alu_out_rsci_wen_comp)
    );
  SDP_X_X_alu_core_core_fsm X_alu_core_core_fsm_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign iExpoWidth_oExpoWidth_prb = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL alu_loop_op_1_X_alu_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL alu_loop_op_1_X_alu_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_1 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL alu_loop_op_1_X_alu_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_1 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_1 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL alu_loop_op_1_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_1 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_2 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL alu_loop_op_2_X_alu_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_2 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_2 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL alu_loop_op_2_X_alu_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_2 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_3 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL alu_loop_op_2_X_alu_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_3 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_3 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL alu_loop_op_2_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_3 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_4 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL alu_loop_op_3_X_alu_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_4 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_4 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL alu_loop_op_3_X_alu_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_4 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_5 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL alu_loop_op_3_X_alu_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_5 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_5 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL alu_loop_op_3_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_5 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_6 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL alu_loop_op_4_X_alu_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_6 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_6 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL alu_loop_op_4_X_alu_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_6 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_7 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL alu_loop_op_4_X_alu_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_7 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_7 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL alu_loop_op_4_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_7 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_8 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL alu_loop_op_5_X_alu_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_8 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_8 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL alu_loop_op_5_X_alu_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_8 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_9 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL alu_loop_op_5_X_alu_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_9 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_9 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL alu_loop_op_5_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_9 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_10 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL alu_loop_op_6_X_alu_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_10 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_10 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL alu_loop_op_6_X_alu_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_10 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_11 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL alu_loop_op_6_X_alu_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_11 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_11 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL alu_loop_op_6_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_11 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_12 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL alu_loop_op_7_X_alu_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_12 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_12 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL alu_loop_op_7_X_alu_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_12 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_13 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL alu_loop_op_7_X_alu_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_13 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_13 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL alu_loop_op_7_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_13 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_14 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL alu_loop_op_8_X_alu_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_14 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_14 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL alu_loop_op_8_X_alu_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_14 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_15 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL alu_loop_op_8_X_alu_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_15 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_15 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL alu_loop_op_8_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_15 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_16 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL alu_loop_op_9_X_alu_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_16 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_16 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL alu_loop_op_9_X_alu_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_16 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_17 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL alu_loop_op_9_X_alu_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_17 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_17 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL alu_loop_op_9_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_17 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_18 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL alu_loop_op_10_X_alu_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_18 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_18 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL alu_loop_op_10_X_alu_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_18 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_19 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL alu_loop_op_10_X_alu_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_19 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_19 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL alu_loop_op_10_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_19 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_20 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL alu_loop_op_11_X_alu_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_20 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_20 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL alu_loop_op_11_X_alu_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_20 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_21 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL alu_loop_op_11_X_alu_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_21 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_21 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL alu_loop_op_11_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_21 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_22 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL alu_loop_op_12_X_alu_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_22 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_22 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL alu_loop_op_12_X_alu_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_22 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_23 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL alu_loop_op_12_X_alu_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_23 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_23 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL alu_loop_op_12_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_23 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_24 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL alu_loop_op_13_X_alu_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_24 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_24 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL alu_loop_op_13_X_alu_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_24 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_25 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL alu_loop_op_13_X_alu_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_25 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_25 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL alu_loop_op_13_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_25 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_26 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL alu_loop_op_14_X_alu_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_26 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_26 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL alu_loop_op_14_X_alu_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_26 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_27 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL alu_loop_op_14_X_alu_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_27 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_27 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL alu_loop_op_14_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_27 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_28 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL alu_loop_op_15_X_alu_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_28 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_28 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL alu_loop_op_15_X_alu_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_28 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_29 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL alu_loop_op_15_X_alu_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_29 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_29 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL alu_loop_op_15_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_29 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_30 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL alu_loop_op_16_X_alu_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_30 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_30 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL alu_loop_op_16_X_alu_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_30 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_31 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL alu_loop_op_16_X_alu_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_31 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_31 = alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_31 } @rose(nvdla_core_clk);
  assign or_4809_cse = ((~(alu_loop_op_else_equal_tmp | alu_loop_op_else_nor_tmp_82))
      & and_1_m1c) | (alu_loop_op_else_equal_tmp & and_1_m1c);
  assign chn_alu_out_and_cse = core_wen & (~(and_dcpl_7 | (~ main_stage_v_4)));
  assign and_149_cse = FpAlu_8U_23U_nor_dfs_79 & nor_7_ssc;
  assign and_150_cse = FpAlu_8U_23U_equal_tmp_235 & nor_7_ssc;
  assign and_151_cse = FpAlu_8U_23U_equal_tmp_237 & nor_7_ssc;
  assign and_152_cse = FpAlu_8U_23U_equal_tmp_239 & nor_7_ssc;
  assign or_cse_2 = (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt;
  assign FpAlu_8U_23U_or_863_cse = (FpAdd_8U_23U_and_ssc & FpAlu_8U_23U_nor_dfs_79)
      | FpAlu_8U_23U_or_831_itm_4;
  assign FpAlu_8U_23U_or_864_cse = (FpAdd_8U_23U_and_2_ssc & FpAlu_8U_23U_nor_dfs_79)
      | FpAlu_8U_23U_or_833_itm_4;
  assign FpAlu_8U_23U_or_865_cse = (FpAdd_8U_23U_and_4_ssc & FpAlu_8U_23U_nor_dfs_79)
      | FpAlu_8U_23U_or_835_itm_4;
  assign FpAlu_8U_23U_or_866_cse = (FpAdd_8U_23U_and_6_ssc & FpAlu_8U_23U_nor_dfs_79)
      | FpAlu_8U_23U_or_837_itm_4;
  assign FpAlu_8U_23U_or_867_cse = (FpAdd_8U_23U_and_8_ssc & FpAlu_8U_23U_nor_dfs_79)
      | FpAlu_8U_23U_or_839_itm_4;
  assign FpAlu_8U_23U_or_868_cse = (FpAdd_8U_23U_and_10_ssc & FpAlu_8U_23U_nor_dfs_79)
      | FpAlu_8U_23U_or_841_itm_4;
  assign FpAlu_8U_23U_or_869_cse = (FpAdd_8U_23U_and_12_ssc & FpAlu_8U_23U_nor_dfs_79)
      | FpAlu_8U_23U_or_843_itm_4;
  assign FpAlu_8U_23U_or_870_cse = (FpAdd_8U_23U_and_14_ssc & FpAlu_8U_23U_nor_dfs_79)
      | FpAlu_8U_23U_or_845_itm_4;
  assign FpAlu_8U_23U_or_871_cse = (FpAdd_8U_23U_and_16_ssc & FpAlu_8U_23U_nor_dfs_79)
      | FpAlu_8U_23U_or_847_itm_4;
  assign FpAlu_8U_23U_or_872_cse = (FpAdd_8U_23U_and_18_ssc & FpAlu_8U_23U_nor_dfs_79)
      | FpAlu_8U_23U_or_849_itm_4;
  assign FpAlu_8U_23U_or_873_cse = (FpAdd_8U_23U_and_20_ssc & FpAlu_8U_23U_nor_dfs_79)
      | FpAlu_8U_23U_or_851_itm_4;
  assign FpAlu_8U_23U_or_874_cse = (FpAdd_8U_23U_and_22_ssc & FpAlu_8U_23U_nor_dfs_79)
      | FpAlu_8U_23U_or_853_itm_4;
  assign FpAlu_8U_23U_or_875_cse = (FpAdd_8U_23U_and_24_ssc & FpAlu_8U_23U_nor_dfs_79)
      | FpAlu_8U_23U_or_855_itm_4;
  assign FpAlu_8U_23U_or_876_cse = (FpAdd_8U_23U_and_26_ssc & FpAlu_8U_23U_nor_dfs_79)
      | FpAlu_8U_23U_or_857_itm_4;
  assign FpAlu_8U_23U_or_877_cse = (FpAdd_8U_23U_and_28_ssc & FpAlu_8U_23U_nor_dfs_79)
      | FpAlu_8U_23U_or_859_itm_4;
  assign FpAlu_8U_23U_or_878_cse = (FpAdd_8U_23U_and_30_ssc & FpAlu_8U_23U_nor_dfs_79)
      | FpAlu_8U_23U_or_861_itm_4;
  assign AluIn_data_and_1_cse = core_wen & and_89_tmp;
  assign FpAdd_8U_23U_is_a_greater_oelse_and_17_cse = core_wen & and_89_tmp & not_tmp_4;
  assign nor_2055_nl = ~(io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2)
      | (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt);
  assign mux_15_nl = MUX_s_1_2_2((nor_2055_nl), (~ io_read_cfg_alu_bypass_rsc_svs_st_1),
      and_89_tmp);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_cse = core_wen & (and_dcpl_29
      | and_dcpl_30) & (mux_15_nl);
  assign and_498_rgt = and_dcpl_21 & and_89_tmp & (~ (cfg_alu_algo_1_sva_st_92[1]));
  assign FpCmp_8U_23U_false_if_and_32_cse = core_wen & (and_498_rgt | and_dcpl_34
      | and_dcpl_36 | and_543_rgt) & (~ mux_16_itm);
  assign FpAdd_8U_23U_is_a_greater_oelse_FpAdd_8U_23U_is_a_greater_oelse_or_21_cse
      = and_dcpl_22 | and_dcpl_23;
  assign FpAdd_8U_23U_is_a_greater_and_17_cse = core_wen & FpAdd_8U_23U_is_a_greater_oelse_FpAdd_8U_23U_is_a_greater_oelse_or_21_cse
      & not_tmp_4;
  assign and_543_rgt = and_89_tmp & (cfg_alu_algo_1_sva_st_92==2'b10);
  assign and_589_rgt = and_dcpl_21 & and_dcpl_122;
  assign FpCmp_8U_23U_false_if_and_39_cse = core_wen & (and_589_rgt | and_dcpl_34
      | and_dcpl_127 | and_543_rgt) & (~ mux_16_itm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_75_cse = core_wen & and_89_tmp
      & (~ mux_127_itm);
  assign or_338_cse = (reg_cfg_alu_algo_1_sva_st_93_cse[0]) | or_tmp_327;
  assign mux_157_cse = MUX_s_1_2_2(mux_tmp_149, or_tmp_329, reg_cfg_alu_algo_1_sva_st_93_cse[0]);
  assign or_343_cse = (cfg_alu_algo_1_sva_st_204!=2'b10) | (~ reg_chn_alu_out_rsci_ld_core_psct_cse)
      | chn_alu_out_rsci_bawt | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign mux_158_nl = MUX_s_1_2_2(mux_157_cse, or_338_cse, or_334_cse);
  assign mux_159_nl = MUX_s_1_2_2(or_343_cse, (mux_158_nl), reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign FpAdd_8U_23U_is_addition_and_cse = core_wen & (~ and_dcpl_7) & (~ (mux_159_nl));
  assign IsZero_8U_23U_1_and_cse = core_wen & (~ and_dcpl_7) & not_tmp_79;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_cse = core_wen & (~ and_dcpl_7);
  assign FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse = (and_dcpl_21
      & or_cse_2) | and_dcpl_241;
  assign FpAdd_8U_23U_b_left_shift_and_32_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & not_tmp_79;
  assign AluIn_data_and_2_cse = core_wen & (~ and_dcpl_7) & mux_tmp_156;
  assign mux_164_nl = MUX_s_1_2_2(mux_tmp_149, or_tmp_327, or_334_cse);
  assign mux_165_nl = MUX_s_1_2_2((mux_164_nl), or_343_cse, or_350_cse);
  assign FpAdd_8U_23U_is_addition_and_33_cse = core_wen & (~ and_dcpl_7) & (~ (mux_165_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_78_cse = core_wen & (~ and_dcpl_7)
      & (~ mux_tmp_149);
  assign and_715_rgt = or_cse_2 & ((~ FpCmp_8U_23U_false_is_a_greater_lpi_1_dfm_7)
      | IsNaN_8U_23U_3_land_lpi_1_dfm_7) & (~ IsNaN_8U_23U_1_land_lpi_1_dfm_8);
  assign nor_1930_cse = ~((~ main_stage_v_3) | (~ FpAlu_8U_23U_equal_tmp_144) | io_read_cfg_alu_bypass_rsc_svs_st_6);
  assign nor_1931_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (~ FpAlu_8U_23U_equal_tmp_235));
  assign mux_250_cse = MUX_s_1_2_2((nor_1931_nl), nor_1930_cse, or_cse_2);
  assign and_719_rgt = ((~(FpCmp_8U_23U_false_is_a_greater_lpi_1_dfm_7 | IsNaN_8U_23U_3_land_lpi_1_dfm_7))
      | IsNaN_8U_23U_1_land_lpi_1_dfm_8) & or_cse_2;
  assign nor_1928_cse = ~((~ main_stage_v_3) | (~ FpAlu_8U_23U_equal_tmp_148) | io_read_cfg_alu_bypass_rsc_svs_st_6);
  assign nor_1929_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (~ FpAlu_8U_23U_equal_tmp_239));
  assign mux_251_cse = MUX_s_1_2_2((nor_1929_nl), nor_1928_cse, or_cse_2);
  assign and_723_rgt = and_dcpl_256 & (IsNaN_8U_23U_3_land_15_lpi_1_dfm_7 | (~ FpCmp_8U_23U_false_is_a_greater_15_lpi_1_dfm_7));
  assign and_726_rgt = ((~(IsNaN_8U_23U_3_land_15_lpi_1_dfm_7 | FpCmp_8U_23U_false_is_a_greater_15_lpi_1_dfm_7))
      | IsNaN_8U_23U_1_land_15_lpi_1_dfm_8) & or_cse_2;
  assign and_730_rgt = and_dcpl_263 & ((~ FpCmp_8U_23U_false_is_a_greater_14_lpi_1_dfm_7)
      | IsNaN_8U_23U_3_land_14_lpi_1_dfm_7);
  assign and_733_rgt = ((~(FpCmp_8U_23U_false_is_a_greater_14_lpi_1_dfm_7 | IsNaN_8U_23U_3_land_14_lpi_1_dfm_7))
      | IsNaN_8U_23U_2_land_14_lpi_1_dfm_8) & or_cse_2;
  assign and_737_rgt = or_cse_2 & ((~ FpCmp_8U_23U_false_is_a_greater_13_lpi_1_dfm_7)
      | IsNaN_8U_23U_3_land_13_lpi_1_dfm_7) & (~ IsNaN_8U_23U_2_land_13_lpi_1_dfm_8);
  assign and_741_rgt = ((~(FpCmp_8U_23U_false_is_a_greater_13_lpi_1_dfm_7 | IsNaN_8U_23U_3_land_13_lpi_1_dfm_7))
      | IsNaN_8U_23U_2_land_13_lpi_1_dfm_8) & or_cse_2;
  assign and_745_rgt = or_cse_2 & (IsNaN_8U_23U_3_land_12_lpi_1_dfm_7 | (~ FpCmp_8U_23U_false_is_a_greater_12_lpi_1_dfm_7))
      & (~ IsNaN_8U_23U_2_land_12_lpi_1_dfm_8);
  assign and_749_rgt = ((~(IsNaN_8U_23U_3_land_12_lpi_1_dfm_7 | FpCmp_8U_23U_false_is_a_greater_12_lpi_1_dfm_7))
      | IsNaN_8U_23U_2_land_12_lpi_1_dfm_8) & or_cse_2;
  assign and_753_rgt = or_cse_2 & ((~ FpCmp_8U_23U_false_is_a_greater_11_lpi_1_dfm_7)
      | IsNaN_8U_23U_3_land_11_lpi_1_dfm_7) & (~ IsNaN_8U_23U_2_land_11_lpi_1_dfm_8);
  assign and_757_rgt = ((~(FpCmp_8U_23U_false_is_a_greater_11_lpi_1_dfm_7 | IsNaN_8U_23U_3_land_11_lpi_1_dfm_7))
      | IsNaN_8U_23U_2_land_11_lpi_1_dfm_8) & or_cse_2;
  assign and_761_rgt = and_dcpl_294 & (IsNaN_8U_23U_3_land_10_lpi_1_dfm_7 | (~ FpCmp_8U_23U_false_is_a_greater_10_lpi_1_dfm_7));
  assign and_764_rgt = ((~(IsNaN_8U_23U_3_land_10_lpi_1_dfm_7 | FpCmp_8U_23U_false_is_a_greater_10_lpi_1_dfm_7))
      | IsNaN_8U_23U_2_land_10_lpi_1_dfm_8) & or_cse_2;
  assign and_768_rgt = or_cse_2 & ((~ FpCmp_8U_23U_false_is_a_greater_9_lpi_1_dfm_7)
      | IsNaN_8U_23U_3_land_9_lpi_1_dfm_7) & (~ IsNaN_8U_23U_2_land_9_lpi_1_dfm_8);
  assign and_772_rgt = ((~(FpCmp_8U_23U_false_is_a_greater_9_lpi_1_dfm_7 | IsNaN_8U_23U_3_land_9_lpi_1_dfm_7))
      | IsNaN_8U_23U_2_land_9_lpi_1_dfm_8) & or_cse_2;
  assign and_776_rgt = and_dcpl_309 & ((~ FpCmp_8U_23U_false_is_a_greater_8_lpi_1_dfm_7)
      | IsNaN_8U_23U_3_land_8_lpi_1_dfm_7);
  assign and_779_rgt = ((~(FpCmp_8U_23U_false_is_a_greater_8_lpi_1_dfm_7 | IsNaN_8U_23U_3_land_8_lpi_1_dfm_7))
      | IsNaN_8U_23U_1_land_8_lpi_1_dfm_8) & or_cse_2;
  assign and_783_rgt = and_dcpl_316 & (IsNaN_8U_23U_3_land_7_lpi_1_dfm_7 | (~ FpCmp_8U_23U_false_is_a_greater_7_lpi_1_dfm_7));
  assign and_786_rgt = ((~(IsNaN_8U_23U_3_land_7_lpi_1_dfm_7 | FpCmp_8U_23U_false_is_a_greater_7_lpi_1_dfm_7))
      | IsNaN_8U_23U_1_land_7_lpi_1_dfm_8) & or_cse_2;
  assign and_790_rgt = or_cse_2 & (IsNaN_8U_23U_3_land_6_lpi_1_dfm_7 | (~ FpCmp_8U_23U_false_is_a_greater_6_lpi_1_dfm_7))
      & (~ IsNaN_8U_23U_2_land_6_lpi_1_dfm_8);
  assign and_794_rgt = ((~(IsNaN_8U_23U_3_land_6_lpi_1_dfm_7 | FpCmp_8U_23U_false_is_a_greater_6_lpi_1_dfm_7))
      | IsNaN_8U_23U_2_land_6_lpi_1_dfm_8) & or_cse_2;
  assign and_798_rgt = or_cse_2 & (IsNaN_8U_23U_3_land_5_lpi_1_dfm_7 | (~ FpCmp_8U_23U_false_is_a_greater_5_lpi_1_dfm_7))
      & (~ IsNaN_8U_23U_2_land_5_lpi_1_dfm_8);
  assign and_802_rgt = ((~(IsNaN_8U_23U_3_land_5_lpi_1_dfm_7 | FpCmp_8U_23U_false_is_a_greater_5_lpi_1_dfm_7))
      | IsNaN_8U_23U_2_land_5_lpi_1_dfm_8) & or_cse_2;
  assign and_806_rgt = or_cse_2 & ((~ FpCmp_8U_23U_false_is_a_greater_4_lpi_1_dfm_7)
      | IsNaN_8U_23U_3_land_4_lpi_1_dfm_7) & (~ IsNaN_8U_23U_2_land_4_lpi_1_dfm_8);
  assign and_810_rgt = ((~(FpCmp_8U_23U_false_is_a_greater_4_lpi_1_dfm_7 | IsNaN_8U_23U_3_land_4_lpi_1_dfm_7))
      | IsNaN_8U_23U_2_land_4_lpi_1_dfm_8) & or_cse_2;
  assign and_814_rgt = and_dcpl_347 & (IsNaN_8U_23U_3_land_3_lpi_1_dfm_7 | (~ FpCmp_8U_23U_false_is_a_greater_3_lpi_1_dfm_7));
  assign and_817_rgt = ((~(IsNaN_8U_23U_3_land_3_lpi_1_dfm_7 | FpCmp_8U_23U_false_is_a_greater_3_lpi_1_dfm_7))
      | IsNaN_8U_23U_1_land_3_lpi_1_dfm_8) & or_cse_2;
  assign and_821_rgt = and_dcpl_354 & ((~ FpCmp_8U_23U_false_is_a_greater_2_lpi_1_dfm_7)
      | IsNaN_8U_23U_3_land_2_lpi_1_dfm_7);
  assign and_824_rgt = ((~(FpCmp_8U_23U_false_is_a_greater_2_lpi_1_dfm_7 | IsNaN_8U_23U_3_land_2_lpi_1_dfm_7))
      | IsNaN_8U_23U_2_land_2_lpi_1_dfm_8) & or_cse_2;
  assign and_828_rgt = and_dcpl_361 & (IsNaN_8U_23U_3_land_1_lpi_1_dfm_7 | (~ FpCmp_8U_23U_false_is_a_greater_1_lpi_1_dfm_7));
  assign and_831_rgt = ((~(IsNaN_8U_23U_3_land_1_lpi_1_dfm_7 | FpCmp_8U_23U_false_is_a_greater_1_lpi_1_dfm_7))
      | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8) & or_cse_2;
  assign nor_1867_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (((cfg_alu_algo_1_sva_7!=2'b01)) & alu_loop_op_else_nor_tmp_82));
  assign mux_285_cse = MUX_s_1_2_2((nor_1867_nl), nor_1862_cse, or_cse_2);
  assign alu_loop_op_else_else_if_and_57_cse = core_wen & (~ and_dcpl_7) & mux_285_cse;
  assign nor_1863_nl = ~((cfg_alu_algo_1_sva_6[0]) | (~ alu_loop_op_else_nor_tmp_81));
  assign mux_286_nl = MUX_s_1_2_2((nor_1863_nl), alu_loop_op_else_nor_tmp_81, cfg_alu_algo_1_sva_6[1]);
  assign nor_1862_cse = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (mux_286_nl));
  assign alu_loop_op_else_else_if_and_60_cse = core_wen & (and_dcpl_369 | and_dcpl_372
      | and_dcpl_375) & mux_285_cse;
  assign alu_loop_op_else_else_if_and_66_cse = core_wen & (and_dcpl_379 | and_dcpl_372
      | and_dcpl_375) & mux_285_cse;
  assign nor_1817_nl = ~(nor_2061_cse | io_read_cfg_alu_bypass_rsc_svs_st_6 | (~
      main_stage_v_3));
  assign mux_348_nl = MUX_s_1_2_2(main_stage_v_4, (~ or_1935_cse), or_cse_2);
  assign mux_349_nl = MUX_s_1_2_2((mux_348_nl), (nor_1817_nl), io_read_cfg_alu_bypass_rsc_svs_7);
  assign FpAlu_8U_23U_and_832_cse = core_wen & (~ and_dcpl_7) & (mux_349_nl);
  assign nor_1815_cse = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (~ alu_loop_op_else_nor_tmp_81));
  assign nor_1816_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (~ alu_loop_op_else_nor_tmp_82));
  assign mux_351_nl = MUX_s_1_2_2((nor_1816_nl), nor_1815_cse, or_cse_2);
  assign AluOut_data_and_cse = core_wen & (~ and_dcpl_7) & (mux_351_nl);
  assign nor_1813_cse = ~((~ main_stage_v_3) | (~ FpAlu_8U_23U_equal_tmp_146) | io_read_cfg_alu_bypass_rsc_svs_st_6);
  assign nor_1814_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (~ FpAlu_8U_23U_equal_tmp_237));
  assign mux_352_nl = MUX_s_1_2_2((nor_1814_nl), nor_1813_cse, or_cse_2);
  assign FpAlu_8U_23U_o_and_cse = core_wen & (~ and_dcpl_7) & (mux_352_nl);
  assign nor_1748_cse = ~((~ FpAlu_8U_23U_or_831_itm_3) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_326_cse = ~((cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_327_cse = ~((cfg_alu_algo_1_sva_st_205!=2'b10));
  assign nor_1743_cse = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1742_cse = ~((cfg_precision!=2'b10) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign and_3766_nl = (~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_st_2
      & (FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm[49]))) & alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm;
  assign mux_387_nl = MUX_s_1_2_2(nor_1743_cse, nor_1742_cse, and_3766_nl);
  assign nor_1744_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & (~(alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2
      & (~(((~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_2)
      | FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_st_3) & (FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49]))))))));
  assign mux_388_nl = MUX_s_1_2_2((nor_1744_nl), (mux_387_nl), or_cse_2);
  assign FpAdd_8U_23U_and_176_cse = core_wen & (~ and_dcpl_7) & (mux_388_nl);
  assign nor_333_cse = ~((cfg_precision!=2'b10));
  assign FpAdd_8U_23U_int_mant_p1_and_16_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (~ mux_393_itm);
  assign nor_1735_nl = ~(FpAdd_8U_23U_mux_2_tmp_49 | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1736_nl = ~(alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm
      | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign mux_394_nl = MUX_s_1_2_2((nor_1736_nl), (nor_1735_nl), nor_333_cse);
  assign nor_1737_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205!=2'b10) | alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2);
  assign mux_395_nl = MUX_s_1_2_2((nor_1737_nl), (mux_394_nl), or_cse_2);
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (mux_395_nl);
  assign nor_1733_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48) | (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_1_lpi_1_dfm_9 | IsNaN_8U_23U_3_land_1_lpi_1_dfm_7);
  assign nor_1734_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_1_lpi_1_dfm_10 | (cfg_alu_algo_1_sva_st_205!=2'b10)
      | (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_9) | IsNaN_8U_23U_land_1_lpi_1_dfm_st_5);
  assign mux_396_nl = MUX_s_1_2_2((nor_1734_nl), (nor_1733_nl), or_cse_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_80_ssc = core_wen & (~ and_dcpl_7)
      & (mux_396_nl);
  assign mux_398_nl = MUX_s_1_2_2(main_stage_v_4, main_stage_v_3, or_cse_2);
  assign AluIn_data_and_3_cse = core_wen & (~ and_dcpl_7) & (mux_398_nl);
  assign or_899_cse = (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7;
  assign nor_338_nl = ~((~ FpAlu_8U_23U_nor_dfs_79) | (cfg_alu_algo_1_sva_st_205!=2'b10));
  assign mux_401_nl = MUX_s_1_2_2(mux_tmp_392, mux_tmp_393, nor_338_nl);
  assign mux_402_nl = MUX_s_1_2_2(mux_tmp_393, (mux_401_nl), FpAlu_8U_23U_equal_tmp_237);
  assign mux_403_nl = MUX_s_1_2_2((mux_402_nl), mux_tmp_392, or_899_cse);
  assign IsNaN_8U_23U_aelse_and_cse = core_wen & (~ and_dcpl_7) & (~ (mux_403_nl));
  assign IsNaN_8U_23U_aelse_and_16_cse = core_wen & (~ and_dcpl_7) & (~ mux_393_itm);
  assign nor_1720_cse = ~((~ FpAlu_8U_23U_or_833_itm_3) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1724_cse = ~((~ FpAlu_8U_23U_or_833_itm_4) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign and_3763_nl = (~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_st_2
      & (FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm[49]))) & alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm;
  assign mux_410_nl = MUX_s_1_2_2(nor_1743_cse, nor_1742_cse, and_3763_nl);
  assign nor_1716_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & (~(alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2
      & (~(((~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_2)
      | FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_st_3) & (FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49]))))))));
  assign mux_411_nl = MUX_s_1_2_2((nor_1716_nl), (mux_410_nl), or_cse_2);
  assign FpAdd_8U_23U_and_178_cse = core_wen & (~ and_dcpl_7) & (mux_411_nl);
  assign FpAdd_8U_23U_int_mant_p1_and_17_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (~ mux_415_itm);
  assign nor_1708_nl = ~(FpAdd_8U_23U_mux_18_tmp_49 | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1709_nl = ~(alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm
      | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign mux_416_nl = MUX_s_1_2_2((nor_1709_nl), (nor_1708_nl), nor_333_cse);
  assign nor_1710_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205!=2'b10) | alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2);
  assign mux_417_nl = MUX_s_1_2_2((nor_1710_nl), (mux_416_nl), or_cse_2);
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_16_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (mux_417_nl);
  assign nor_1706_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48) | (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_2_lpi_1_dfm_9 | IsNaN_8U_23U_2_land_2_lpi_1_dfm_8);
  assign nor_1707_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_2_lpi_1_dfm_10 | (cfg_alu_algo_1_sva_st_205!=2'b10)
      | (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_9) | IsNaN_8U_23U_land_2_lpi_1_dfm_st_5);
  assign mux_418_nl = MUX_s_1_2_2((nor_1707_nl), (nor_1706_nl), or_cse_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_81_ssc = core_wen & (~ and_dcpl_7)
      & (mux_418_nl);
  assign IsNaN_8U_23U_aelse_and_18_cse = core_wen & (~ and_dcpl_7) & (~ mux_415_itm);
  assign nor_1693_cse = ~((~ FpAlu_8U_23U_or_835_itm_3) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1697_cse = ~((~ FpAlu_8U_23U_or_835_itm_4) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign and_3760_nl = (~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_st_2
      & (FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm[49]))) & alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm;
  assign mux_431_nl = MUX_s_1_2_2(nor_1743_cse, nor_1742_cse, and_3760_nl);
  assign nor_1689_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & (~(alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2
      & (~(((~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_2)
      | FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_st_3) & (FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49]))))))));
  assign mux_432_nl = MUX_s_1_2_2((nor_1689_nl), (mux_431_nl), or_cse_2);
  assign FpAdd_8U_23U_and_180_cse = core_wen & (~ and_dcpl_7) & (mux_432_nl);
  assign nor_1681_nl = ~(FpAdd_8U_23U_mux_34_tmp_49 | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1682_nl = ~(alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm
      | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign mux_437_nl = MUX_s_1_2_2((nor_1682_nl), (nor_1681_nl), nor_333_cse);
  assign nor_1683_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205!=2'b10) | alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2);
  assign mux_438_nl = MUX_s_1_2_2((nor_1683_nl), (mux_437_nl), or_cse_2);
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_17_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (mux_438_nl);
  assign nor_1679_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48) | (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_3_lpi_1_dfm_9 | IsNaN_8U_23U_3_land_3_lpi_1_dfm_7);
  assign nor_1680_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_3_lpi_1_dfm_10 | (cfg_alu_algo_1_sva_st_205!=2'b10)
      | (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_9) | IsNaN_8U_23U_land_3_lpi_1_dfm_st_5);
  assign mux_439_nl = MUX_s_1_2_2((nor_1680_nl), (nor_1679_nl), or_cse_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_82_ssc = core_wen & (~ and_dcpl_7)
      & (mux_439_nl);
  assign nor_1666_cse = ~((~ FpAlu_8U_23U_or_837_itm_3) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1670_cse = ~((~ FpAlu_8U_23U_or_837_itm_4) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign and_3757_nl = (~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_4_sva_st_2
      & (FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm[49]))) & alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm;
  assign mux_452_nl = MUX_s_1_2_2(nor_1743_cse, nor_1742_cse, and_3757_nl);
  assign nor_1662_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & (~(alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2
      & (~(((~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_4_sva_2)
      | FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_4_sva_st_3) & (FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_5[49]))))))));
  assign mux_453_nl = MUX_s_1_2_2((nor_1662_nl), (mux_452_nl), or_cse_2);
  assign FpAdd_8U_23U_and_182_cse = core_wen & (~ and_dcpl_7) & (mux_453_nl);
  assign nor_1654_nl = ~(FpAdd_8U_23U_mux_50_tmp_49 | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1655_nl = ~(alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm
      | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign mux_458_nl = MUX_s_1_2_2((nor_1655_nl), (nor_1654_nl), nor_333_cse);
  assign nor_1656_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205!=2'b10) | alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2);
  assign mux_459_nl = MUX_s_1_2_2((nor_1656_nl), (mux_458_nl), or_cse_2);
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_18_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (mux_459_nl);
  assign nor_1652_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48) | (~ IsNaN_8U_23U_1_land_4_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_4_lpi_1_dfm_9 | IsNaN_8U_23U_2_land_4_lpi_1_dfm_8);
  assign nor_1653_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_4_lpi_1_dfm_10 | (cfg_alu_algo_1_sva_st_205!=2'b10)
      | (~ IsNaN_8U_23U_1_land_4_lpi_1_dfm_9) | IsNaN_8U_23U_land_4_lpi_1_dfm_st_5);
  assign mux_460_nl = MUX_s_1_2_2((nor_1653_nl), (nor_1652_nl), or_cse_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_83_ssc = core_wen & (~ and_dcpl_7)
      & (mux_460_nl);
  assign nor_1639_cse = ~((~ FpAlu_8U_23U_or_839_itm_3) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1643_cse = ~((~ FpAlu_8U_23U_or_839_itm_4) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign and_3754_nl = (~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_5_sva_st_2
      & (FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm[49]))) & alu_loop_op_5_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm;
  assign mux_473_nl = MUX_s_1_2_2(nor_1743_cse, nor_1742_cse, and_3754_nl);
  assign nor_1635_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & (~(alu_loop_op_5_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2
      & (~(((~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_5_sva_2)
      | FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_5_sva_st_3) & (FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_5[49]))))))));
  assign mux_474_nl = MUX_s_1_2_2((nor_1635_nl), (mux_473_nl), or_cse_2);
  assign FpAdd_8U_23U_and_184_cse = core_wen & (~ and_dcpl_7) & (mux_474_nl);
  assign FpAdd_8U_23U_int_mant_p1_and_20_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (~ mux_478_itm);
  assign nor_1627_nl = ~(FpAdd_8U_23U_mux_66_tmp_49 | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1628_nl = ~(alu_loop_op_5_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm
      | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign mux_479_nl = MUX_s_1_2_2((nor_1628_nl), (nor_1627_nl), nor_333_cse);
  assign nor_1629_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205!=2'b10) | alu_loop_op_5_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2);
  assign mux_480_nl = MUX_s_1_2_2((nor_1629_nl), (mux_479_nl), or_cse_2);
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_19_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (mux_480_nl);
  assign nor_1625_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48) | (~ IsNaN_8U_23U_1_land_5_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_5_lpi_1_dfm_9 | IsNaN_8U_23U_2_land_5_lpi_1_dfm_8);
  assign nor_1626_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_5_lpi_1_dfm_10 | (cfg_alu_algo_1_sva_st_205!=2'b10)
      | (~ IsNaN_8U_23U_1_land_5_lpi_1_dfm_9) | IsNaN_8U_23U_land_5_lpi_1_dfm_st_5);
  assign mux_481_nl = MUX_s_1_2_2((nor_1626_nl), (nor_1625_nl), or_cse_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_84_ssc = core_wen & (~ and_dcpl_7)
      & (mux_481_nl);
  assign IsNaN_8U_23U_aelse_and_24_cse = core_wen & (~ and_dcpl_7) & (~ mux_478_itm);
  assign nor_1612_cse = ~((~ FpAlu_8U_23U_or_841_itm_3) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1616_cse = ~((~ FpAlu_8U_23U_or_841_itm_4) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign and_3751_nl = (~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_6_sva_st_2
      & (FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm[49]))) & alu_loop_op_6_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm;
  assign mux_494_nl = MUX_s_1_2_2(nor_1743_cse, nor_1742_cse, and_3751_nl);
  assign nor_1608_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & (~(alu_loop_op_6_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2
      & (~(((~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_6_sva_2)
      | FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_6_sva_st_3) & (FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_5[49]))))))));
  assign mux_495_nl = MUX_s_1_2_2((nor_1608_nl), (mux_494_nl), or_cse_2);
  assign FpAdd_8U_23U_and_186_cse = core_wen & (~ and_dcpl_7) & (mux_495_nl);
  assign nor_1600_nl = ~(FpAdd_8U_23U_mux_82_tmp_49 | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1601_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | alu_loop_op_6_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm);
  assign mux_500_nl = MUX_s_1_2_2((nor_1601_nl), (nor_1600_nl), nor_333_cse);
  assign nor_1602_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205!=2'b10) | alu_loop_op_6_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2);
  assign mux_501_nl = MUX_s_1_2_2((nor_1602_nl), (mux_500_nl), or_cse_2);
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_20_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (mux_501_nl);
  assign nor_1598_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48) | (~ IsNaN_8U_23U_1_land_6_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_6_lpi_1_dfm_9 | IsNaN_8U_23U_2_land_6_lpi_1_dfm_8);
  assign nor_1599_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_6_lpi_1_dfm_10 | (cfg_alu_algo_1_sva_st_205!=2'b10)
      | (~ IsNaN_8U_23U_1_land_6_lpi_1_dfm_9) | IsNaN_8U_23U_land_6_lpi_1_dfm_st_5);
  assign mux_502_nl = MUX_s_1_2_2((nor_1599_nl), (nor_1598_nl), or_cse_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_85_ssc = core_wen & (~ and_dcpl_7)
      & (mux_502_nl);
  assign nor_1585_cse = ~((~ FpAlu_8U_23U_or_843_itm_3) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1589_cse = ~((~ FpAlu_8U_23U_or_843_itm_4) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign and_3747_nl = nor_1743_cse & (~(alu_loop_op_7_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm
      & or_22_cse));
  assign and_3748_nl = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_7_sva_st_2
      & (FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm[49]);
  assign mux_515_nl = MUX_s_1_2_2((and_3747_nl), nor_1743_cse, and_3748_nl);
  assign nor_1581_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & (~(alu_loop_op_7_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2
      & (~(((~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_7_sva_2)
      | FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_7_sva_st_3) & (FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_5[49]))))))));
  assign mux_516_nl = MUX_s_1_2_2((nor_1581_nl), (mux_515_nl), or_cse_2);
  assign FpAdd_8U_23U_and_188_cse = core_wen & (~ and_dcpl_7) & (mux_516_nl);
  assign nor_1574_nl = ~(FpAdd_8U_23U_mux_98_tmp_49 | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1575_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | alu_loop_op_7_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm);
  assign mux_521_nl = MUX_s_1_2_2((nor_1575_nl), (nor_1574_nl), nor_333_cse);
  assign nor_1576_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205!=2'b10) | alu_loop_op_7_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2);
  assign mux_522_nl = MUX_s_1_2_2((nor_1576_nl), (mux_521_nl), or_cse_2);
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_21_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (mux_522_nl);
  assign nor_1572_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48) | (~ IsNaN_8U_23U_1_land_7_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_7_lpi_1_dfm_9 | IsNaN_8U_23U_3_land_7_lpi_1_dfm_7);
  assign nor_1573_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_7_lpi_1_dfm_10 | (cfg_alu_algo_1_sva_st_205!=2'b10)
      | (~ IsNaN_8U_23U_1_land_7_lpi_1_dfm_9) | IsNaN_8U_23U_land_7_lpi_1_dfm_st_5);
  assign mux_523_nl = MUX_s_1_2_2((nor_1573_nl), (nor_1572_nl), or_cse_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_86_ssc = core_wen & (~ and_dcpl_7)
      & (mux_523_nl);
  assign nor_1559_cse = ~((~ FpAlu_8U_23U_or_845_itm_3) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1563_cse = ~((~ FpAlu_8U_23U_or_845_itm_4) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign and_3743_nl = nor_1743_cse & (~(alu_loop_op_8_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm
      & or_22_cse));
  assign and_3744_nl = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_8_sva_st_2
      & (FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm[49]);
  assign mux_536_nl = MUX_s_1_2_2((and_3743_nl), nor_1743_cse, and_3744_nl);
  assign nor_1555_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & (~(alu_loop_op_8_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2
      & (~(((~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_8_sva_2)
      | FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_8_sva_st_3) & (FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_5[49]))))))));
  assign mux_537_nl = MUX_s_1_2_2((nor_1555_nl), (mux_536_nl), or_cse_2);
  assign FpAdd_8U_23U_and_190_cse = core_wen & (~ and_dcpl_7) & (mux_537_nl);
  assign nor_1548_nl = ~(FpAdd_8U_23U_mux_114_tmp_49 | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1549_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | alu_loop_op_8_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm);
  assign mux_542_nl = MUX_s_1_2_2((nor_1549_nl), (nor_1548_nl), nor_333_cse);
  assign nor_1550_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205!=2'b10) | alu_loop_op_8_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2);
  assign mux_543_nl = MUX_s_1_2_2((nor_1550_nl), (mux_542_nl), or_cse_2);
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_22_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (mux_543_nl);
  assign nor_1546_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48) | (~ IsNaN_8U_23U_1_land_8_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_8_lpi_1_dfm_9 | IsNaN_8U_23U_3_land_8_lpi_1_dfm_7);
  assign nor_1547_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_8_lpi_1_dfm_10 | (cfg_alu_algo_1_sva_st_205!=2'b10)
      | (~ IsNaN_8U_23U_1_land_8_lpi_1_dfm_9) | IsNaN_8U_23U_land_8_lpi_1_dfm_st_5);
  assign mux_544_nl = MUX_s_1_2_2((nor_1547_nl), (nor_1546_nl), or_cse_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_87_ssc = core_wen & (~ and_dcpl_7)
      & (mux_544_nl);
  assign nor_1533_cse = ~((~ FpAlu_8U_23U_or_847_itm_3) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1537_cse = ~((~ FpAlu_8U_23U_or_847_itm_4) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign and_3739_nl = nor_1743_cse & (~(alu_loop_op_9_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm
      & or_22_cse));
  assign and_3740_nl = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_9_sva_st_2
      & (FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm[49]);
  assign mux_557_nl = MUX_s_1_2_2((and_3739_nl), nor_1743_cse, and_3740_nl);
  assign nor_1529_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & (~(alu_loop_op_9_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2
      & (~(((~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_9_sva_2)
      | FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_9_sva_st_3) & (FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_5[49]))))))));
  assign mux_558_nl = MUX_s_1_2_2((nor_1529_nl), (mux_557_nl), or_cse_2);
  assign FpAdd_8U_23U_and_192_cse = core_wen & (~ and_dcpl_7) & (mux_558_nl);
  assign nor_1522_nl = ~(FpAdd_8U_23U_mux_130_tmp_49 | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1523_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | alu_loop_op_9_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm);
  assign mux_563_nl = MUX_s_1_2_2((nor_1523_nl), (nor_1522_nl), nor_333_cse);
  assign nor_1524_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205!=2'b10) | alu_loop_op_9_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2);
  assign mux_564_nl = MUX_s_1_2_2((nor_1524_nl), (mux_563_nl), or_cse_2);
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_23_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (mux_564_nl);
  assign nor_1520_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48) | (~ IsNaN_8U_23U_1_land_9_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_9_lpi_1_dfm_9 | IsNaN_8U_23U_2_land_9_lpi_1_dfm_8);
  assign nor_1521_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_9_lpi_1_dfm_10 | (cfg_alu_algo_1_sva_st_205!=2'b10)
      | (~ IsNaN_8U_23U_1_land_9_lpi_1_dfm_9) | IsNaN_8U_23U_land_9_lpi_1_dfm_st_5);
  assign mux_565_nl = MUX_s_1_2_2((nor_1521_nl), (nor_1520_nl), or_cse_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_88_ssc = core_wen & (~ and_dcpl_7)
      & (mux_565_nl);
  assign nor_1507_cse = ~((~ FpAlu_8U_23U_or_849_itm_3) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1511_cse = ~((~ FpAlu_8U_23U_or_849_itm_4) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign and_3735_nl = nor_1743_cse & (~(alu_loop_op_10_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm
      & or_22_cse));
  assign and_3736_nl = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_10_sva_st_2
      & (FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm[49]);
  assign mux_578_nl = MUX_s_1_2_2((and_3735_nl), nor_1743_cse, and_3736_nl);
  assign nor_1503_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & (~(alu_loop_op_10_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2
      & (~(((~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_10_sva_2)
      | FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_10_sva_st_3) &
      (FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_5[49]))))))));
  assign mux_579_nl = MUX_s_1_2_2((nor_1503_nl), (mux_578_nl), or_cse_2);
  assign FpAdd_8U_23U_and_194_cse = core_wen & (~ and_dcpl_7) & (mux_579_nl);
  assign nor_1496_nl = ~(FpAdd_8U_23U_mux_146_tmp_49 | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1497_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | alu_loop_op_10_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm);
  assign mux_584_nl = MUX_s_1_2_2((nor_1497_nl), (nor_1496_nl), nor_333_cse);
  assign nor_1498_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205!=2'b10) | alu_loop_op_10_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2);
  assign mux_585_nl = MUX_s_1_2_2((nor_1498_nl), (mux_584_nl), or_cse_2);
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_24_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (mux_585_nl);
  assign nor_1494_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48) | (~ IsNaN_8U_23U_1_land_10_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_10_lpi_1_dfm_9 | IsNaN_8U_23U_2_land_10_lpi_1_dfm_8);
  assign nor_1495_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_10_lpi_1_dfm_10 | (cfg_alu_algo_1_sva_st_205!=2'b10)
      | (~ IsNaN_8U_23U_1_land_10_lpi_1_dfm_9) | IsNaN_8U_23U_land_10_lpi_1_dfm_st_5);
  assign mux_586_nl = MUX_s_1_2_2((nor_1495_nl), (nor_1494_nl), or_cse_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_89_ssc = core_wen & (~ and_dcpl_7)
      & (mux_586_nl);
  assign nor_1481_cse = ~((~ FpAlu_8U_23U_or_851_itm_3) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1485_cse = ~((~ FpAlu_8U_23U_or_851_itm_4) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign and_3731_nl = nor_1743_cse & (~(alu_loop_op_11_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm
      & or_22_cse));
  assign and_3732_nl = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_11_sva_st_2
      & (FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm[49]);
  assign mux_599_nl = MUX_s_1_2_2((and_3731_nl), nor_1743_cse, and_3732_nl);
  assign nor_1477_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & (~(alu_loop_op_11_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2
      & (~(((~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_11_sva_2)
      | FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_11_sva_st_3) &
      (FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_5[49]))))))));
  assign mux_600_nl = MUX_s_1_2_2((nor_1477_nl), (mux_599_nl), or_cse_2);
  assign FpAdd_8U_23U_and_196_cse = core_wen & (~ and_dcpl_7) & (mux_600_nl);
  assign FpAdd_8U_23U_int_mant_p1_and_26_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (~ mux_604_itm);
  assign nor_1470_nl = ~(FpAdd_8U_23U_mux_162_tmp_49 | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1471_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | alu_loop_op_11_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm);
  assign mux_605_nl = MUX_s_1_2_2((nor_1471_nl), (nor_1470_nl), nor_333_cse);
  assign nor_1472_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205!=2'b10) | alu_loop_op_11_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2);
  assign mux_606_nl = MUX_s_1_2_2((nor_1472_nl), (mux_605_nl), or_cse_2);
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_25_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (mux_606_nl);
  assign nor_1468_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48) | (~ IsNaN_8U_23U_1_land_11_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_11_lpi_1_dfm_9 | IsNaN_8U_23U_2_land_11_lpi_1_dfm_8);
  assign nor_1469_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_11_lpi_1_dfm_10 | (cfg_alu_algo_1_sva_st_205!=2'b10)
      | (~ IsNaN_8U_23U_1_land_11_lpi_1_dfm_9) | IsNaN_8U_23U_land_11_lpi_1_dfm_st_5);
  assign mux_607_nl = MUX_s_1_2_2((nor_1469_nl), (nor_1468_nl), or_cse_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_90_ssc = core_wen & (~ and_dcpl_7)
      & (mux_607_nl);
  assign IsNaN_8U_23U_aelse_and_36_cse = core_wen & (~ and_dcpl_7) & (~ mux_604_itm);
  assign nor_1455_cse = ~((~ FpAlu_8U_23U_or_853_itm_3) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1459_cse = ~((~ FpAlu_8U_23U_or_853_itm_4) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign and_3727_nl = nor_1743_cse & (~(alu_loop_op_12_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm
      & or_22_cse));
  assign and_3728_nl = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_12_sva_st_2
      & (FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm[49]);
  assign mux_620_nl = MUX_s_1_2_2((and_3727_nl), nor_1743_cse, and_3728_nl);
  assign nor_1451_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & (~(alu_loop_op_12_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2
      & (~(((~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_12_sva_2)
      | FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_12_sva_st_3) &
      (FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_5[49]))))))));
  assign mux_621_nl = MUX_s_1_2_2((nor_1451_nl), (mux_620_nl), or_cse_2);
  assign FpAdd_8U_23U_and_198_cse = core_wen & (~ and_dcpl_7) & (mux_621_nl);
  assign nor_1444_nl = ~(FpAdd_8U_23U_mux_178_tmp_49 | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1445_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | alu_loop_op_12_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm);
  assign mux_626_nl = MUX_s_1_2_2((nor_1445_nl), (nor_1444_nl), nor_333_cse);
  assign nor_1446_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205!=2'b10) | alu_loop_op_12_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2);
  assign mux_627_nl = MUX_s_1_2_2((nor_1446_nl), (mux_626_nl), or_cse_2);
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_26_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (mux_627_nl);
  assign nor_1442_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48) | (~ IsNaN_8U_23U_1_land_12_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_12_lpi_1_dfm_9 | IsNaN_8U_23U_2_land_12_lpi_1_dfm_8);
  assign nor_1443_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_12_lpi_1_dfm_10 | (cfg_alu_algo_1_sva_st_205!=2'b10)
      | (~ IsNaN_8U_23U_1_land_12_lpi_1_dfm_9) | IsNaN_8U_23U_land_12_lpi_1_dfm_st_5);
  assign mux_628_nl = MUX_s_1_2_2((nor_1443_nl), (nor_1442_nl), or_cse_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_91_ssc = core_wen & (~ and_dcpl_7)
      & (mux_628_nl);
  assign nor_1429_cse = ~((~ FpAlu_8U_23U_or_855_itm_3) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1433_cse = ~((~ FpAlu_8U_23U_or_855_itm_4) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign and_3723_nl = nor_1743_cse & (~(alu_loop_op_13_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm
      & or_22_cse));
  assign and_3724_nl = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_13_sva_st_2
      & (FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm[49]);
  assign mux_641_nl = MUX_s_1_2_2((and_3723_nl), nor_1743_cse, and_3724_nl);
  assign nor_1425_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & (~(alu_loop_op_13_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2
      & (~(((~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_13_sva_2)
      | FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_13_sva_st_3) &
      (FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_5[49]))))))));
  assign mux_642_nl = MUX_s_1_2_2((nor_1425_nl), (mux_641_nl), or_cse_2);
  assign FpAdd_8U_23U_and_200_cse = core_wen & (~ and_dcpl_7) & (mux_642_nl);
  assign nor_1418_nl = ~(FpAdd_8U_23U_mux_194_tmp_49 | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1419_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | alu_loop_op_13_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm);
  assign mux_647_nl = MUX_s_1_2_2((nor_1419_nl), (nor_1418_nl), nor_333_cse);
  assign nor_1420_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205!=2'b10) | alu_loop_op_13_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2);
  assign mux_648_nl = MUX_s_1_2_2((nor_1420_nl), (mux_647_nl), or_cse_2);
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_27_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (mux_648_nl);
  assign nor_1416_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48) | (~ IsNaN_8U_23U_1_land_13_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_13_lpi_1_dfm_9 | IsNaN_8U_23U_2_land_13_lpi_1_dfm_8);
  assign nor_1417_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_13_lpi_1_dfm_10 | (cfg_alu_algo_1_sva_st_205!=2'b10)
      | (~ IsNaN_8U_23U_1_land_13_lpi_1_dfm_9) | IsNaN_8U_23U_land_13_lpi_1_dfm_st_5);
  assign mux_649_nl = MUX_s_1_2_2((nor_1417_nl), (nor_1416_nl), or_cse_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_92_ssc = core_wen & (~ and_dcpl_7)
      & (mux_649_nl);
  assign nor_1403_cse = ~((~ FpAlu_8U_23U_or_857_itm_3) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1407_cse = ~((~ FpAlu_8U_23U_or_857_itm_4) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign and_3719_nl = nor_1743_cse & (~(alu_loop_op_14_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm
      & or_22_cse));
  assign and_3720_nl = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_14_sva_st_2
      & (FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm[49]);
  assign mux_662_nl = MUX_s_1_2_2((and_3719_nl), nor_1743_cse, and_3720_nl);
  assign nor_1399_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & (~(alu_loop_op_14_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2
      & (~(((~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_14_sva_2)
      | FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_14_sva_st_3) &
      (FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_5[49]))))))));
  assign mux_663_nl = MUX_s_1_2_2((nor_1399_nl), (mux_662_nl), or_cse_2);
  assign FpAdd_8U_23U_and_202_cse = core_wen & (~ and_dcpl_7) & (mux_663_nl);
  assign nor_1392_nl = ~(FpAdd_8U_23U_mux_210_tmp_49 | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1393_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | alu_loop_op_14_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm);
  assign mux_668_nl = MUX_s_1_2_2((nor_1393_nl), (nor_1392_nl), nor_333_cse);
  assign nor_1394_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205!=2'b10) | alu_loop_op_14_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2);
  assign mux_669_nl = MUX_s_1_2_2((nor_1394_nl), (mux_668_nl), or_cse_2);
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_28_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (mux_669_nl);
  assign nor_1390_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48) | (~ IsNaN_8U_23U_1_land_14_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_14_lpi_1_dfm_9 | IsNaN_8U_23U_2_land_14_lpi_1_dfm_8);
  assign nor_1391_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_14_lpi_1_dfm_10 | (cfg_alu_algo_1_sva_st_205!=2'b10)
      | (~ IsNaN_8U_23U_1_land_14_lpi_1_dfm_9) | IsNaN_8U_23U_land_14_lpi_1_dfm_st_5);
  assign mux_670_nl = MUX_s_1_2_2((nor_1391_nl), (nor_1390_nl), or_cse_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_93_ssc = core_wen & (~ and_dcpl_7)
      & (mux_670_nl);
  assign nor_1378_cse = ~((~ FpAlu_8U_23U_or_859_itm_3) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign and_3715_nl = nor_1743_cse & (~(alu_loop_op_15_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm
      & or_22_cse));
  assign and_3716_nl = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_15_sva_st_2
      & (FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm[49]);
  assign mux_682_nl = MUX_s_1_2_2((and_3715_nl), nor_1743_cse, and_3716_nl);
  assign nor_1374_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & (~(alu_loop_op_15_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2
      & (~(((~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_15_sva_2)
      | FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_15_sva_st_3) &
      (FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_5[49]))))))));
  assign mux_683_nl = MUX_s_1_2_2((nor_1374_nl), (mux_682_nl), or_cse_2);
  assign FpAdd_8U_23U_and_204_cse = core_wen & (~ and_dcpl_7) & (mux_683_nl);
  assign nor_1367_nl = ~(FpAdd_8U_23U_mux_226_tmp_49 | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1368_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | alu_loop_op_15_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm);
  assign mux_688_nl = MUX_s_1_2_2((nor_1368_nl), (nor_1367_nl), nor_333_cse);
  assign nor_1369_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205!=2'b10) | alu_loop_op_15_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2);
  assign mux_689_nl = MUX_s_1_2_2((nor_1369_nl), (mux_688_nl), or_cse_2);
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_29_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (mux_689_nl);
  assign nor_1365_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48) | (~ IsNaN_8U_23U_1_land_15_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_15_lpi_1_dfm_9 | IsNaN_8U_23U_3_land_15_lpi_1_dfm_7);
  assign nor_1366_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_15_lpi_1_dfm_10 | (cfg_alu_algo_1_sva_st_205!=2'b10)
      | (~ IsNaN_8U_23U_1_land_15_lpi_1_dfm_9) | IsNaN_8U_23U_land_15_lpi_1_dfm_st_5);
  assign mux_690_nl = MUX_s_1_2_2((nor_1366_nl), (nor_1365_nl), or_cse_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_94_ssc = core_wen & (~ and_dcpl_7)
      & (mux_690_nl);
  assign nor_1353_cse = ~((~ FpAlu_8U_23U_or_861_itm_3) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign and_3711_nl = nor_1743_cse & (~(alu_loop_op_16_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm
      & or_22_cse));
  assign and_3712_nl = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_st_2
      & (FpAdd_8U_23U_int_mant_p1_lpi_1_dfm[49]);
  assign mux_702_nl = MUX_s_1_2_2((and_3711_nl), nor_1743_cse, and_3712_nl);
  assign nor_1349_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & (~(alu_loop_op_16_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2
      & (~(((~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_2) |
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_st_3) & (FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49]))))))));
  assign mux_703_nl = MUX_s_1_2_2((nor_1349_nl), (mux_702_nl), or_cse_2);
  assign FpAdd_8U_23U_and_206_cse = core_wen & (~ and_dcpl_7) & (mux_703_nl);
  assign nor_1342_nl = ~(FpAdd_8U_23U_mux_242_tmp_49 | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1343_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | alu_loop_op_16_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm);
  assign mux_708_nl = MUX_s_1_2_2((nor_1343_nl), (nor_1342_nl), nor_333_cse);
  assign nor_1344_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205!=2'b10) | alu_loop_op_16_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2);
  assign mux_709_nl = MUX_s_1_2_2((nor_1344_nl), (mux_708_nl), or_cse_2);
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_30_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (mux_709_nl);
  assign nor_1340_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48) | (~ IsNaN_8U_23U_1_land_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_lpi_1_dfm_9 | IsNaN_8U_23U_3_land_lpi_1_dfm_7);
  assign nor_1341_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_lpi_1_dfm_10 | (cfg_alu_algo_1_sva_st_205!=2'b10)
      | (~ IsNaN_8U_23U_1_land_lpi_1_dfm_9) | IsNaN_8U_23U_land_lpi_1_dfm_st_5);
  assign mux_710_nl = MUX_s_1_2_2((nor_1341_nl), (nor_1340_nl), or_cse_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_95_ssc = core_wen & (~ and_dcpl_7)
      & (mux_710_nl);
  assign or_1811_nl = FpAlu_8U_23U_equal_tmp_237 | io_read_cfg_alu_bypass_rsc_svs_7
      | (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt | (~ main_stage_v_4);
  assign or_1812_nl = FpAlu_8U_23U_equal_tmp_237 | io_read_cfg_alu_bypass_rsc_svs_7;
  assign mux_718_nl = MUX_s_1_2_2(mux_tmp_339, or_tmp_670, or_1812_nl);
  assign mux_719_nl = MUX_s_1_2_2((mux_718_nl), (or_1811_nl), FpAlu_8U_23U_equal_tmp_146);
  assign FpAlu_8U_23U_and_849_cse = core_wen & (~ and_dcpl_7) & (~ (mux_719_nl));
  assign cfg_alu_algo_and_115_cse = core_wen & (~ and_dcpl_7) & (~ mux_tmp_339);
  assign or_1827_cse = io_read_cfg_alu_bypass_rsc_svs_7 | (~ reg_chn_alu_out_rsci_ld_core_psct_cse)
      | chn_alu_out_rsci_bawt | (~ main_stage_v_4);
  assign or_1825_nl = FpAlu_8U_23U_equal_tmp_146 | or_tmp_670;
  assign mux_347_nl = MUX_s_1_2_2(mux_tmp_339, or_tmp_670, io_read_cfg_alu_bypass_rsc_svs_7);
  assign mux_728_nl = MUX_s_1_2_2((mux_347_nl), or_1827_cse, FpAlu_8U_23U_equal_tmp_146);
  assign mux_729_nl = MUX_s_1_2_2((mux_728_nl), (or_1825_nl), FpAlu_8U_23U_equal_tmp_237);
  assign FpAlu_8U_23U_and_889_cse = core_wen & (~ and_dcpl_7) & (~ (mux_729_nl));
  assign AluIn_data_and_cse = core_wen & (~((~ and_91_tmp) | (fsm_output[0])));
  assign IsNaN_8U_23U_2_aelse_and_cse = core_wen & (~ (fsm_output[0]));
  assign and_3707_cse = (cfg_alu_algo_1_sva_st_15==2'b11);
  assign IsNaN_8U_23U_aelse_IsNaN_8U_23U_2_aelse_or_15_cse = and_dcpl_394 | and_dcpl_395;
  assign or_1861_nl = cfg_alu_bypass_rsci_d | ((cfg_alu_algo_rsci_d==2'b11) & (cfg_precision==2'b10));
  assign mux_750_nl = MUX_s_1_2_2((or_1861_nl), or_tmp_1848, and_3707_cse);
  assign mux_751_nl = MUX_s_1_2_2(or_tmp_20, (mux_750_nl), and_91_tmp);
  assign IsNaN_8U_23U_2_aelse_and_48_cse = IsNaN_8U_23U_2_aelse_and_cse & IsNaN_8U_23U_aelse_IsNaN_8U_23U_2_aelse_or_15_cse
      & (~ (mux_751_nl));
  assign cfg_alu_algo_and_132_cse = IsNaN_8U_23U_2_aelse_and_cse & IsNaN_8U_23U_aelse_IsNaN_8U_23U_2_aelse_or_15_cse
      & (~ mux_782_itm);
  assign cfg_alu_src_and_cse = IsNaN_8U_23U_2_aelse_and_cse & and_91_tmp & (~ mux_782_itm);
  assign FpAdd_8U_23U_and_208_cse = core_wen & (and_dcpl_402 | and_dcpl_407 | and_dcpl_408)
      & mux_tmp_156;
  assign FpNormalize_8U_49U_if_and_31_cse = IsNaN_8U_23U_2_aelse_and_cse & (~ or_dcpl_137)
      & (~ mux_tmp_778);
  assign FpAdd_8U_23U_int_mant_p1_and_cse = core_wen & (~(or_22_cse | io_read_cfg_alu_bypass_rsc_svs_st_6
      | and_dcpl_7 | (~ main_stage_v_3)));
  assign FpAdd_8U_23U_if_3_and_cse = core_wen & (~ or_dcpl_137);
  assign FpAdd_8U_23U_and_210_cse = core_wen & (and_dcpl_417 | and_dcpl_422 | and_dcpl_408)
      & mux_tmp_156;
  assign FpNormalize_8U_49U_if_and_32_cse = IsNaN_8U_23U_2_aelse_and_cse & (~ or_dcpl_137)
      & (~ mux_tmp_779);
  assign FpAdd_8U_23U_and_212_cse = core_wen & (and_dcpl_432 | and_dcpl_437 | and_dcpl_408)
      & mux_tmp_156;
  assign FpNormalize_8U_49U_if_and_33_cse = IsNaN_8U_23U_2_aelse_and_cse & (~ or_dcpl_137)
      & (~ mux_tmp_781);
  assign FpAdd_8U_23U_and_214_cse = core_wen & (and_dcpl_447 | and_dcpl_452 | and_dcpl_408)
      & mux_tmp_156;
  assign FpNormalize_8U_49U_if_and_34_cse = IsNaN_8U_23U_2_aelse_and_cse & (~ or_dcpl_137)
      & (~ mux_tmp_782);
  assign FpNormalize_8U_49U_if_and_35_cse = IsNaN_8U_23U_2_aelse_and_cse & (~ or_dcpl_137)
      & (~ mux_tmp_783);
  assign FpNormalize_8U_49U_if_and_36_cse = IsNaN_8U_23U_2_aelse_and_cse & (~ or_dcpl_137)
      & (~ mux_tmp_785);
  assign FpNormalize_8U_49U_if_and_37_cse = IsNaN_8U_23U_2_aelse_and_cse & (~ or_dcpl_137)
      & (~ mux_tmp_786);
  assign FpAdd_8U_23U_and_216_cse = core_wen & (and_dcpl_474 | and_dcpl_479 | and_dcpl_408)
      & mux_tmp_156;
  assign FpNormalize_8U_49U_if_and_38_cse = IsNaN_8U_23U_2_aelse_and_cse & (~ or_dcpl_137)
      & (~ mux_tmp_787);
  assign FpNormalize_8U_49U_if_and_39_cse = IsNaN_8U_23U_2_aelse_and_cse & (~ or_dcpl_137)
      & (~ mux_tmp_788);
  assign FpNormalize_8U_49U_if_and_40_cse = IsNaN_8U_23U_2_aelse_and_cse & (~ or_dcpl_137)
      & (~ mux_tmp_789);
  assign FpNormalize_8U_49U_if_and_41_cse = IsNaN_8U_23U_2_aelse_and_cse & (~ or_dcpl_137)
      & (~ mux_tmp_790);
  assign FpNormalize_8U_49U_if_and_42_cse = IsNaN_8U_23U_2_aelse_and_cse & (~ or_dcpl_137)
      & (~ mux_tmp_791);
  assign FpAdd_8U_23U_and_218_cse = core_wen & (and_dcpl_505 | and_dcpl_510 | and_dcpl_408)
      & mux_tmp_156;
  assign FpNormalize_8U_49U_if_and_43_cse = IsNaN_8U_23U_2_aelse_and_cse & (~ or_dcpl_137)
      & (~ mux_tmp_792);
  assign FpAdd_8U_23U_and_220_cse = core_wen & (and_dcpl_520 | and_dcpl_525 | and_dcpl_408)
      & mux_tmp_156;
  assign FpNormalize_8U_49U_if_and_44_cse = IsNaN_8U_23U_2_aelse_and_cse & (~ or_dcpl_137)
      & (~ mux_tmp_793);
  assign FpAdd_8U_23U_and_222_cse = core_wen & (and_dcpl_535 | and_dcpl_540 | and_dcpl_408)
      & mux_tmp_156;
  assign FpNormalize_8U_49U_if_and_45_cse = IsNaN_8U_23U_2_aelse_and_cse & (~ or_dcpl_137)
      & (~ mux_tmp_795);
  assign FpAdd_8U_23U_and_224_cse = core_wen & (and_dcpl_550 | and_dcpl_555 | and_dcpl_408)
      & mux_tmp_156;
  assign FpNormalize_8U_49U_if_and_46_cse = IsNaN_8U_23U_2_aelse_and_cse & (~ or_dcpl_137)
      & (~ mux_tmp_796);
  assign alu_loop_op_else_if_and_cse = core_wen & (~(or_dcpl_219 | and_dcpl_7 | or_dcpl_116));
  assign alu_loop_op_else_else_if_and_cse = core_wen & (~(or_dcpl_219 | and_dcpl_7
      | or_dcpl_113));
  assign FpAdd_8U_23U_and_226_cse = core_wen & (and_dcpl_565 | and_dcpl_570 | and_dcpl_408)
      & mux_tmp_156;
  assign FpAdd_8U_23U_and_228_cse = core_wen & (and_dcpl_576 | and_dcpl_581 | and_dcpl_408)
      & mux_tmp_156;
  assign FpAdd_8U_23U_and_230_cse = core_wen & (and_dcpl_587 | and_dcpl_592 | and_dcpl_408)
      & mux_tmp_156;
  assign FpAdd_8U_23U_and_232_cse = core_wen & (and_dcpl_598 | and_dcpl_603 | and_dcpl_408)
      & mux_tmp_156;
  assign FpAdd_8U_23U_and_234_cse = core_wen & (and_dcpl_609 | and_dcpl_614 | and_dcpl_408)
      & mux_tmp_156;
  assign FpAdd_8U_23U_and_236_cse = core_wen & (and_dcpl_620 | and_dcpl_625 | and_dcpl_408)
      & mux_tmp_156;
  assign FpAdd_8U_23U_and_238_cse = core_wen & (and_dcpl_631 | and_dcpl_636 | and_dcpl_408)
      & mux_tmp_156;
  assign FpAdd_8U_23U_b_left_shift_and_cse = core_wen & (~(or_22_cse | (~ main_stage_v_2)
      | io_read_cfg_alu_bypass_rsc_svs_st_5 | and_dcpl_7 | or_350_cse));
  assign and_1106_rgt = (or_dcpl_14 | (cfg_alu_algo_1_sva_st_92!=2'b10)) & and_89_tmp;
  assign and_1105_cse = and_dcpl_638 & and_543_rgt;
  assign IsZero_8U_23U_1_and_24_cse = core_wen & (and_1105_cse | and_1106_rgt);
  assign and_1108_rgt = (or_dcpl_14 | or_dcpl_295) & and_89_tmp;
  assign IsZero_8U_23U_1_and_25_cse = core_wen & (and_1105_cse | and_1108_rgt);
  assign or_1935_cse = io_read_cfg_alu_bypass_rsc_svs_st_6 | (~ main_stage_v_3);
  assign or_1923_cse = (~ (cfg_alu_algo_1_sva_5[0])) | (reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign and_1135_rgt = or_cse_2 & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b01);
  assign nor_577_cse = ~(FpAlu_8U_23U_equal_tmp_2 | (~ (reg_cfg_alu_algo_1_sva_st_93_cse[0])));
  assign or_1938_cse = (~ FpAlu_8U_23U_equal_tmp_144) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign IsNaN_8U_23U_1_aelse_or_5_cse = and_1318_cse | and_1135_rgt;
  assign IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_1_aelse_or_5_cse = and_1141_cse | and_1318_cse
      | and_1135_rgt;
  assign or_1922_nl = (cfg_alu_algo_1_sva_5[0]) | (reg_cfg_alu_algo_1_sva_st_93_cse!=2'b10)
      | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign or_1927_nl = (~ (reg_cfg_alu_algo_1_sva_st_93_cse[0])) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign mux_804_nl = MUX_s_1_2_2((or_1927_nl), or_tmp_1915, or_1923_cse);
  assign mux_805_cse = MUX_s_1_2_2((mux_804_nl), (or_1922_nl), cfg_alu_algo_1_sva_5[1]);
  assign or_1931_nl = nor_577_cse | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign nand_448_nl = ~(FpAlu_8U_23U_equal_tmp_2 & (reg_cfg_alu_algo_1_sva_st_93_cse[0])
      & (~ io_read_cfg_alu_bypass_rsc_svs_st_5) & main_stage_v_2);
  assign mux_807_cse = MUX_s_1_2_2((nand_448_nl), (or_1931_nl), FpAlu_8U_23U_equal_tmp);
  assign or_1937_nl = (~ FpAlu_8U_23U_equal_tmp_148) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_811_cse = MUX_s_1_2_2(or_1938_cse, (or_1937_nl), cfg_alu_algo_1_sva_st_204[0]);
  assign and_3689_cse = (cfg_alu_algo_1_sva_5==2'b11);
  assign nor_1317_cse = ~(io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign nor_1315_nl = ~(and_3689_cse | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~
      main_stage_v_2));
  assign nor_1316_nl = ~((reg_cfg_alu_algo_1_sva_st_93_cse!=2'b10) | (~ FpAlu_8U_23U_nor_dfs)
      | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_814_nl = MUX_s_1_2_2(nor_1317_cse, (nor_1316_nl), FpAlu_8U_23U_equal_tmp_1);
  assign mux_815_nl = MUX_s_1_2_2((mux_814_nl), (nor_1315_nl), nor_333_cse);
  assign nor_1318_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (FpAlu_8U_23U_equal_tmp_146 & ((cfg_alu_algo_1_sva_st_204[0]) | (~((cfg_alu_algo_1_sva_st_204[1])
      & FpAlu_8U_23U_nor_dfs_48)))));
  assign mux_816_nl = MUX_s_1_2_2((nor_1318_nl), (mux_815_nl), or_cse_2);
  assign IsNaN_8U_23U_aelse_and_47_cse = core_wen & (~ and_dcpl_7) & (mux_816_nl);
  assign nor_1305_nl = ~((cfg_alu_algo_1_sva_5[1]) | (reg_cfg_alu_algo_1_sva_st_93_cse[0])
      | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign nor_1306_nl = ~((cfg_alu_algo_1_sva_5[1]) | (~ (reg_cfg_alu_algo_1_sva_st_93_cse[0]))
      | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_817_nl = MUX_s_1_2_2((nor_1306_nl), (nor_1305_nl), reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign nor_1307_nl = ~((~((reg_cfg_alu_algo_1_sva_st_93_cse[1]) | (~ (cfg_alu_algo_1_sva_5[1]))))
      | (reg_cfg_alu_algo_1_sva_st_93_cse[0]) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (~ main_stage_v_2));
  assign mux_818_cse = MUX_s_1_2_2((nor_1307_nl), (mux_817_nl), cfg_alu_algo_1_sva_5[0]);
  assign nor_1309_nl = ~(nor_577_cse | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign and_4250_nl = FpAlu_8U_23U_equal_tmp_2 & (reg_cfg_alu_algo_1_sva_st_93_cse[0])
      & (~ io_read_cfg_alu_bypass_rsc_svs_st_5) & main_stage_v_2;
  assign mux_819_cse = MUX_s_1_2_2((and_4250_nl), (nor_1309_nl), FpAlu_8U_23U_equal_tmp);
  assign mux_823_cse = MUX_s_1_2_2(nor_1930_cse, nor_1928_cse, cfg_alu_algo_1_sva_st_204[0]);
  assign nor_1312_cse = ~((cfg_alu_algo_1_sva_st_204[0]) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign IsNaN_8U_23U_1_aelse_and_34_cse = core_wen & (~ and_dcpl_7) & (~ mux_tmp_823);
  assign and_1141_cse = or_cse_2 & (reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign IsNaN_8U_23U_1_aelse_or_3_cse = and_1421_cse | and_1135_rgt;
  assign IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_1_aelse_or_3_cse = and_1141_cse | and_1421_cse
      | and_1135_rgt;
  assign nor_1222_nl = ~((~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (~ alu_loop_op_else_nor_tmp_80));
  assign mux_912_nl = MUX_s_1_2_2(nor_1815_cse, (nor_1222_nl), or_cse_2);
  assign AluOut_data_and_16_cse = core_wen & (~ and_dcpl_7) & (mux_912_nl);
  assign mux_1631_cse = MUX_s_1_2_2(FpAlu_8U_23U_equal_tmp_1, and_3689_cse, nor_333_cse);
  assign and_3670_nl = main_stage_v_2 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5) &
      mux_1631_cse;
  assign mux_930_nl = MUX_s_1_2_2(nor_1813_cse, (and_3670_nl), or_cse_2);
  assign FpAlu_8U_23U_o_and_16_cse = core_wen & (~ and_dcpl_7) & (mux_930_nl);
  assign nor_1173_nl = ~((cfg_alu_algo_1_sva_5[0]) | (~ alu_loop_op_else_nor_tmp_80));
  assign mux_976_nl = MUX_s_1_2_2((nor_1173_nl), alu_loop_op_else_nor_tmp_80, cfg_alu_algo_1_sva_5[1]);
  assign nor_1172_nl = ~((~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (mux_976_nl));
  assign mux_980_cse = MUX_s_1_2_2(nor_1862_cse, (nor_1172_nl), or_cse_2);
  assign alu_loop_op_else_else_if_and_105_cse = core_wen & (and_dcpl_698 | and_dcpl_701
      | and_dcpl_704 | and_dcpl_707) & mux_980_cse;
  assign alu_loop_op_else_else_if_and_108_cse = core_wen & (and_dcpl_711 | and_dcpl_714
      | and_dcpl_704 | and_dcpl_707) & mux_980_cse;
  assign alu_loop_op_else_else_if_and_111_cse = core_wen & (and_dcpl_722 | and_dcpl_725
      | and_dcpl_704 | and_dcpl_707) & mux_980_cse;
  assign alu_loop_op_else_else_if_and_114_cse = core_wen & (and_dcpl_733 | and_dcpl_736
      | and_dcpl_704 | and_dcpl_707) & mux_980_cse;
  assign alu_loop_op_else_else_if_and_117_cse = core_wen & (and_dcpl_744 | and_dcpl_747
      | and_dcpl_704 | and_dcpl_707) & mux_980_cse;
  assign alu_loop_op_else_else_if_and_120_cse = core_wen & (and_dcpl_755 | and_dcpl_758
      | and_dcpl_704 | and_dcpl_707) & mux_980_cse;
  assign alu_loop_op_else_else_if_and_123_cse = core_wen & (and_dcpl_766 | and_dcpl_769
      | and_dcpl_704 | and_dcpl_707) & mux_980_cse;
  assign alu_loop_op_else_else_if_and_126_cse = core_wen & (and_dcpl_777 | and_dcpl_780
      | and_dcpl_704 | and_dcpl_707) & mux_980_cse;
  assign alu_loop_op_else_else_if_and_129_cse = core_wen & (and_dcpl_788 | and_dcpl_791
      | and_dcpl_704 | and_dcpl_707) & mux_980_cse;
  assign alu_loop_op_else_else_if_and_132_cse = core_wen & (and_dcpl_799 | and_dcpl_802
      | and_dcpl_704 | and_dcpl_707) & mux_980_cse;
  assign alu_loop_op_else_else_if_and_135_cse = core_wen & (and_dcpl_810 | and_dcpl_813
      | and_dcpl_704 | and_dcpl_707) & mux_980_cse;
  assign alu_loop_op_else_else_if_and_138_cse = core_wen & (and_dcpl_821 | and_dcpl_824
      | and_dcpl_704 | and_dcpl_707) & mux_980_cse;
  assign alu_loop_op_else_else_if_and_141_cse = core_wen & (and_dcpl_832 | and_dcpl_834
      | and_dcpl_704 | and_dcpl_707) & mux_980_cse;
  assign nor_1122_nl = ~(io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2)
      | mux_1631_cse);
  assign nor_1123_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign mux_1042_nl = MUX_s_1_2_2((nor_1123_nl), (nor_1122_nl), or_cse_2);
  assign FpAlu_8U_23U_and_976_cse = core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
      & (mux_1042_nl);
  assign FpAlu_8U_23U_FpAlu_8U_23U_or_79_cse = (and_dcpl_398 & or_cse_2) | and_dcpl_840;
  assign FpAlu_8U_23U_and_1040_cse = core_wen & FpAlu_8U_23U_FpAlu_8U_23U_or_79_cse
      & (~ mux_tmp_823);
  assign FpAlu_8U_23U_and_1056_cse = core_wen & FpAlu_8U_23U_FpAlu_8U_23U_or_79_cse
      & mux_tmp_156;
  assign and_1308_rgt = or_cse_2 & and_dcpl_397;
  assign and_1307_cse = or_cse_2 & (reg_cfg_alu_algo_1_sva_st_93_cse[0]);
  assign mux_1076_nl = MUX_s_1_2_2((~ or_1923_cse), or_1923_cse, reg_cfg_alu_algo_1_sva_st_93_cse[0]);
  assign mux_1077_nl = MUX_s_1_2_2((mux_1076_nl), or_350_cse, cfg_alu_algo_1_sva_5[1]);
  assign or_2484_nl = (~ FpAlu_8U_23U_equal_tmp_2) | (reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign nor_1088_nl = ~(FpAlu_8U_23U_equal_tmp | (reg_cfg_alu_algo_1_sva_st_93_cse[1]));
  assign mux_1078_nl = MUX_s_1_2_2((nor_1088_nl), (or_2484_nl), reg_cfg_alu_algo_1_sva_st_93_cse[0]);
  assign mux_1079_nl = MUX_s_1_2_2((mux_1078_nl), (mux_1077_nl), nor_333_cse);
  assign nor_1087_nl = ~(io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2)
      | (mux_1079_nl));
  assign or_2487_nl = (~ FpAlu_8U_23U_equal_tmp_148) | (cfg_alu_algo_1_sva_st_204[1]);
  assign nor_1090_nl = ~(FpAlu_8U_23U_equal_tmp_144 | (cfg_alu_algo_1_sva_st_204[1]));
  assign mux_1081_nl = MUX_s_1_2_2((nor_1090_nl), (or_2487_nl), cfg_alu_algo_1_sva_st_204[0]);
  assign nor_1089_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (mux_1081_nl));
  assign mux_1082_cse = MUX_s_1_2_2((nor_1089_nl), (nor_1087_nl), or_cse_2);
  assign IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_15_cse = and_1318_cse | and_1307_cse
      | and_1308_rgt;
  assign IsNaN_8U_23U_3_aelse_and_cse = core_wen & IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_15_cse
      & mux_1082_cse;
  assign and_1311_rgt = and_dcpl_844 & and_dcpl_843;
  assign and_1313_rgt = and_dcpl_846 & and_dcpl_843;
  assign and_1315_rgt = and_dcpl_844 & and_dcpl_848;
  assign and_1316_rgt = and_dcpl_846 & and_dcpl_848;
  assign mux_1085_nl = MUX_s_1_2_2((reg_cfg_alu_algo_1_sva_st_93_cse[0]), (~ (reg_cfg_alu_algo_1_sva_st_93_cse[0])),
      cfg_alu_algo_1_sva_5[0]);
  assign nor_1085_nl = ~((cfg_alu_algo_1_sva_5[1]) | (mux_1085_nl));
  assign mux_1086_nl = MUX_s_1_2_2(mux_tmp_1077, (nor_1085_nl), cfg_precision[1]);
  assign mux_1087_nl = MUX_s_1_2_2((mux_1086_nl), mux_tmp_1077, cfg_precision[0]);
  assign nor_1084_nl = ~(io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ (mux_1087_nl)));
  assign mux_1088_nl = MUX_s_1_2_2((nor_1084_nl), (~ (reg_cfg_alu_algo_1_sva_st_93_cse[0])),
      reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign and_3622_nl = nor_1317_cse & (mux_1088_nl);
  assign mux_1090_nl = MUX_s_1_2_2(FpAlu_8U_23U_equal_tmp_144, FpAlu_8U_23U_equal_tmp_148,
      cfg_alu_algo_1_sva_st_204[0]);
  assign mux_1091_nl = MUX_s_1_2_2((mux_1090_nl), (~ (cfg_alu_algo_1_sva_st_204[0])),
      cfg_alu_algo_1_sva_st_204[1]);
  assign and_4266_nl = main_stage_v_3 & (~ io_read_cfg_alu_bypass_rsc_svs_st_6) &
      (mux_1091_nl);
  assign mux_1092_cse = MUX_s_1_2_2((and_4266_nl), (and_3622_nl), or_cse_2);
  assign and_1318_cse = or_cse_2 & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b00);
  assign IsNaN_8U_23U_3_aelse_and_1_cse = core_wen & IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_15_cse
      & mux_1092_cse;
  assign and_1323_rgt = and_dcpl_856 & and_dcpl_843;
  assign and_1325_rgt = and_dcpl_858 & and_dcpl_843;
  assign and_1327_rgt = and_dcpl_856 & and_dcpl_848;
  assign and_1328_rgt = and_dcpl_858 & and_dcpl_848;
  assign IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_13_cse = and_1421_cse | and_1307_cse
      | and_1308_rgt;
  assign IsNaN_8U_23U_3_aelse_and_2_cse = core_wen & IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_13_cse
      & mux_1082_cse;
  assign and_1333_rgt = or_cse_2 & (AluIn_data_sva_501[95]) & (reg_cfg_alu_algo_1_sva_st_93_cse[0]);
  assign and_1335_rgt = or_cse_2 & (~ (AluIn_data_sva_501[95])) & (reg_cfg_alu_algo_1_sva_st_93_cse[0]);
  assign and_1337_rgt = or_cse_2 & (AluIn_data_sva_501[95]) & and_dcpl_676;
  assign and_1339_rgt = or_cse_2 & (~ (AluIn_data_sva_501[95])) & and_dcpl_676;
  assign and_1346_rgt = and_dcpl_879 & (~ (cfg_precision[0])) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10);
  assign and_1347_rgt = and_dcpl_241 & and_dcpl_397;
  assign and_1351_rgt = and_dcpl_884 & and_dcpl_843;
  assign and_1353_rgt = and_dcpl_886 & and_dcpl_843;
  assign and_1355_rgt = and_dcpl_884 & and_dcpl_848;
  assign and_1356_rgt = and_dcpl_886 & and_dcpl_848;
  assign and_1364_rgt = and_dcpl_897 & and_dcpl_843;
  assign and_1366_rgt = and_dcpl_899 & and_dcpl_843;
  assign and_1368_rgt = and_dcpl_897 & and_dcpl_848;
  assign and_1369_rgt = and_dcpl_899 & and_dcpl_848;
  assign IsNaN_8U_23U_3_aelse_or_1_cse = and_1421_cse | and_1307_cse;
  assign IsNaN_8U_23U_3_aelse_and_5_cse = core_wen & (and_1421_cse | and_1307_cse
      | and_1346_rgt | and_1347_rgt) & mux_1092_cse;
  assign and_1380_rgt = or_cse_2 & (AluIn_data_sva_501[191]) & (reg_cfg_alu_algo_1_sva_st_93_cse[0]);
  assign and_1382_rgt = or_cse_2 & (~ (AluIn_data_sva_501[191])) & (reg_cfg_alu_algo_1_sva_st_93_cse[0]);
  assign and_1384_rgt = or_cse_2 & (AluIn_data_sva_501[191]) & and_dcpl_676;
  assign and_1386_rgt = or_cse_2 & (~ (AluIn_data_sva_501[191])) & and_dcpl_676;
  assign and_1391_rgt = and_dcpl_924 & and_dcpl_843;
  assign and_1393_rgt = and_dcpl_926 & and_dcpl_843;
  assign and_1395_rgt = and_dcpl_924 & and_dcpl_848;
  assign and_1396_rgt = and_dcpl_926 & and_dcpl_848;
  assign and_1400_rgt = or_cse_2 & (AluIn_data_sva_501[255]) & (reg_cfg_alu_algo_1_sva_st_93_cse[0]);
  assign and_1402_rgt = or_cse_2 & (~ (AluIn_data_sva_501[255])) & (reg_cfg_alu_algo_1_sva_st_93_cse[0]);
  assign and_1404_rgt = or_cse_2 & (AluIn_data_sva_501[255]) & and_dcpl_676;
  assign and_1406_rgt = or_cse_2 & (~ (AluIn_data_sva_501[255])) & and_dcpl_676;
  assign and_1413_rgt = and_dcpl_946 & and_dcpl_843;
  assign and_1415_rgt = and_dcpl_948 & and_dcpl_843;
  assign and_1417_rgt = and_dcpl_946 & and_dcpl_848;
  assign and_1418_rgt = and_dcpl_948 & and_dcpl_848;
  assign and_1421_cse = or_cse_2 & and_dcpl_676;
  assign IsNaN_8U_23U_3_aelse_and_9_cse = core_wen & IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_13_cse
      & mux_1092_cse;
  assign and_1425_rgt = or_cse_2 & (AluIn_data_sva_501[319]) & (reg_cfg_alu_algo_1_sva_st_93_cse[0]);
  assign and_1427_rgt = or_cse_2 & (~ (AluIn_data_sva_501[319])) & (reg_cfg_alu_algo_1_sva_st_93_cse[0]);
  assign and_1429_rgt = or_cse_2 & (AluIn_data_sva_501[319]) & and_dcpl_676;
  assign and_1431_rgt = or_cse_2 & (~ (AluIn_data_sva_501[319])) & and_dcpl_676;
  assign and_1438_rgt = and_dcpl_971 & (AluIn_data_sva_501[351]) & (cfg_alu_algo_1_sva_5[0]);
  assign and_1440_rgt = and_dcpl_971 & (~ (AluIn_data_sva_501[351])) & (cfg_alu_algo_1_sva_5[0]);
  assign and_1442_rgt = and_dcpl_971 & (AluIn_data_sva_501[351]) & (~ (cfg_alu_algo_1_sva_5[0]));
  assign and_1444_rgt = and_dcpl_971 & (~ (AluIn_data_sva_501[351])) & (~ (cfg_alu_algo_1_sva_5[0]));
  assign and_1452_rgt = and_dcpl_971 & (AluIn_data_sva_501[383]) & (cfg_alu_algo_1_sva_5[0]);
  assign and_1454_rgt = and_dcpl_971 & (~ (AluIn_data_sva_501[383])) & (cfg_alu_algo_1_sva_5[0]);
  assign and_1456_rgt = and_dcpl_971 & (AluIn_data_sva_501[383]) & (~ (cfg_alu_algo_1_sva_5[0]));
  assign and_1458_rgt = and_dcpl_971 & (~ (AluIn_data_sva_501[383])) & (~ (cfg_alu_algo_1_sva_5[0]));
  assign and_1469_rgt = or_cse_2 & (AluIn_data_sva_501[415]) & (reg_cfg_alu_algo_1_sva_st_93_cse[0]);
  assign and_1471_rgt = or_cse_2 & (~ (AluIn_data_sva_501[415])) & (reg_cfg_alu_algo_1_sva_st_93_cse[0]);
  assign and_1473_rgt = or_cse_2 & (AluIn_data_sva_501[415]) & and_dcpl_676;
  assign and_1475_rgt = or_cse_2 & (~ (AluIn_data_sva_501[415])) & and_dcpl_676;
  assign and_1481_rgt = or_cse_2 & (AluIn_data_sva_501[447]) & (reg_cfg_alu_algo_1_sva_st_93_cse[0]);
  assign and_1483_rgt = or_cse_2 & (~ (AluIn_data_sva_501[447])) & (reg_cfg_alu_algo_1_sva_st_93_cse[0]);
  assign and_1485_rgt = or_cse_2 & (AluIn_data_sva_501[447]) & and_dcpl_676;
  assign and_1487_rgt = or_cse_2 & (~ (AluIn_data_sva_501[447])) & and_dcpl_676;
  assign and_1492_rgt = and_dcpl_971 & (AluIn_data_sva_501[479]) & (cfg_alu_algo_1_sva_5[0]);
  assign and_1494_rgt = and_dcpl_971 & (~ (AluIn_data_sva_501[479])) & (cfg_alu_algo_1_sva_5[0]);
  assign and_1496_rgt = and_dcpl_971 & (AluIn_data_sva_501[479]) & (~ (cfg_alu_algo_1_sva_5[0]));
  assign and_1498_rgt = and_dcpl_971 & (~ (AluIn_data_sva_501[479])) & (~ (cfg_alu_algo_1_sva_5[0]));
  assign and_1503_rgt = and_dcpl_1036 & and_dcpl_843;
  assign and_1505_rgt = and_dcpl_1038 & and_dcpl_843;
  assign and_1507_rgt = and_dcpl_1036 & and_dcpl_848;
  assign and_1508_rgt = and_dcpl_1038 & and_dcpl_848;
  assign or_2817_nl = (reg_cfg_alu_algo_1_sva_st_110_cse[1]) | (~ reg_chn_alu_out_rsci_ld_core_psct_cse)
      | chn_alu_out_rsci_bawt | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign mux_1348_nl = MUX_s_1_2_2(mux_tmp_149, or_tmp_327, reg_cfg_alu_algo_1_sva_st_110_cse[1]);
  assign mux_1349_cse = MUX_s_1_2_2((mux_1348_nl), (or_2817_nl), reg_cfg_alu_algo_1_sva_st_157_cse[1]);
  assign alu_loop_op_else_else_if_and_144_cse = core_wen & (and_dcpl_1044 | and_dcpl_1046
      | and_dcpl_1048 | and_dcpl_1050) & (~ mux_1349_cse);
  assign alu_loop_op_else_else_if_and_147_cse = core_wen & (and_dcpl_1052 | and_dcpl_1054
      | and_dcpl_1048 | and_dcpl_1050) & (~ mux_1349_cse);
  assign or_2819_nl = (reg_cfg_alu_algo_1_sva_st_157_cse[1]) | or_tmp_327;
  assign mux_1352_nl = MUX_s_1_2_2(mux_tmp_149, or_tmp_329, reg_cfg_alu_algo_1_sva_st_157_cse[1]);
  assign mux_1353_nl = MUX_s_1_2_2((mux_1352_nl), (or_2819_nl), reg_cfg_alu_algo_1_sva_st_110_cse[1]);
  assign alu_loop_op_else_else_if_and_150_cse = core_wen & (and_dcpl_1060 | and_dcpl_1062
      | and_dcpl_1048 | and_dcpl_1050) & (~ (mux_1353_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_14_cse = core_wen & ((and_dcpl_1073
      & and_dcpl_1070 & (else_mux_2_tmp[1]) & and_89_tmp & (~ IsNaN_5U_23U_nor_tmp)
      & (fsm_output[1])) | or_tmp_3190);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_15_cse = core_wen & (~(or_dcpl_393
      | (fsm_output[0])));
  assign FpAdd_8U_23U_is_a_greater_and_cse = core_wen & (~(or_dcpl_14 | or_dcpl_394
      | (~ (cfg_alu_algo_1_sva_st_92[1]))));
  assign FpCmp_8U_23U_true_if_and_cse = core_wen & (~(or_dcpl_14 | or_dcpl_394 |
      (cfg_alu_algo_1_sva_st_92[1]) | (fsm_output[0])));
  assign FpCmp_8U_23U_false_if_and_cse = core_wen & (~(or_dcpl_14 | (~ and_89_tmp)
      | (cfg_alu_algo_1_sva_st_92!=2'b01)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_17_cse = core_wen & ((and_dcpl_1087
      & and_dcpl_1084 & (else_mux_5_tmp[0]) & and_89_tmp & (~ IsNaN_5U_23U_nor_1_tmp)
      & (fsm_output[1])) | or_tmp_3201);
  assign FpAdd_8U_23U_is_a_greater_and_1_cse = core_wen & (~ or_dcpl_414);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_20_cse = core_wen & ((and_dcpl_1101
      & and_dcpl_1098 & (else_mux_8_tmp[0]) & and_89_tmp & (~ IsNaN_5U_23U_nor_2_tmp)
      & (fsm_output[1])) | or_tmp_3212);
  assign FpAdd_8U_23U_is_a_greater_and_3_cse = core_wen & (~(or_dcpl_14 | or_dcpl_413));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_23_cse = core_wen & ((and_dcpl_1115
      & and_dcpl_1112 & (else_mux_11_tmp[0]) & and_89_tmp & (~ IsNaN_5U_23U_nor_3_tmp)
      & (fsm_output[1])) | or_tmp_3223);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_26_cse = core_wen & ((and_dcpl_1129
      & and_dcpl_1126 & and_dcpl_1123 & and_89_tmp & (fsm_output[1])) | or_tmp_3234);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_29_cse = core_wen & ((and_dcpl_638
      & or_dcpl_477 & (else_mux_17_tmp==5'b11111) & (~ IsNaN_5U_23U_nor_5_tmp) &
      and_89_tmp & (fsm_output[1])) | or_tmp_3245);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_32_cse = core_wen & ((and_dcpl_638
      & or_dcpl_495 & (else_mux_20_tmp==5'b11111) & (~ IsNaN_5U_23U_nor_6_tmp) &
      and_89_tmp & (fsm_output[1])) | or_tmp_3256);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_35_cse = core_wen & ((and_dcpl_638
      & or_dcpl_513 & (else_mux_23_tmp==5'b11111) & (~ IsNaN_5U_23U_nor_7_tmp) &
      and_89_tmp & (fsm_output[1])) | or_tmp_3267);
  assign FpAdd_8U_23U_is_a_greater_and_8_cse = core_wen & (~(or_dcpl_14 | or_dcpl_520));
  assign FpCmp_8U_23U_true_if_and_7_cse = core_wen & (~(or_dcpl_14 | (cfg_alu_algo_1_sva_st_92!=2'b00)
      | (~ and_89_tmp) | (fsm_output[0])));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_38_cse = core_wen & ((and_dcpl_638
      & or_dcpl_531 & (else_mux_26_tmp==5'b11111) & (~ IsNaN_5U_23U_nor_8_tmp) &
      and_89_tmp & (fsm_output[1])) | or_tmp_3278);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_41_cse = core_wen & ((and_dcpl_1214
      & and_dcpl_1211 & (else_mux_29_tmp[4]) & and_89_tmp & (~ IsNaN_5U_23U_nor_9_tmp)
      & (fsm_output[1])) | or_tmp_3289);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_44_cse = core_wen & ((and_dcpl_638
      & or_dcpl_567 & (else_mux_32_tmp==5'b11111) & (~ IsNaN_5U_23U_nor_10_tmp) &
      and_89_tmp & (fsm_output[1])) | or_tmp_3300);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_47_cse = core_wen & ((and_dcpl_638
      & or_dcpl_585 & (else_mux_35_tmp==5'b11111) & (~ IsNaN_5U_23U_nor_11_tmp) &
      and_89_tmp & (fsm_output[1])) | or_tmp_3311);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_50_cse = core_wen & ((and_dcpl_638
      & or_dcpl_603 & (else_mux_38_tmp==5'b11111) & (~ IsNaN_5U_23U_nor_12_tmp) &
      and_89_tmp & (fsm_output[1])) | or_tmp_3322);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_53_cse = core_wen & ((and_dcpl_1283
      & and_dcpl_1279 & (else_mux_41_tmp[0]) & and_89_tmp & (~ IsNaN_5U_23U_nor_13_tmp)
      & (fsm_output[1])) | or_tmp_3333);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_56_cse = core_wen & ((and_dcpl_638
      & or_dcpl_639 & (else_mux_44_tmp==5'b11111) & (~ IsNaN_5U_23U_nor_14_tmp) &
      and_89_tmp & (fsm_output[1])) | or_tmp_3344);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_59_cse = core_wen & ((and_dcpl_638
      & or_dcpl_657 & (else_mux_47_tmp==5'b11111) & (~ IsNaN_5U_23U_nor_15_tmp) &
      and_89_tmp & (fsm_output[1])) | or_tmp_3355);
  assign nor_920_nl = ~(cfg_alu_bypass_rsci_d | (cfg_alu_algo_rsci_d!=2'b11) | (cfg_precision!=2'b10));
  assign mux_1390_nl = MUX_s_1_2_2((nor_920_nl), or_tmp_1848, and_3707_cse);
  assign mux_1391_nl = MUX_s_1_2_2(and_3707_cse, (mux_1390_nl), and_91_tmp);
  assign IsNaN_8U_23U_2_aelse_and_74_cse = IsNaN_8U_23U_2_aelse_and_cse & (~ or_dcpl_675)
      & (~ (mux_1391_nl));
  assign FpAdd_8U_23U_and_144_cse = core_wen & ((and_dcpl_401 & and_dcpl_1329 & (~
      io_read_cfg_alu_bypass_rsc_svs_st_5) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10))
      | and_dcpl_1335);
  assign FpAdd_8U_23U_and_146_cse = core_wen & ((and_dcpl_416 & and_dcpl_1329 & (~
      io_read_cfg_alu_bypass_rsc_svs_st_5) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10))
      | and_dcpl_1341);
  assign FpAdd_8U_23U_and_148_cse = core_wen & ((and_dcpl_431 & and_dcpl_1329 & (~
      io_read_cfg_alu_bypass_rsc_svs_st_5) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10))
      | and_dcpl_1347);
  assign FpAdd_8U_23U_and_150_cse = core_wen & ((and_dcpl_446 & and_dcpl_1329 & (~
      io_read_cfg_alu_bypass_rsc_svs_st_5) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10))
      | and_dcpl_1353);
  assign FpAdd_8U_23U_and_152_cse = core_wen & ((and_dcpl_564 & and_dcpl_1329 & (~
      io_read_cfg_alu_bypass_rsc_svs_st_5) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10))
      | and_dcpl_1359);
  assign FpAdd_8U_23U_and_154_cse = core_wen & ((and_dcpl_575 & and_dcpl_1329 & (~
      io_read_cfg_alu_bypass_rsc_svs_st_5) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10))
      | and_dcpl_1365);
  assign FpAdd_8U_23U_and_156_cse = core_wen & ((and_dcpl_586 & and_dcpl_1329 & (~
      io_read_cfg_alu_bypass_rsc_svs_st_5) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10))
      | and_dcpl_1371);
  assign FpAdd_8U_23U_and_158_cse = core_wen & ((and_dcpl_473 & and_dcpl_1329 & (~
      io_read_cfg_alu_bypass_rsc_svs_st_5) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10))
      | and_dcpl_1377);
  assign FpAdd_8U_23U_and_160_cse = core_wen & ((and_dcpl_597 & and_dcpl_1329 & (~
      io_read_cfg_alu_bypass_rsc_svs_st_5) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10))
      | and_dcpl_1383);
  assign FpAdd_8U_23U_and_162_cse = core_wen & ((and_dcpl_608 & and_dcpl_1329 & (~
      io_read_cfg_alu_bypass_rsc_svs_st_5) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10))
      | and_dcpl_1389);
  assign FpAdd_8U_23U_and_164_cse = core_wen & ((and_dcpl_619 & and_dcpl_1329 & (~
      io_read_cfg_alu_bypass_rsc_svs_st_5) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10))
      | and_dcpl_1395);
  assign FpAdd_8U_23U_and_166_cse = core_wen & ((and_dcpl_630 & and_dcpl_1329 & (~
      io_read_cfg_alu_bypass_rsc_svs_st_5) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10))
      | and_dcpl_1401);
  assign FpAdd_8U_23U_and_168_cse = core_wen & ((and_dcpl_504 & and_dcpl_1329 & (~
      io_read_cfg_alu_bypass_rsc_svs_st_5) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10))
      | and_dcpl_1407);
  assign FpAdd_8U_23U_and_170_cse = core_wen & ((and_dcpl_519 & and_dcpl_1329 & (~
      io_read_cfg_alu_bypass_rsc_svs_st_5) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10))
      | and_dcpl_1413);
  assign FpAdd_8U_23U_and_172_cse = core_wen & ((and_dcpl_534 & and_dcpl_1329 & (~
      io_read_cfg_alu_bypass_rsc_svs_st_5) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10))
      | and_dcpl_1419);
  assign FpAdd_8U_23U_and_174_cse = core_wen & ((and_dcpl_549 & and_dcpl_1329 & (~
      io_read_cfg_alu_bypass_rsc_svs_st_5) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10))
      | and_dcpl_1425);
  assign nor_2190_nl = ~((cfg_alu_algo_1_sva_5[1]) | or_tmp_2842);
  assign nand_444_nl = ~((cfg_alu_algo_1_sva_5[1]) & (~ or_tmp_2842));
  assign mux_1422_nl = MUX_s_1_2_2((nand_444_nl), (nor_2190_nl), FpAlu_8U_23U_equal_tmp_1);
  assign nand_445_nl = ~(FpAlu_8U_23U_equal_tmp_1 & or_tmp_2842);
  assign mux_1423_nl = MUX_s_1_2_2((nand_445_nl), (mux_1422_nl), cfg_alu_algo_1_sva_5[0]);
  assign FpAlu_8U_23U_and_1120_cse = IsNaN_8U_23U_2_aelse_and_cse & (~ or_dcpl_678)
      & (mux_1423_nl);
  assign FpAlu_8U_23U_and_692_cse = core_wen & (~ or_dcpl_678);
  assign and_1895_rgt = (or_dcpl_14 | or_dcpl_679) & and_89_tmp;
  assign and_1899_rgt = (or_dcpl_14 | or_dcpl_681) & and_89_tmp;
  assign and_1903_rgt = (or_dcpl_14 | or_dcpl_683) & and_89_tmp;
  assign and_1907_rgt = (or_dcpl_14 | or_dcpl_686) & and_89_tmp;
  assign and_1911_rgt = (or_dcpl_14 | or_dcpl_688) & and_89_tmp;
  assign and_1921_rgt = (or_dcpl_14 | or_dcpl_692) & and_89_tmp;
  assign and_1925_rgt = (or_dcpl_14 | or_dcpl_694) & and_89_tmp;
  assign and_1929_rgt = (or_dcpl_14 | or_dcpl_696) & and_89_tmp;
  assign and_1933_rgt = (or_dcpl_14 | or_dcpl_699) & and_89_tmp;
  assign alu_loop_op_else_if_and_9_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_1_else_if_acc_itm_32_1 & and_dcpl_1468) | and_dcpl_1476);
  assign alu_loop_op_else_else_if_and_9_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_1_else_else_if_acc_itm_32_1 & and_dcpl_1477) | and_dcpl_1483);
  assign alu_loop_op_else_if_and_12_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_2_else_if_acc_1_itm_32_1 & and_dcpl_1468) | and_dcpl_1490);
  assign alu_loop_op_else_else_if_and_12_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_2_else_else_if_acc_1_itm_32_1 & and_dcpl_1477) | and_dcpl_1497);
  assign alu_loop_op_else_if_and_15_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_3_else_if_acc_itm_32_1 & and_dcpl_1468) | and_dcpl_1504);
  assign alu_loop_op_else_else_if_and_15_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_3_else_else_if_acc_itm_32_1 & and_dcpl_1477) | and_dcpl_1511);
  assign alu_loop_op_else_if_and_18_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_4_else_if_acc_1_itm_32_1 & and_dcpl_1468) | and_dcpl_1518);
  assign alu_loop_op_else_else_if_and_18_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_4_else_else_if_acc_1_itm_32_1 & and_dcpl_1477) | and_dcpl_1525);
  assign alu_loop_op_else_if_and_21_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_5_else_if_acc_itm_32_1 & and_dcpl_1468) | and_dcpl_1532);
  assign alu_loop_op_else_else_if_and_21_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_5_else_else_if_acc_itm_32_1 & and_dcpl_1477) | and_dcpl_1539);
  assign alu_loop_op_else_if_and_24_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_6_else_if_acc_1_itm_32_1 & and_dcpl_1468) | and_dcpl_1546);
  assign alu_loop_op_else_else_if_and_24_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_6_else_else_if_acc_1_itm_32_1 & and_dcpl_1477) | and_dcpl_1553);
  assign alu_loop_op_else_if_and_27_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_7_else_if_acc_itm_32_1 & and_dcpl_1468) | and_dcpl_1560);
  assign alu_loop_op_else_else_if_and_27_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_7_else_else_if_acc_itm_32_1 & and_dcpl_1477) | and_dcpl_1567);
  assign alu_loop_op_else_if_and_30_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_8_else_if_acc_1_itm_32_1 & and_dcpl_1468) | and_dcpl_1574);
  assign alu_loop_op_else_else_if_and_30_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_8_else_else_if_acc_1_itm_32_1 & and_dcpl_1477) | and_dcpl_1581);
  assign alu_loop_op_else_if_and_33_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_9_else_if_acc_itm_32_1 & and_dcpl_1468) | and_dcpl_1588);
  assign alu_loop_op_else_else_if_and_33_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_9_else_else_if_acc_itm_32_1 & and_dcpl_1477) | and_dcpl_1595);
  assign alu_loop_op_else_if_and_36_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_10_else_if_acc_1_itm_32_1 & and_dcpl_1468) | and_dcpl_1602);
  assign alu_loop_op_else_else_if_and_36_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_10_else_else_if_acc_1_itm_32_1 & and_dcpl_1477) | and_dcpl_1609);
  assign alu_loop_op_else_if_and_39_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_11_else_if_acc_itm_32_1 & and_dcpl_1468) | and_dcpl_1616);
  assign alu_loop_op_else_else_if_and_39_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_11_else_else_if_acc_itm_32_1 & and_dcpl_1477) | and_dcpl_1623);
  assign alu_loop_op_else_if_and_42_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_12_else_if_acc_1_itm_32_1 & and_dcpl_1468) | and_dcpl_1630);
  assign alu_loop_op_else_else_if_and_42_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_12_else_else_if_acc_1_itm_32_1 & and_dcpl_1477) | and_dcpl_1637);
  assign alu_loop_op_else_if_and_45_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_13_else_if_acc_itm_32_1 & and_dcpl_1468) | and_dcpl_1644);
  assign alu_loop_op_else_else_if_and_45_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_13_else_else_if_acc_itm_32_1 & and_dcpl_1477) | and_dcpl_1651);
  assign alu_loop_op_else_if_and_48_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_14_else_if_acc_1_itm_32_1 & and_dcpl_1468) | and_dcpl_1658);
  assign alu_loop_op_else_else_if_and_48_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_14_else_else_if_acc_1_itm_32_1 & and_dcpl_1477) | and_dcpl_1665);
  assign alu_loop_op_else_if_and_51_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_15_else_if_acc_itm_32_1 & and_dcpl_1468) | and_dcpl_1672);
  assign alu_loop_op_else_else_if_and_51_cse = core_wen & ((and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & alu_loop_op_15_else_else_if_acc_itm_32_1 & and_dcpl_1477) | and_dcpl_1679);
  assign alu_loop_op_else_if_and_54_cse = core_wen & ((and_dcpl_1682 & (~ (reg_cfg_alu_algo_1_sva_st_157_cse[0]))
      & alu_loop_op_16_else_if_acc_1_itm_32_1 & or_cse_2) | and_dcpl_1686);
  assign alu_loop_op_else_else_if_and_54_cse = core_wen & ((and_dcpl_1682 & nor_tmp_847
      & or_cse_2) | and_dcpl_1691);
  assign and_2163_rgt = (or_dcpl_14 | or_dcpl_295 | IsNaN_8U_23U_2_land_12_lpi_1_dfm_st_1)
      & and_89_tmp;
  assign and_2167_rgt = (or_dcpl_14 | or_dcpl_775) & and_89_tmp;
  assign and_2171_rgt = (or_dcpl_14 | or_dcpl_777) & and_89_tmp;
  assign and_2175_rgt = (or_dcpl_14 | or_dcpl_780) & and_89_tmp;
  assign and_2179_rgt = (or_dcpl_14 | or_dcpl_783) & and_89_tmp;
  assign and_2183_rgt = (or_dcpl_14 | or_dcpl_785) & and_89_tmp;
  assign alu_nan_to_zero_op_sign_and_25_cse = core_wen & FpAdd_8U_23U_is_a_greater_oelse_FpAdd_8U_23U_is_a_greater_oelse_or_21_cse
      & (~ mux_127_itm);
  assign and_2185_rgt = and_dcpl_23 & (cfg_alu_algo_1_sva_st_92==2'b10);
  assign FpCmp_8U_23U_false_if_and_48_cse = core_wen & (and_dcpl_22 | and_dcpl_34
      | and_dcpl_36 | and_2185_rgt) & (~ mux_16_itm);
  assign and_2186_rgt = and_dcpl_23 & and_dcpl_1426;
  assign FpCmp_8U_23U_false_if_and_49_cse = core_wen & (and_dcpl_22 | and_dcpl_34
      | and_dcpl_36 | and_2186_rgt) & (~ mux_16_itm);
  assign alu_nan_to_zero_op_sign_and_cse = core_wen & FpAdd_8U_23U_is_a_greater_oelse_FpAdd_8U_23U_is_a_greater_oelse_or_21_cse;
  assign and_2193_rgt = and_dcpl_126 & (cfg_alu_algo_1_sva_st_92[1]) & and_89_tmp;
  assign and_2198_rgt = and_dcpl_126 & and_dcpl_1692;
  assign or_2856_nl = (~ alu_loop_op_else_nor_tmp_16) | io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign mux_1456_cse = MUX_s_1_2_2(io_read_cfg_alu_bypass_rsc_svs_st_1, (or_2856_nl),
      cfg_alu_algo_1_sva_st_96[1]);
  assign or_2858_nl = (~ alu_loop_op_else_nor_tmp_80) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt | (~ main_stage_v_2);
  assign mux_1457_nl = MUX_s_1_2_2(or_tmp_263, (or_2858_nl), reg_cfg_alu_algo_1_sva_st_157_cse[1]);
  assign mux_1458_nl = MUX_s_1_2_2((mux_1457_nl), mux_1456_cse, and_89_tmp);
  assign IntShiftLeft_16U_6U_32U_and_48_cse = core_wen & FpAdd_8U_23U_is_a_greater_oelse_FpAdd_8U_23U_is_a_greater_oelse_or_21_cse
      & (~ (mux_1458_nl));
  assign or_2905_nl = (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt
      | (reg_cfg_alu_algo_1_sva_st_157_cse[1]) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign or_2903_nl = (~ alu_loop_op_else_nor_tmp_80) | io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign mux_1502_nl = MUX_s_1_2_2(or_tmp_263, (or_2905_nl), or_2903_nl);
  assign mux_1503_nl = MUX_s_1_2_2((mux_1502_nl), mux_1456_cse, and_89_tmp);
  assign IntShiftLeft_16U_6U_32U_and_93_cse = core_wen & FpAdd_8U_23U_is_a_greater_oelse_FpAdd_8U_23U_is_a_greater_oelse_or_21_cse
      & (~ (mux_1503_nl));
  assign IsZero_8U_23U_and_cse = core_wen & ((and_dcpl_21 & (cfg_alu_algo_rsci_d==2'b10)
      & and_91_tmp & (~ cfg_alu_bypass_rsci_d) & (fsm_output[1])) | or_tmp_3479);
  assign IntShiftLeft_16U_6U_32U_and_cse = core_wen & (~(and_dcpl_21 | io_read_cfg_alu_bypass_rsc_svs_st_1
      | (~ and_89_tmp) | (fsm_output[0])));
  assign IsZero_8U_23U_and_16_cse = core_wen & (~(or_dcpl_901 | (~ (cfg_alu_algo_rsci_d[1]))
      | (~ and_91_tmp) | cfg_alu_bypass_rsci_d | (fsm_output[0])));
  assign and_469_nl = (cfg_precision==2'b10) & (~ cfg_alu_bypass_rsci_d) & and_91_tmp
      & (fsm_output[1]);
  assign alu_loop_op_16_X_alu_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_469_nl);
  assign alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0 = (AluIn_data_sva_1[30:23])
      == ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_mx0w0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w0});
  assign nl_alu_loop_op_1_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl = conv_u2u_3_4({2'b11
      , (alu_nan_to_zero_op_expo_1_lpi_1_dfm[4])}) + 4'b1;
  assign alu_loop_op_1_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl = nl_alu_loop_op_1_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl[3:0];
  assign IsZero_5U_23U_aelse_IsZero_5U_23U_or_15_nl = (alu_nan_to_zero_op_mant_1_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_1_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_2_nl =
      MUX_v_4_2_2(4'b0000, (alu_loop_op_1_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl),
      (IsZero_5U_23U_aelse_IsZero_5U_23U_or_15_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_144_nl = MUX_v_4_2_2(({2'b1 , (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_1_sva[5:4])}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_2_nl), FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_144_nl)
      | ({{3{IsInf_5U_23U_land_1_lpi_1_dfm}}, IsInf_5U_23U_land_1_lpi_1_dfm}) | ({{3{IsNaN_5U_23U_land_1_lpi_1_dfm}},
      IsNaN_5U_23U_land_1_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_nl =
      MUX1HOT_v_4_3_2((alu_nan_to_zero_op_expo_1_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_1_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_ssc
      , IsDenorm_5U_23U_land_1_lpi_1_dfm , IsInf_5U_23U_land_1_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_nl),
      4'b1111, IsNaN_5U_23U_land_1_lpi_1_dfm);
  assign alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0 = (AluIn_data_sva_1[62:55])
      == ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_mx0w0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w0});
  assign nl_alu_loop_op_2_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl = conv_u2u_3_4({2'b11
      , (alu_nan_to_zero_op_expo_2_lpi_1_dfm[4])}) + 4'b1;
  assign alu_loop_op_2_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl = nl_alu_loop_op_2_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl[3:0];
  assign IsZero_5U_23U_aelse_IsZero_5U_23U_or_14_nl = (alu_nan_to_zero_op_mant_2_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_2_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_6_nl =
      MUX_v_4_2_2(4'b0000, (alu_loop_op_2_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl),
      (IsZero_5U_23U_aelse_IsZero_5U_23U_or_14_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_146_nl = MUX_v_4_2_2(({2'b1 , (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_2_sva[5:4])}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_6_nl), FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_146_nl)
      | ({{3{IsInf_5U_23U_land_2_lpi_1_dfm}}, IsInf_5U_23U_land_2_lpi_1_dfm}) | ({{3{IsNaN_5U_23U_land_2_lpi_1_dfm}},
      IsNaN_5U_23U_land_2_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_1_nl
      = MUX1HOT_v_4_3_2((alu_nan_to_zero_op_expo_2_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_2_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_ssc
      , IsDenorm_5U_23U_land_2_lpi_1_dfm , IsInf_5U_23U_land_2_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_1_nl),
      4'b1111, IsNaN_5U_23U_land_2_lpi_1_dfm);
  assign alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0 = (AluIn_data_sva_1[94:87])
      == ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_mx0w0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w0});
  assign nl_alu_loop_op_3_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl = conv_u2u_3_4({2'b11
      , (alu_nan_to_zero_op_expo_3_lpi_1_dfm[4])}) + 4'b1;
  assign alu_loop_op_3_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl = nl_alu_loop_op_3_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl[3:0];
  assign IsZero_5U_23U_aelse_IsZero_5U_23U_or_13_nl = (alu_nan_to_zero_op_mant_3_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_3_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_10_nl
      = MUX_v_4_2_2(4'b0000, (alu_loop_op_3_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl),
      (IsZero_5U_23U_aelse_IsZero_5U_23U_or_13_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_148_nl = MUX_v_4_2_2(({2'b1 , (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_3_sva[5:4])}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_10_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_148_nl)
      | ({{3{IsInf_5U_23U_land_3_lpi_1_dfm}}, IsInf_5U_23U_land_3_lpi_1_dfm}) | ({{3{IsNaN_5U_23U_land_3_lpi_1_dfm}},
      IsNaN_5U_23U_land_3_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_2_nl
      = MUX1HOT_v_4_3_2((alu_nan_to_zero_op_expo_3_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_3_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_ssc
      , IsDenorm_5U_23U_land_3_lpi_1_dfm , IsInf_5U_23U_land_3_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_2_nl),
      4'b1111, IsNaN_5U_23U_land_3_lpi_1_dfm);
  assign alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0 = (AluIn_data_sva_1[126:119])
      == ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_mx0w0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3_mx0w0});
  assign nl_alu_loop_op_4_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl = conv_u2u_3_4({2'b11
      , (alu_nan_to_zero_op_expo_4_lpi_1_dfm[4])}) + 4'b1;
  assign alu_loop_op_4_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl = nl_alu_loop_op_4_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl[3:0];
  assign IsZero_5U_23U_aelse_IsZero_5U_23U_or_12_nl = (alu_nan_to_zero_op_mant_4_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_4_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_14_nl
      = MUX_v_4_2_2(4'b0000, (alu_loop_op_4_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl),
      (IsZero_5U_23U_aelse_IsZero_5U_23U_or_12_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_150_nl = MUX_v_4_2_2(({2'b1 , (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_4_sva[5:4])}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_14_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_150_nl)
      | ({{3{IsInf_5U_23U_land_4_lpi_1_dfm}}, IsInf_5U_23U_land_4_lpi_1_dfm}) | ({{3{IsNaN_5U_23U_land_4_lpi_1_dfm}},
      IsNaN_5U_23U_land_4_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_3_nl
      = MUX1HOT_v_4_3_2((alu_nan_to_zero_op_expo_4_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_4_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_ssc
      , IsDenorm_5U_23U_land_4_lpi_1_dfm , IsInf_5U_23U_land_4_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_3_nl),
      4'b1111, IsNaN_5U_23U_land_4_lpi_1_dfm);
  assign alu_loop_op_5_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0 = (AluIn_data_sva_1[158:151])
      == ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_mx0w0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3_mx0w0});
  assign nl_alu_loop_op_5_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl = conv_u2u_3_4({2'b11
      , (alu_nan_to_zero_op_expo_5_lpi_1_dfm[4])}) + 4'b1;
  assign alu_loop_op_5_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl = nl_alu_loop_op_5_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl[3:0];
  assign IsZero_5U_23U_aelse_IsZero_5U_23U_or_11_nl = (alu_nan_to_zero_op_mant_5_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_5_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_18_nl
      = MUX_v_4_2_2(4'b0000, (alu_loop_op_5_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl),
      (IsZero_5U_23U_aelse_IsZero_5U_23U_or_11_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_152_nl = MUX_v_4_2_2(({2'b1 , (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_5_sva[5:4])}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_18_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_152_nl)
      | ({{3{IsInf_5U_23U_land_5_lpi_1_dfm}}, IsInf_5U_23U_land_5_lpi_1_dfm}) | ({{3{IsNaN_5U_23U_land_5_lpi_1_dfm}},
      IsNaN_5U_23U_land_5_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_4_nl
      = MUX1HOT_v_4_3_2((alu_nan_to_zero_op_expo_5_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_5_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_ssc
      , IsDenorm_5U_23U_land_5_lpi_1_dfm , IsInf_5U_23U_land_5_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_4_nl),
      4'b1111, IsNaN_5U_23U_land_5_lpi_1_dfm);
  assign alu_loop_op_6_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0 = (AluIn_data_sva_1[190:183])
      == ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_mx0w0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3_mx0w0});
  assign nl_alu_loop_op_6_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl = conv_u2u_3_4({2'b11
      , (alu_nan_to_zero_op_expo_6_lpi_1_dfm[4])}) + 4'b1;
  assign alu_loop_op_6_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl = nl_alu_loop_op_6_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl[3:0];
  assign IsZero_5U_23U_aelse_IsZero_5U_23U_or_10_nl = (alu_nan_to_zero_op_mant_6_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_6_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_22_nl
      = MUX_v_4_2_2(4'b0000, (alu_loop_op_6_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl),
      (IsZero_5U_23U_aelse_IsZero_5U_23U_or_10_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_154_nl = MUX_v_4_2_2(({2'b1 , (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_6_sva[5:4])}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_22_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_154_nl)
      | ({{3{IsInf_5U_23U_land_6_lpi_1_dfm}}, IsInf_5U_23U_land_6_lpi_1_dfm}) | ({{3{IsNaN_5U_23U_land_6_lpi_1_dfm}},
      IsNaN_5U_23U_land_6_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_5_nl
      = MUX1HOT_v_4_3_2((alu_nan_to_zero_op_expo_6_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_6_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_ssc
      , IsDenorm_5U_23U_land_6_lpi_1_dfm , IsInf_5U_23U_land_6_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_5_nl),
      4'b1111, IsNaN_5U_23U_land_6_lpi_1_dfm);
  assign alu_loop_op_7_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0 = (AluIn_data_sva_1[222:215])
      == ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_mx0w0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3_mx0w0});
  assign nl_alu_loop_op_7_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl = conv_u2u_3_4({2'b11
      , (alu_nan_to_zero_op_expo_7_lpi_1_dfm[4])}) + 4'b1;
  assign alu_loop_op_7_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl = nl_alu_loop_op_7_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl[3:0];
  assign IsZero_5U_23U_aelse_IsZero_5U_23U_or_9_nl = (alu_nan_to_zero_op_mant_7_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_7_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_26_nl
      = MUX_v_4_2_2(4'b0000, (alu_loop_op_7_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl),
      (IsZero_5U_23U_aelse_IsZero_5U_23U_or_9_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_156_nl = MUX_v_4_2_2(({2'b1 , (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_7_sva[5:4])}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_26_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_156_nl)
      | ({{3{IsInf_5U_23U_land_7_lpi_1_dfm}}, IsInf_5U_23U_land_7_lpi_1_dfm}) | ({{3{IsNaN_5U_23U_land_7_lpi_1_dfm}},
      IsNaN_5U_23U_land_7_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_6_nl
      = MUX1HOT_v_4_3_2((alu_nan_to_zero_op_expo_7_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_7_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_ssc
      , IsDenorm_5U_23U_land_7_lpi_1_dfm , IsInf_5U_23U_land_7_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_6_nl),
      4'b1111, IsNaN_5U_23U_land_7_lpi_1_dfm);
  assign alu_loop_op_8_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0 = (AluIn_data_sva_1[254:247])
      == ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_mx0w0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3_mx0w0});
  assign nl_alu_loop_op_8_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl = conv_u2u_3_4({2'b11
      , (alu_nan_to_zero_op_expo_8_lpi_1_dfm[4])}) + 4'b1;
  assign alu_loop_op_8_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl = nl_alu_loop_op_8_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl[3:0];
  assign IsZero_5U_23U_aelse_IsZero_5U_23U_or_8_nl = (alu_nan_to_zero_op_mant_8_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_8_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_30_nl
      = MUX_v_4_2_2(4'b0000, (alu_loop_op_8_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl),
      (IsZero_5U_23U_aelse_IsZero_5U_23U_or_8_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_158_nl = MUX_v_4_2_2(({2'b1 , (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_8_sva[5:4])}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_30_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_158_nl)
      | ({{3{IsInf_5U_23U_land_8_lpi_1_dfm}}, IsInf_5U_23U_land_8_lpi_1_dfm}) | ({{3{IsNaN_5U_23U_land_8_lpi_1_dfm}},
      IsNaN_5U_23U_land_8_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_7_nl
      = MUX1HOT_v_4_3_2((alu_nan_to_zero_op_expo_8_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_8_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_ssc
      , IsDenorm_5U_23U_land_8_lpi_1_dfm , IsInf_5U_23U_land_8_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_7_nl),
      4'b1111, IsNaN_5U_23U_land_8_lpi_1_dfm);
  assign alu_loop_op_9_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0 = (AluIn_data_sva_1[286:279])
      == ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_mx0w0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3_mx0w0});
  assign nl_alu_loop_op_9_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl = conv_u2u_3_4({2'b11
      , (alu_nan_to_zero_op_expo_9_lpi_1_dfm[4])}) + 4'b1;
  assign alu_loop_op_9_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl = nl_alu_loop_op_9_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl[3:0];
  assign IsZero_5U_23U_aelse_IsZero_5U_23U_or_7_nl = (alu_nan_to_zero_op_mant_9_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_9_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_34_nl
      = MUX_v_4_2_2(4'b0000, (alu_loop_op_9_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl),
      (IsZero_5U_23U_aelse_IsZero_5U_23U_or_7_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_160_nl = MUX_v_4_2_2(({2'b1 , (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_9_sva[5:4])}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_34_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_16_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_160_nl)
      | ({{3{IsInf_5U_23U_land_9_lpi_1_dfm}}, IsInf_5U_23U_land_9_lpi_1_dfm}) | ({{3{IsNaN_5U_23U_land_9_lpi_1_dfm}},
      IsNaN_5U_23U_land_9_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_8_nl
      = MUX1HOT_v_4_3_2((alu_nan_to_zero_op_expo_9_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_9_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_16_ssc
      , IsDenorm_5U_23U_land_9_lpi_1_dfm , IsInf_5U_23U_land_9_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_8_nl),
      4'b1111, IsNaN_5U_23U_land_9_lpi_1_dfm);
  assign alu_loop_op_10_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0 = (AluIn_data_sva_1[318:311])
      == ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_mx0w0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3_mx0w0});
  assign nl_alu_loop_op_10_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl = conv_u2u_3_4({2'b11
      , (alu_nan_to_zero_op_expo_10_lpi_1_dfm[4])}) + 4'b1;
  assign alu_loop_op_10_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl = nl_alu_loop_op_10_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl[3:0];
  assign IsZero_5U_23U_aelse_IsZero_5U_23U_or_6_nl = (alu_nan_to_zero_op_mant_10_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_10_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_38_nl
      = MUX_v_4_2_2(4'b0000, (alu_loop_op_10_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl),
      (IsZero_5U_23U_aelse_IsZero_5U_23U_or_6_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_162_nl = MUX_v_4_2_2(({2'b1 , (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_10_sva[5:4])}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_38_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_18_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_162_nl)
      | ({{3{IsInf_5U_23U_land_10_lpi_1_dfm}}, IsInf_5U_23U_land_10_lpi_1_dfm}) |
      ({{3{IsNaN_5U_23U_land_10_lpi_1_dfm}}, IsNaN_5U_23U_land_10_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_9_nl
      = MUX1HOT_v_4_3_2((alu_nan_to_zero_op_expo_10_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_10_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_18_ssc
      , IsDenorm_5U_23U_land_10_lpi_1_dfm , IsInf_5U_23U_land_10_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_9_nl),
      4'b1111, IsNaN_5U_23U_land_10_lpi_1_dfm);
  assign alu_loop_op_11_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0 = (AluIn_data_sva_1[350:343])
      == ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_mx0w0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3_mx0w0});
  assign nl_alu_loop_op_11_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl = conv_u2u_3_4({2'b11
      , (alu_nan_to_zero_op_expo_11_lpi_1_dfm[4])}) + 4'b1;
  assign alu_loop_op_11_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl = nl_alu_loop_op_11_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl[3:0];
  assign IsZero_5U_23U_aelse_IsZero_5U_23U_or_5_nl = (alu_nan_to_zero_op_mant_11_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_11_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_42_nl
      = MUX_v_4_2_2(4'b0000, (alu_loop_op_11_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl),
      (IsZero_5U_23U_aelse_IsZero_5U_23U_or_5_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_164_nl = MUX_v_4_2_2(({2'b1 , (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_11_sva[5:4])}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_42_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_20_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_164_nl)
      | ({{3{IsInf_5U_23U_land_11_lpi_1_dfm}}, IsInf_5U_23U_land_11_lpi_1_dfm}) |
      ({{3{IsNaN_5U_23U_land_11_lpi_1_dfm}}, IsNaN_5U_23U_land_11_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_10_nl
      = MUX1HOT_v_4_3_2((alu_nan_to_zero_op_expo_11_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_11_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_20_ssc
      , IsDenorm_5U_23U_land_11_lpi_1_dfm , IsInf_5U_23U_land_11_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_10_nl),
      4'b1111, IsNaN_5U_23U_land_11_lpi_1_dfm);
  assign alu_loop_op_12_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0 = (AluIn_data_sva_1[382:375])
      == ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_mx0w0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3_mx0w0});
  assign nl_alu_loop_op_12_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl = conv_u2u_3_4({2'b11
      , (alu_nan_to_zero_op_expo_12_lpi_1_dfm[4])}) + 4'b1;
  assign alu_loop_op_12_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl = nl_alu_loop_op_12_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl[3:0];
  assign IsZero_5U_23U_aelse_IsZero_5U_23U_or_4_nl = (alu_nan_to_zero_op_mant_12_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_12_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_46_nl
      = MUX_v_4_2_2(4'b0000, (alu_loop_op_12_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl),
      (IsZero_5U_23U_aelse_IsZero_5U_23U_or_4_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_166_nl = MUX_v_4_2_2(({2'b1 , (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_12_sva[5:4])}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_46_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_22_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_166_nl)
      | ({{3{IsInf_5U_23U_land_12_lpi_1_dfm}}, IsInf_5U_23U_land_12_lpi_1_dfm}) |
      ({{3{IsNaN_5U_23U_land_12_lpi_1_dfm}}, IsNaN_5U_23U_land_12_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_11_nl
      = MUX1HOT_v_4_3_2((alu_nan_to_zero_op_expo_12_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_12_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_22_ssc
      , IsDenorm_5U_23U_land_12_lpi_1_dfm , IsInf_5U_23U_land_12_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_11_nl),
      4'b1111, IsNaN_5U_23U_land_12_lpi_1_dfm);
  assign alu_loop_op_13_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0 = (AluIn_data_sva_1[414:407])
      == ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_mx0w0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3_mx0w0});
  assign nl_alu_loop_op_13_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl = conv_u2u_3_4({2'b11
      , (alu_nan_to_zero_op_expo_13_lpi_1_dfm[4])}) + 4'b1;
  assign alu_loop_op_13_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl = nl_alu_loop_op_13_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl[3:0];
  assign IsZero_5U_23U_aelse_IsZero_5U_23U_or_3_nl = (alu_nan_to_zero_op_mant_13_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_13_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_50_nl
      = MUX_v_4_2_2(4'b0000, (alu_loop_op_13_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl),
      (IsZero_5U_23U_aelse_IsZero_5U_23U_or_3_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_168_nl = MUX_v_4_2_2(({2'b1 , (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_13_sva[5:4])}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_50_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_24_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_168_nl)
      | ({{3{IsInf_5U_23U_land_13_lpi_1_dfm}}, IsInf_5U_23U_land_13_lpi_1_dfm}) |
      ({{3{IsNaN_5U_23U_land_13_lpi_1_dfm}}, IsNaN_5U_23U_land_13_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_12_nl
      = MUX1HOT_v_4_3_2((alu_nan_to_zero_op_expo_13_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_13_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_24_ssc
      , IsDenorm_5U_23U_land_13_lpi_1_dfm , IsInf_5U_23U_land_13_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_12_nl),
      4'b1111, IsNaN_5U_23U_land_13_lpi_1_dfm);
  assign alu_loop_op_14_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0 = (AluIn_data_sva_1[446:439])
      == ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_mx0w0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3_mx0w0});
  assign nl_alu_loop_op_14_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl = conv_u2u_3_4({2'b11
      , (alu_nan_to_zero_op_expo_14_lpi_1_dfm[4])}) + 4'b1;
  assign alu_loop_op_14_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl = nl_alu_loop_op_14_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl[3:0];
  assign IsZero_5U_23U_aelse_IsZero_5U_23U_or_2_nl = (alu_nan_to_zero_op_mant_14_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_14_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_54_nl
      = MUX_v_4_2_2(4'b0000, (alu_loop_op_14_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl),
      (IsZero_5U_23U_aelse_IsZero_5U_23U_or_2_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_170_nl = MUX_v_4_2_2(({2'b1 , (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_14_sva[5:4])}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_54_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_26_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_170_nl)
      | ({{3{IsInf_5U_23U_land_14_lpi_1_dfm}}, IsInf_5U_23U_land_14_lpi_1_dfm}) |
      ({{3{IsNaN_5U_23U_land_14_lpi_1_dfm}}, IsNaN_5U_23U_land_14_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_13_nl
      = MUX1HOT_v_4_3_2((alu_nan_to_zero_op_expo_14_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_14_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_26_ssc
      , IsDenorm_5U_23U_land_14_lpi_1_dfm , IsInf_5U_23U_land_14_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_13_nl),
      4'b1111, IsNaN_5U_23U_land_14_lpi_1_dfm);
  assign alu_loop_op_15_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0 = (AluIn_data_sva_1[478:471])
      == ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_mx0w0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3_mx0w0});
  assign nl_alu_loop_op_15_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl = conv_u2u_3_4({2'b11
      , (alu_nan_to_zero_op_expo_15_lpi_1_dfm[4])}) + 4'b1;
  assign alu_loop_op_15_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl = nl_alu_loop_op_15_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl[3:0];
  assign IsZero_5U_23U_aelse_IsZero_5U_23U_or_1_nl = (alu_nan_to_zero_op_mant_15_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_15_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_58_nl
      = MUX_v_4_2_2(4'b0000, (alu_loop_op_15_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_nl),
      (IsZero_5U_23U_aelse_IsZero_5U_23U_or_1_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_172_nl = MUX_v_4_2_2(({2'b1 , (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_15_sva[5:4])}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_58_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_28_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_172_nl)
      | ({{3{IsInf_5U_23U_land_15_lpi_1_dfm}}, IsInf_5U_23U_land_15_lpi_1_dfm}) |
      ({{3{IsNaN_5U_23U_land_15_lpi_1_dfm}}, IsNaN_5U_23U_land_15_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_14_nl
      = MUX1HOT_v_4_3_2((alu_nan_to_zero_op_expo_15_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_15_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_28_ssc
      , IsDenorm_5U_23U_land_15_lpi_1_dfm , IsInf_5U_23U_land_15_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_14_nl),
      4'b1111, IsNaN_5U_23U_land_15_lpi_1_dfm);
  assign alu_loop_op_16_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0 = (AluIn_data_sva_1[510:503])
      == ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_mx0w0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w0});
  assign nl_alu_loop_op_16_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl = conv_u2u_3_4({2'b11
      , (alu_nan_to_zero_op_expo_lpi_1_dfm[4])}) + 4'b1;
  assign alu_loop_op_16_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl = nl_alu_loop_op_16_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl[3:0];
  assign IsZero_5U_23U_aelse_IsZero_5U_23U_or_nl = (alu_nan_to_zero_op_mant_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_62_nl
      = MUX_v_4_2_2(4'b0000, (alu_loop_op_16_FpExpoWidthInc_5U_8U_23U_1U_1U_else_acc_1_nl),
      (IsZero_5U_23U_aelse_IsZero_5U_23U_or_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_174_nl = MUX_v_4_2_2(({2'b1 , (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_sva[5:4])}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_62_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_30_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_174_nl)
      | ({{3{IsInf_5U_23U_land_lpi_1_dfm}}, IsInf_5U_23U_land_lpi_1_dfm}) | ({{3{IsNaN_5U_23U_land_lpi_1_dfm}},
      IsNaN_5U_23U_land_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_15_nl
      = MUX1HOT_v_4_3_2((alu_nan_to_zero_op_expo_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_30_ssc
      , IsDenorm_5U_23U_land_lpi_1_dfm , IsInf_5U_23U_land_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_15_nl),
      4'b1111, IsNaN_5U_23U_land_lpi_1_dfm);
  assign nl_alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0 = ({1'b1 , (~ (FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0 = nl_alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0[7:0];
  assign nl_alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0 = ({1'b1 , (~ (FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0 = nl_alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0[7:0];
  assign nl_alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0 = nl_alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0[7:0];
  assign nl_alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0 = nl_alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0[7:0];
  assign nl_alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0 = ({1'b1 , (~ (FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0 = nl_alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0[7:0];
  assign nl_alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0 = ({1'b1 , (~ (FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0 = nl_alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0[7:0];
  assign nl_alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_b_right_shift_qr_4_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0 = nl_alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0[7:0];
  assign nl_alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_a_right_shift_qr_4_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0 = nl_alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0[7:0];
  assign nl_alu_loop_op_5_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0 = ({1'b1 , (~ (FpAdd_8U_23U_b_right_shift_qr_5_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign alu_loop_op_5_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0 = nl_alu_loop_op_5_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0[7:0];
  assign nl_alu_loop_op_5_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0 = ({1'b1 , (~ (FpAdd_8U_23U_a_right_shift_qr_5_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign alu_loop_op_5_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0 = nl_alu_loop_op_5_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0[7:0];
  assign nl_alu_loop_op_6_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_b_right_shift_qr_6_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_6_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0 = nl_alu_loop_op_6_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0[7:0];
  assign nl_alu_loop_op_6_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_a_right_shift_qr_6_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_6_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0 = nl_alu_loop_op_6_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0[7:0];
  assign nl_alu_loop_op_7_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0 = ({1'b1 , (~ (FpAdd_8U_23U_b_right_shift_qr_7_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign alu_loop_op_7_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0 = nl_alu_loop_op_7_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0[7:0];
  assign nl_alu_loop_op_7_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0 = ({1'b1 , (~ (FpAdd_8U_23U_a_right_shift_qr_7_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign alu_loop_op_7_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0 = nl_alu_loop_op_7_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0[7:0];
  assign nl_alu_loop_op_8_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_b_right_shift_qr_8_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_8_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0 = nl_alu_loop_op_8_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0[7:0];
  assign nl_alu_loop_op_8_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_a_right_shift_qr_8_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_8_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0 = nl_alu_loop_op_8_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0[7:0];
  assign nl_alu_loop_op_9_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0 = ({1'b1 , (~ (FpAdd_8U_23U_b_right_shift_qr_9_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign alu_loop_op_9_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0 = nl_alu_loop_op_9_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0[7:0];
  assign nl_alu_loop_op_9_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0 = ({1'b1 , (~ (FpAdd_8U_23U_a_right_shift_qr_9_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign alu_loop_op_9_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0 = nl_alu_loop_op_9_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0[7:0];
  assign nl_alu_loop_op_10_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_b_right_shift_qr_10_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_10_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0 = nl_alu_loop_op_10_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0[7:0];
  assign nl_alu_loop_op_10_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_a_right_shift_qr_10_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_10_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0 = nl_alu_loop_op_10_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0[7:0];
  assign nl_alu_loop_op_11_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_b_right_shift_qr_11_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_11_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0 = nl_alu_loop_op_11_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0[7:0];
  assign nl_alu_loop_op_11_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_a_right_shift_qr_11_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_11_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0 = nl_alu_loop_op_11_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0[7:0];
  assign nl_alu_loop_op_12_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_b_right_shift_qr_12_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_12_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0 = nl_alu_loop_op_12_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0[7:0];
  assign nl_alu_loop_op_12_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_a_right_shift_qr_12_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_12_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0 = nl_alu_loop_op_12_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0[7:0];
  assign nl_alu_loop_op_13_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_b_right_shift_qr_13_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_13_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0 = nl_alu_loop_op_13_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0[7:0];
  assign nl_alu_loop_op_13_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_a_right_shift_qr_13_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_13_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0 = nl_alu_loop_op_13_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0[7:0];
  assign nl_alu_loop_op_14_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_b_right_shift_qr_14_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_14_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0 = nl_alu_loop_op_14_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0[7:0];
  assign nl_alu_loop_op_14_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_a_right_shift_qr_14_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_14_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0 = nl_alu_loop_op_14_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0[7:0];
  assign nl_alu_loop_op_15_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_b_right_shift_qr_15_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_15_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0 = nl_alu_loop_op_15_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0[7:0];
  assign nl_alu_loop_op_15_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_a_right_shift_qr_15_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_15_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0 = nl_alu_loop_op_15_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0[7:0];
  assign nl_alu_loop_op_16_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_16_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0 = nl_alu_loop_op_16_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0[7:0];
  assign nl_alu_loop_op_16_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0 = ({1'b1 , (~
      (FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm[7:1]))}) + 8'b1101;
  assign alu_loop_op_16_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0 = nl_alu_loop_op_16_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0[7:0];
  assign FpAdd_8U_23U_o_expo_1_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_1_lpi_1_dfm_1[3:0]),
      FpAdd_8U_23U_qr_2_lpi_1_dfm_5_3_0_1, (z_out[3:0]), {(~ (FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_256 , FpAdd_8U_23U_asn_258});
  assign FpAdd_8U_23U_and_ssc = IsNaN_8U_23U_1_land_1_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_1_lpi_1_dfm_10);
  assign FpAdd_8U_23U_and_51_ssc = FpAdd_8U_23U_and_32_tmp & (~ FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0)
      & alu_loop_op_if_alu_loop_op_if_nor_cse;
  assign FpAdd_8U_23U_and_113_ssc = FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0 & alu_loop_op_if_alu_loop_op_if_nor_cse;
  assign FpNormalize_8U_49U_if_or_itm_mx0w0 = (FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_mx2[48:0]!=49'b0000000000000000000000000000000000000000000000000);
  assign nl_alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl = ({1'b1 , FpAdd_8U_23U_qr_2_lpi_1_dfm_4_7_4_1
      , (FpAdd_8U_23U_qr_2_lpi_1_dfm_4_3_0_1[3:1])}) + 8'b1;
  assign alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl = nl_alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl[7:0];
  assign alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_itm_7 = readslicef_8_1_7((alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl));
  assign FpAdd_8U_23U_o_expo_2_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_2_lpi_1_dfm_1[3:0]),
      FpAdd_8U_23U_qr_3_lpi_1_dfm_5_3_0_1, (z_out_1[3:0]), {(~ (FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_260 , FpAdd_8U_23U_asn_262});
  assign FpAdd_8U_23U_and_2_ssc = IsNaN_8U_23U_1_land_2_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_2_lpi_1_dfm_10);
  assign FpAdd_8U_23U_and_55_ssc = FpAdd_8U_23U_and_33_tmp & (~ FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0)
      & alu_loop_op_if_alu_loop_op_if_nor_1_cse;
  assign FpAdd_8U_23U_and_115_ssc = FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0 & alu_loop_op_if_alu_loop_op_if_nor_1_cse;
  assign FpNormalize_8U_49U_if_or_1_itm_mx0w0 = (FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_mx2[48:0]!=49'b0000000000000000000000000000000000000000000000000);
  assign nl_alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_2_nl = ({1'b1 , FpAdd_8U_23U_qr_3_lpi_1_dfm_4_7_4_1
      , (FpAdd_8U_23U_qr_3_lpi_1_dfm_4_3_0_1[3:1])}) + 8'b1;
  assign alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_2_nl = nl_alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_2_nl[7:0];
  assign alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_2_itm_7 = readslicef_8_1_7((alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_2_nl));
  assign FpAdd_8U_23U_o_expo_3_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_3_lpi_1_dfm_1[3:0]),
      FpAdd_8U_23U_qr_4_lpi_1_dfm_5_3_0_1, (z_out_2[3:0]), {(~ (FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_264 , FpAdd_8U_23U_asn_266});
  assign FpAdd_8U_23U_and_4_ssc = IsNaN_8U_23U_1_land_3_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_3_lpi_1_dfm_10);
  assign FpAdd_8U_23U_and_59_ssc = FpAdd_8U_23U_and_34_tmp & (~ FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0)
      & alu_loop_op_if_alu_loop_op_if_nor_2_cse;
  assign FpAdd_8U_23U_and_117_ssc = FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0 & alu_loop_op_if_alu_loop_op_if_nor_2_cse;
  assign FpNormalize_8U_49U_if_or_2_itm_mx0w0 = (FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_mx2[48:0]!=49'b0000000000000000000000000000000000000000000000000);
  assign nl_alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_1_nl = ({1'b1 , FpAdd_8U_23U_qr_4_lpi_1_dfm_4_7_4_1
      , (FpAdd_8U_23U_qr_4_lpi_1_dfm_4_3_0_1[3:1])}) + 8'b1;
  assign alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_1_nl = nl_alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_1_nl[7:0];
  assign alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_1_itm_7 = readslicef_8_1_7((alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_1_nl));
  assign FpAdd_8U_23U_o_expo_4_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_4_lpi_1_dfm_1[3:0]),
      FpAdd_8U_23U_qr_5_lpi_1_dfm_5_3_0_1, (z_out_3[3:0]), {(~ (FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_268 , FpAdd_8U_23U_asn_270});
  assign FpAdd_8U_23U_and_6_ssc = IsNaN_8U_23U_1_land_4_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_4_lpi_1_dfm_10);
  assign FpAdd_8U_23U_and_63_ssc = FpAdd_8U_23U_and_35_tmp & (~ FpAdd_8U_23U_is_inf_4_lpi_1_dfm_2_mx0)
      & alu_loop_op_if_alu_loop_op_if_nor_3_cse;
  assign FpAdd_8U_23U_and_119_ssc = FpAdd_8U_23U_is_inf_4_lpi_1_dfm_2_mx0 & alu_loop_op_if_alu_loop_op_if_nor_3_cse;
  assign FpNormalize_8U_49U_if_or_3_itm_mx0w0 = (FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_mx2[48:0]!=49'b0000000000000000000000000000000000000000000000000);
  assign nl_alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_2_nl = ({1'b1 , FpAdd_8U_23U_qr_5_lpi_1_dfm_4_7_4_1
      , (FpAdd_8U_23U_qr_5_lpi_1_dfm_4_3_0_1[3:1])}) + 8'b1;
  assign alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_2_nl = nl_alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_2_nl[7:0];
  assign alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_2_itm_7 = readslicef_8_1_7((alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_2_nl));
  assign FpAdd_8U_23U_o_expo_5_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_5_lpi_1_dfm_1[3:0]),
      FpAdd_8U_23U_qr_6_lpi_1_dfm_5_3_0_1, (z_out_4[3:0]), {(~ (FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_272 , FpAdd_8U_23U_asn_274});
  assign FpAdd_8U_23U_and_8_ssc = IsNaN_8U_23U_1_land_5_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_5_lpi_1_dfm_10);
  assign FpAdd_8U_23U_and_67_ssc = FpAdd_8U_23U_and_36_tmp & (~ FpAdd_8U_23U_is_inf_5_lpi_1_dfm_2_mx0)
      & alu_loop_op_if_alu_loop_op_if_nor_4_cse;
  assign FpAdd_8U_23U_and_121_ssc = FpAdd_8U_23U_is_inf_5_lpi_1_dfm_2_mx0 & alu_loop_op_if_alu_loop_op_if_nor_4_cse;
  assign FpNormalize_8U_49U_if_or_4_itm_mx0w0 = (FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_mx2[48:0]!=49'b0000000000000000000000000000000000000000000000000);
  assign nl_alu_loop_op_5_FpAdd_8U_23U_if_3_if_acc_1_nl = ({1'b1 , FpAdd_8U_23U_qr_6_lpi_1_dfm_4_7_4_1
      , (FpAdd_8U_23U_qr_6_lpi_1_dfm_4_3_0_1[3:1])}) + 8'b1;
  assign alu_loop_op_5_FpAdd_8U_23U_if_3_if_acc_1_nl = nl_alu_loop_op_5_FpAdd_8U_23U_if_3_if_acc_1_nl[7:0];
  assign alu_loop_op_5_FpAdd_8U_23U_if_3_if_acc_1_itm_7 = readslicef_8_1_7((alu_loop_op_5_FpAdd_8U_23U_if_3_if_acc_1_nl));
  assign FpAdd_8U_23U_o_expo_6_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_6_lpi_1_dfm_1[3:0]),
      FpAdd_8U_23U_qr_7_lpi_1_dfm_5_3_0_1, (z_out_5[3:0]), {(~ (FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_276 , FpAdd_8U_23U_asn_278});
  assign FpAdd_8U_23U_and_10_ssc = IsNaN_8U_23U_1_land_6_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_6_lpi_1_dfm_10);
  assign FpAdd_8U_23U_and_71_ssc = FpAdd_8U_23U_and_37_tmp & (~ FpAdd_8U_23U_is_inf_6_lpi_1_dfm_2_mx0)
      & alu_loop_op_if_alu_loop_op_if_nor_5_cse;
  assign FpAdd_8U_23U_and_123_ssc = FpAdd_8U_23U_is_inf_6_lpi_1_dfm_2_mx0 & alu_loop_op_if_alu_loop_op_if_nor_5_cse;
  assign FpNormalize_8U_49U_if_or_5_itm_mx0w0 = (FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_mx2[48:0]!=49'b0000000000000000000000000000000000000000000000000);
  assign nl_alu_loop_op_6_FpAdd_8U_23U_if_3_if_acc_2_nl = ({1'b1 , FpAdd_8U_23U_qr_7_lpi_1_dfm_4_7_4_1
      , (FpAdd_8U_23U_qr_7_lpi_1_dfm_4_3_0_1[3:1])}) + 8'b1;
  assign alu_loop_op_6_FpAdd_8U_23U_if_3_if_acc_2_nl = nl_alu_loop_op_6_FpAdd_8U_23U_if_3_if_acc_2_nl[7:0];
  assign alu_loop_op_6_FpAdd_8U_23U_if_3_if_acc_2_itm_7 = readslicef_8_1_7((alu_loop_op_6_FpAdd_8U_23U_if_3_if_acc_2_nl));
  assign FpAdd_8U_23U_o_expo_7_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_7_lpi_1_dfm_1[3:0]),
      FpAdd_8U_23U_qr_8_lpi_1_dfm_5_3_0_1, (z_out_6[3:0]), {(~ (FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_280 , FpAdd_8U_23U_asn_282});
  assign FpAdd_8U_23U_and_12_ssc = IsNaN_8U_23U_1_land_7_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_7_lpi_1_dfm_10);
  assign FpAdd_8U_23U_and_75_ssc = FpAdd_8U_23U_and_38_tmp & (~ FpAdd_8U_23U_is_inf_7_lpi_1_dfm_2_mx0)
      & alu_loop_op_if_alu_loop_op_if_nor_6_cse;
  assign FpAdd_8U_23U_and_125_ssc = FpAdd_8U_23U_is_inf_7_lpi_1_dfm_2_mx0 & alu_loop_op_if_alu_loop_op_if_nor_6_cse;
  assign FpNormalize_8U_49U_if_or_6_itm_mx0w0 = (FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_mx2[48:0]!=49'b0000000000000000000000000000000000000000000000000);
  assign nl_alu_loop_op_7_FpAdd_8U_23U_if_3_if_acc_1_nl = ({1'b1 , FpAdd_8U_23U_qr_8_lpi_1_dfm_4_7_4_1
      , (FpAdd_8U_23U_qr_8_lpi_1_dfm_4_3_0_1[3:1])}) + 8'b1;
  assign alu_loop_op_7_FpAdd_8U_23U_if_3_if_acc_1_nl = nl_alu_loop_op_7_FpAdd_8U_23U_if_3_if_acc_1_nl[7:0];
  assign alu_loop_op_7_FpAdd_8U_23U_if_3_if_acc_1_itm_7 = readslicef_8_1_7((alu_loop_op_7_FpAdd_8U_23U_if_3_if_acc_1_nl));
  assign FpAdd_8U_23U_o_expo_8_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_8_lpi_1_dfm_1[3:0]),
      FpAdd_8U_23U_qr_9_lpi_1_dfm_5_3_0_1, (z_out_7[3:0]), {(~ (FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_284 , FpAdd_8U_23U_asn_286});
  assign FpAdd_8U_23U_and_14_ssc = IsNaN_8U_23U_1_land_8_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_8_lpi_1_dfm_10);
  assign FpAdd_8U_23U_and_79_ssc = FpAdd_8U_23U_and_39_tmp & (~ FpAdd_8U_23U_is_inf_8_lpi_1_dfm_2_mx0)
      & alu_loop_op_if_alu_loop_op_if_nor_7_cse;
  assign FpAdd_8U_23U_and_127_ssc = FpAdd_8U_23U_is_inf_8_lpi_1_dfm_2_mx0 & alu_loop_op_if_alu_loop_op_if_nor_7_cse;
  assign FpNormalize_8U_49U_if_or_7_itm_mx0w0 = (FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_mx2[48:0]!=49'b0000000000000000000000000000000000000000000000000);
  assign nl_alu_loop_op_8_FpAdd_8U_23U_if_3_if_acc_2_nl = ({1'b1 , FpAdd_8U_23U_qr_9_lpi_1_dfm_4_7_4_1
      , (FpAdd_8U_23U_qr_9_lpi_1_dfm_4_3_0_1[3:1])}) + 8'b1;
  assign alu_loop_op_8_FpAdd_8U_23U_if_3_if_acc_2_nl = nl_alu_loop_op_8_FpAdd_8U_23U_if_3_if_acc_2_nl[7:0];
  assign alu_loop_op_8_FpAdd_8U_23U_if_3_if_acc_2_itm_7 = readslicef_8_1_7((alu_loop_op_8_FpAdd_8U_23U_if_3_if_acc_2_nl));
  assign FpAdd_8U_23U_o_expo_9_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_9_lpi_1_dfm_1[3:0]),
      FpAdd_8U_23U_qr_10_lpi_1_dfm_5_3_0_1, (z_out_8[3:0]), {(~ (FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_288 , FpAdd_8U_23U_asn_290});
  assign FpAdd_8U_23U_and_16_ssc = IsNaN_8U_23U_1_land_9_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_9_lpi_1_dfm_10);
  assign FpAdd_8U_23U_and_83_ssc = FpAdd_8U_23U_and_40_tmp & (~ FpAdd_8U_23U_is_inf_9_lpi_1_dfm_2_mx0)
      & alu_loop_op_if_alu_loop_op_if_nor_8_cse;
  assign FpAdd_8U_23U_and_129_ssc = FpAdd_8U_23U_is_inf_9_lpi_1_dfm_2_mx0 & alu_loop_op_if_alu_loop_op_if_nor_8_cse;
  assign FpNormalize_8U_49U_if_or_8_itm_mx0w0 = (FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_mx2[48:0]!=49'b0000000000000000000000000000000000000000000000000);
  assign nl_alu_loop_op_9_FpAdd_8U_23U_if_3_if_acc_1_nl = ({1'b1 , FpAdd_8U_23U_qr_10_lpi_1_dfm_4_7_4_1
      , (FpAdd_8U_23U_qr_10_lpi_1_dfm_4_3_0_1[3:1])}) + 8'b1;
  assign alu_loop_op_9_FpAdd_8U_23U_if_3_if_acc_1_nl = nl_alu_loop_op_9_FpAdd_8U_23U_if_3_if_acc_1_nl[7:0];
  assign alu_loop_op_9_FpAdd_8U_23U_if_3_if_acc_1_itm_7 = readslicef_8_1_7((alu_loop_op_9_FpAdd_8U_23U_if_3_if_acc_1_nl));
  assign FpAdd_8U_23U_o_expo_10_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_10_lpi_1_dfm_1[3:0]),
      FpAdd_8U_23U_qr_11_lpi_1_dfm_5_3_0_1, (z_out_9[3:0]), {(~ (FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_292 , FpAdd_8U_23U_asn_294});
  assign FpAdd_8U_23U_and_18_ssc = IsNaN_8U_23U_1_land_10_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_10_lpi_1_dfm_10);
  assign FpAdd_8U_23U_and_87_ssc = FpAdd_8U_23U_and_41_tmp & (~ FpAdd_8U_23U_is_inf_10_lpi_1_dfm_2_mx0)
      & alu_loop_op_if_alu_loop_op_if_nor_9_cse;
  assign FpAdd_8U_23U_and_131_ssc = FpAdd_8U_23U_is_inf_10_lpi_1_dfm_2_mx0 & alu_loop_op_if_alu_loop_op_if_nor_9_cse;
  assign FpNormalize_8U_49U_if_or_9_itm_mx0w0 = (FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_mx2[48:0]!=49'b0000000000000000000000000000000000000000000000000);
  assign nl_alu_loop_op_10_FpAdd_8U_23U_if_3_if_acc_2_nl = ({1'b1 , FpAdd_8U_23U_qr_11_lpi_1_dfm_4_7_4_1
      , (FpAdd_8U_23U_qr_11_lpi_1_dfm_4_3_0_1[3:1])}) + 8'b1;
  assign alu_loop_op_10_FpAdd_8U_23U_if_3_if_acc_2_nl = nl_alu_loop_op_10_FpAdd_8U_23U_if_3_if_acc_2_nl[7:0];
  assign alu_loop_op_10_FpAdd_8U_23U_if_3_if_acc_2_itm_7 = readslicef_8_1_7((alu_loop_op_10_FpAdd_8U_23U_if_3_if_acc_2_nl));
  assign FpAdd_8U_23U_o_expo_11_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_11_lpi_1_dfm_1[3:0]),
      FpAdd_8U_23U_qr_12_lpi_1_dfm_5_3_0_1, (z_out_10[3:0]), {(~ (FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_296 , FpAdd_8U_23U_asn_298});
  assign FpAdd_8U_23U_and_20_ssc = IsNaN_8U_23U_1_land_11_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_11_lpi_1_dfm_10);
  assign FpAdd_8U_23U_and_91_ssc = FpAdd_8U_23U_and_42_tmp & (~ FpAdd_8U_23U_is_inf_11_lpi_1_dfm_2_mx0)
      & alu_loop_op_if_alu_loop_op_if_nor_10_cse;
  assign FpAdd_8U_23U_and_133_ssc = FpAdd_8U_23U_is_inf_11_lpi_1_dfm_2_mx0 & alu_loop_op_if_alu_loop_op_if_nor_10_cse;
  assign FpNormalize_8U_49U_if_or_10_itm_mx0w0 = (FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_mx2[48:0]!=49'b0000000000000000000000000000000000000000000000000);
  assign nl_alu_loop_op_11_FpAdd_8U_23U_if_3_if_acc_1_nl = ({1'b1 , FpAdd_8U_23U_qr_12_lpi_1_dfm_4_7_4_1
      , (FpAdd_8U_23U_qr_12_lpi_1_dfm_4_3_0_1[3:1])}) + 8'b1;
  assign alu_loop_op_11_FpAdd_8U_23U_if_3_if_acc_1_nl = nl_alu_loop_op_11_FpAdd_8U_23U_if_3_if_acc_1_nl[7:0];
  assign alu_loop_op_11_FpAdd_8U_23U_if_3_if_acc_1_itm_7 = readslicef_8_1_7((alu_loop_op_11_FpAdd_8U_23U_if_3_if_acc_1_nl));
  assign FpAdd_8U_23U_o_expo_12_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_12_lpi_1_dfm_1[3:0]),
      FpAdd_8U_23U_qr_13_lpi_1_dfm_5_3_0_1, (z_out_11[3:0]), {(~ (FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_300 , FpAdd_8U_23U_asn_302});
  assign FpAdd_8U_23U_and_22_ssc = IsNaN_8U_23U_1_land_12_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_12_lpi_1_dfm_10);
  assign FpAdd_8U_23U_and_95_ssc = FpAdd_8U_23U_and_43_tmp & (~ FpAdd_8U_23U_is_inf_12_lpi_1_dfm_2_mx0)
      & alu_loop_op_if_alu_loop_op_if_nor_11_cse;
  assign FpAdd_8U_23U_and_135_ssc = FpAdd_8U_23U_is_inf_12_lpi_1_dfm_2_mx0 & alu_loop_op_if_alu_loop_op_if_nor_11_cse;
  assign FpNormalize_8U_49U_if_or_11_itm_mx0w0 = (FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_mx2[48:0]!=49'b0000000000000000000000000000000000000000000000000);
  assign nl_alu_loop_op_12_FpAdd_8U_23U_if_3_if_acc_2_nl = ({1'b1 , FpAdd_8U_23U_qr_13_lpi_1_dfm_4_7_4_1
      , (FpAdd_8U_23U_qr_13_lpi_1_dfm_4_3_0_1[3:1])}) + 8'b1;
  assign alu_loop_op_12_FpAdd_8U_23U_if_3_if_acc_2_nl = nl_alu_loop_op_12_FpAdd_8U_23U_if_3_if_acc_2_nl[7:0];
  assign alu_loop_op_12_FpAdd_8U_23U_if_3_if_acc_2_itm_7 = readslicef_8_1_7((alu_loop_op_12_FpAdd_8U_23U_if_3_if_acc_2_nl));
  assign FpAdd_8U_23U_o_expo_13_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_13_lpi_1_dfm_1[3:0]),
      FpAdd_8U_23U_qr_14_lpi_1_dfm_5_3_0_1, (z_out_12[3:0]), {(~ (FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_304 , FpAdd_8U_23U_asn_306});
  assign FpAdd_8U_23U_and_24_ssc = IsNaN_8U_23U_1_land_13_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_13_lpi_1_dfm_10);
  assign FpAdd_8U_23U_and_99_ssc = FpAdd_8U_23U_and_44_tmp & (~ FpAdd_8U_23U_is_inf_13_lpi_1_dfm_2_mx0)
      & alu_loop_op_if_alu_loop_op_if_nor_12_cse;
  assign FpAdd_8U_23U_and_137_ssc = FpAdd_8U_23U_is_inf_13_lpi_1_dfm_2_mx0 & alu_loop_op_if_alu_loop_op_if_nor_12_cse;
  assign FpNormalize_8U_49U_if_or_12_itm_mx0w0 = (FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_mx2[48:0]!=49'b0000000000000000000000000000000000000000000000000);
  assign nl_alu_loop_op_13_FpAdd_8U_23U_if_3_if_acc_1_nl = ({1'b1 , FpAdd_8U_23U_qr_14_lpi_1_dfm_4_7_4_1
      , (FpAdd_8U_23U_qr_14_lpi_1_dfm_4_3_0_1[3:1])}) + 8'b1;
  assign alu_loop_op_13_FpAdd_8U_23U_if_3_if_acc_1_nl = nl_alu_loop_op_13_FpAdd_8U_23U_if_3_if_acc_1_nl[7:0];
  assign alu_loop_op_13_FpAdd_8U_23U_if_3_if_acc_1_itm_7 = readslicef_8_1_7((alu_loop_op_13_FpAdd_8U_23U_if_3_if_acc_1_nl));
  assign FpAdd_8U_23U_o_expo_14_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_14_lpi_1_dfm_1[3:0]),
      FpAdd_8U_23U_qr_15_lpi_1_dfm_5_3_0_1, (z_out_13[3:0]), {(~ (FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_308 , FpAdd_8U_23U_asn_310});
  assign FpAdd_8U_23U_and_26_ssc = IsNaN_8U_23U_1_land_14_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_14_lpi_1_dfm_10);
  assign FpAdd_8U_23U_and_103_ssc = FpAdd_8U_23U_and_45_tmp & (~ FpAdd_8U_23U_is_inf_14_lpi_1_dfm_2_mx0)
      & alu_loop_op_if_alu_loop_op_if_nor_13_cse;
  assign FpAdd_8U_23U_and_139_ssc = FpAdd_8U_23U_is_inf_14_lpi_1_dfm_2_mx0 & alu_loop_op_if_alu_loop_op_if_nor_13_cse;
  assign FpNormalize_8U_49U_if_or_13_itm_mx0w0 = (FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_mx2[48:0]!=49'b0000000000000000000000000000000000000000000000000);
  assign nl_alu_loop_op_14_FpAdd_8U_23U_if_3_if_acc_2_nl = ({1'b1 , FpAdd_8U_23U_qr_15_lpi_1_dfm_4_7_4_1
      , (FpAdd_8U_23U_qr_15_lpi_1_dfm_4_3_0_1[3:1])}) + 8'b1;
  assign alu_loop_op_14_FpAdd_8U_23U_if_3_if_acc_2_nl = nl_alu_loop_op_14_FpAdd_8U_23U_if_3_if_acc_2_nl[7:0];
  assign alu_loop_op_14_FpAdd_8U_23U_if_3_if_acc_2_itm_7 = readslicef_8_1_7((alu_loop_op_14_FpAdd_8U_23U_if_3_if_acc_2_nl));
  assign FpAdd_8U_23U_o_expo_15_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_15_lpi_1_dfm_1[3:0]),
      FpAdd_8U_23U_qr_16_lpi_1_dfm_5_3_0_1, (z_out_14[3:0]), {(~ (FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_312 , FpAdd_8U_23U_asn_314});
  assign FpAdd_8U_23U_and_28_ssc = IsNaN_8U_23U_1_land_15_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_15_lpi_1_dfm_10);
  assign FpAdd_8U_23U_and_107_ssc = FpAdd_8U_23U_and_46_tmp & (~ FpAdd_8U_23U_is_inf_15_lpi_1_dfm_2_mx0)
      & alu_loop_op_if_alu_loop_op_if_nor_14_cse;
  assign FpAdd_8U_23U_and_141_ssc = FpAdd_8U_23U_is_inf_15_lpi_1_dfm_2_mx0 & alu_loop_op_if_alu_loop_op_if_nor_14_cse;
  assign FpNormalize_8U_49U_if_or_14_itm_mx0w0 = (FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_mx2[48:0]!=49'b0000000000000000000000000000000000000000000000000);
  assign nl_alu_loop_op_15_FpAdd_8U_23U_if_3_if_acc_1_nl = ({1'b1 , FpAdd_8U_23U_qr_16_lpi_1_dfm_4_7_4_1
      , (FpAdd_8U_23U_qr_16_lpi_1_dfm_4_3_0_1[3:1])}) + 8'b1;
  assign alu_loop_op_15_FpAdd_8U_23U_if_3_if_acc_1_nl = nl_alu_loop_op_15_FpAdd_8U_23U_if_3_if_acc_1_nl[7:0];
  assign alu_loop_op_15_FpAdd_8U_23U_if_3_if_acc_1_itm_7 = readslicef_8_1_7((alu_loop_op_15_FpAdd_8U_23U_if_3_if_acc_1_nl));
  assign FpAdd_8U_23U_o_expo_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_lpi_1_dfm_1[3:0]),
      FpAdd_8U_23U_qr_lpi_1_dfm_5_3_0_1, (z_out_15[3:0]), {(~ (FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_316 , FpAdd_8U_23U_asn_318});
  assign FpAdd_8U_23U_and_30_ssc = IsNaN_8U_23U_1_land_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_lpi_1_dfm_10);
  assign FpAdd_8U_23U_and_111_ssc = FpAdd_8U_23U_and_47_tmp & (~ FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0)
      & alu_loop_op_if_alu_loop_op_if_nor_15_cse;
  assign FpAdd_8U_23U_and_143_ssc = FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0 & alu_loop_op_if_alu_loop_op_if_nor_15_cse;
  assign FpNormalize_8U_49U_if_or_15_itm_mx0w0 = (FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_mx2[48:0]!=49'b0000000000000000000000000000000000000000000000000);
  assign nl_alu_loop_op_16_FpAdd_8U_23U_if_3_if_acc_2_nl = ({1'b1 , FpAdd_8U_23U_qr_lpi_1_dfm_4_7_4_1
      , (FpAdd_8U_23U_qr_lpi_1_dfm_4_3_0_1[3:1])}) + 8'b1;
  assign alu_loop_op_16_FpAdd_8U_23U_if_3_if_acc_2_nl = nl_alu_loop_op_16_FpAdd_8U_23U_if_3_if_acc_2_nl[7:0];
  assign alu_loop_op_16_FpAdd_8U_23U_if_3_if_acc_2_itm_7 = readslicef_8_1_7((alu_loop_op_16_FpAdd_8U_23U_if_3_if_acc_2_nl));
  assign nl_FpAdd_8U_23U_asn_76_mx1w1 = ({1'b1 , (~ FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_mx0) + 50'b1;
  assign FpAdd_8U_23U_asn_76_mx1w1 = nl_FpAdd_8U_23U_asn_76_mx1w1[49:0];
  assign and_876_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & reg_alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign and_878_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & (~ reg_alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse)
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_mx1 = MUX1HOT_v_50_3_2(FpAdd_8U_23U_int_mant_p1_1_sva,
      FpAdd_8U_23U_asn_76_mx1w1, FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm, {(and_876_nl)
      , (and_878_nl) , or_334_cse});
  assign FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_mx2 = MUX_v_50_2_2(FpAdd_8U_23U_asn_76_mx1w1,
      FpAdd_8U_23U_int_mant_p1_1_sva, reg_alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse);
  assign nl_FpAdd_8U_23U_asn_73_mx1w1 = ({1'b1 , (~ FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_mx0) + 50'b1;
  assign FpAdd_8U_23U_asn_73_mx1w1 = nl_FpAdd_8U_23U_asn_73_mx1w1[49:0];
  assign and_891_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & reg_alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign and_893_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & (~ reg_alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse)
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_mx1 = MUX1HOT_v_50_3_2(FpAdd_8U_23U_int_mant_p1_2_sva,
      FpAdd_8U_23U_asn_73_mx1w1, FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm, {(and_891_nl)
      , (and_893_nl) , or_334_cse});
  assign FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_mx2 = MUX_v_50_2_2(FpAdd_8U_23U_asn_73_mx1w1,
      FpAdd_8U_23U_int_mant_p1_2_sva, reg_alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse);
  assign nl_FpAdd_8U_23U_asn_70_mx1w1 = ({1'b1 , (~ FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_mx0) + 50'b1;
  assign FpAdd_8U_23U_asn_70_mx1w1 = nl_FpAdd_8U_23U_asn_70_mx1w1[49:0];
  assign and_906_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & reg_alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign and_908_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & (~ reg_alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse)
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_mx1 = MUX1HOT_v_50_3_2(FpAdd_8U_23U_int_mant_p1_3_sva,
      FpAdd_8U_23U_asn_70_mx1w1, FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm, {(and_906_nl)
      , (and_908_nl) , or_334_cse});
  assign FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_mx2 = MUX_v_50_2_2(FpAdd_8U_23U_asn_70_mx1w1,
      FpAdd_8U_23U_int_mant_p1_3_sva, reg_alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse);
  assign nl_FpAdd_8U_23U_asn_67_mx1w1 = ({1'b1 , (~ FpAdd_8U_23U_addend_smaller_qr_4_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_4_lpi_1_dfm_mx0) + 50'b1;
  assign FpAdd_8U_23U_asn_67_mx1w1 = nl_FpAdd_8U_23U_asn_67_mx1w1[49:0];
  assign and_921_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & reg_alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign and_923_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & (~ reg_alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse)
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_mx1 = MUX1HOT_v_50_3_2(FpAdd_8U_23U_int_mant_p1_4_sva,
      FpAdd_8U_23U_asn_67_mx1w1, FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm, {(and_921_nl)
      , (and_923_nl) , or_334_cse});
  assign FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_mx2 = MUX_v_50_2_2(FpAdd_8U_23U_asn_67_mx1w1,
      FpAdd_8U_23U_int_mant_p1_4_sva, reg_alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse);
  assign nl_FpAdd_8U_23U_asn_64_mx1w1 = ({1'b1 , (~ FpAdd_8U_23U_addend_smaller_qr_5_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_5_lpi_1_dfm_mx0) + 50'b1;
  assign FpAdd_8U_23U_asn_64_mx1w1 = nl_FpAdd_8U_23U_asn_64_mx1w1[49:0];
  assign and_925_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & reg_alu_loop_op_5_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign and_927_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & (~ reg_alu_loop_op_5_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse)
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_mx1 = MUX1HOT_v_50_3_2(FpAdd_8U_23U_int_mant_p1_5_sva,
      FpAdd_8U_23U_asn_64_mx1w1, FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm, {(and_925_nl)
      , (and_927_nl) , or_334_cse});
  assign FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_mx2 = MUX_v_50_2_2(FpAdd_8U_23U_asn_64_mx1w1,
      FpAdd_8U_23U_int_mant_p1_5_sva, reg_alu_loop_op_5_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse);
  assign nl_FpAdd_8U_23U_asn_61_mx1w1 = ({1'b1 , (~ FpAdd_8U_23U_addend_smaller_qr_6_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_6_lpi_1_dfm_mx0) + 50'b1;
  assign FpAdd_8U_23U_asn_61_mx1w1 = nl_FpAdd_8U_23U_asn_61_mx1w1[49:0];
  assign and_929_nl = reg_alu_loop_op_6_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
      & (cfg_alu_algo_1_sva_st_204==2'b10);
  assign and_931_nl = (~ reg_alu_loop_op_6_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse)
      & (cfg_alu_algo_1_sva_st_204==2'b10);
  assign FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_mx1 = MUX1HOT_v_50_3_2(FpAdd_8U_23U_int_mant_p1_6_sva,
      FpAdd_8U_23U_asn_61_mx1w1, FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm, {(and_929_nl)
      , (and_931_nl) , or_334_cse});
  assign FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_mx2 = MUX_v_50_2_2(FpAdd_8U_23U_asn_61_mx1w1,
      FpAdd_8U_23U_int_mant_p1_6_sva, reg_alu_loop_op_6_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse);
  assign nl_FpAdd_8U_23U_asn_58_mx1w1 = ({1'b1 , (~ FpAdd_8U_23U_addend_smaller_qr_7_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_7_lpi_1_dfm_mx0) + 50'b1;
  assign FpAdd_8U_23U_asn_58_mx1w1 = nl_FpAdd_8U_23U_asn_58_mx1w1[49:0];
  assign and_933_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & reg_alu_loop_op_7_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign and_935_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & (~ reg_alu_loop_op_7_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse)
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_mx1 = MUX1HOT_v_50_3_2(FpAdd_8U_23U_int_mant_p1_7_sva,
      FpAdd_8U_23U_asn_58_mx1w1, FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm, {(and_933_nl)
      , (and_935_nl) , or_334_cse});
  assign FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_mx2 = MUX_v_50_2_2(FpAdd_8U_23U_asn_58_mx1w1,
      FpAdd_8U_23U_int_mant_p1_7_sva, reg_alu_loop_op_7_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse);
  assign nl_FpAdd_8U_23U_asn_55_mx1w1 = ({1'b1 , (~ FpAdd_8U_23U_addend_smaller_qr_8_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_8_lpi_1_dfm_mx0) + 50'b1;
  assign FpAdd_8U_23U_asn_55_mx1w1 = nl_FpAdd_8U_23U_asn_55_mx1w1[49:0];
  assign and_948_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & reg_alu_loop_op_8_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign and_950_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & (~ reg_alu_loop_op_8_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse)
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_mx1 = MUX1HOT_v_50_3_2(FpAdd_8U_23U_int_mant_p1_8_sva,
      FpAdd_8U_23U_asn_55_mx1w1, FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm, {(and_948_nl)
      , (and_950_nl) , or_334_cse});
  assign FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_mx2 = MUX_v_50_2_2(FpAdd_8U_23U_asn_55_mx1w1,
      FpAdd_8U_23U_int_mant_p1_8_sva, reg_alu_loop_op_8_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse);
  assign nl_FpAdd_8U_23U_asn_52_mx1w1 = ({1'b1 , (~ FpAdd_8U_23U_addend_smaller_qr_9_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_9_lpi_1_dfm_mx0) + 50'b1;
  assign FpAdd_8U_23U_asn_52_mx1w1 = nl_FpAdd_8U_23U_asn_52_mx1w1[49:0];
  assign and_952_nl = reg_alu_loop_op_9_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
      & (cfg_alu_algo_1_sva_st_204==2'b10);
  assign and_954_nl = (~ reg_alu_loop_op_9_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse)
      & (cfg_alu_algo_1_sva_st_204==2'b10);
  assign FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_mx1 = MUX1HOT_v_50_3_2(FpAdd_8U_23U_int_mant_p1_9_sva,
      FpAdd_8U_23U_asn_52_mx1w1, FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm, {(and_952_nl)
      , (and_954_nl) , or_334_cse});
  assign FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_mx2 = MUX_v_50_2_2(FpAdd_8U_23U_asn_52_mx1w1,
      FpAdd_8U_23U_int_mant_p1_9_sva, reg_alu_loop_op_9_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse);
  assign nl_FpAdd_8U_23U_asn_49_mx1w1 = ({1'b1 , (~ FpAdd_8U_23U_addend_smaller_qr_10_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_10_lpi_1_dfm_mx0) + 50'b1;
  assign FpAdd_8U_23U_asn_49_mx1w1 = nl_FpAdd_8U_23U_asn_49_mx1w1[49:0];
  assign and_956_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & reg_alu_loop_op_10_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign and_958_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & (~ reg_alu_loop_op_10_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse)
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_mx1 = MUX1HOT_v_50_3_2(FpAdd_8U_23U_int_mant_p1_10_sva,
      FpAdd_8U_23U_asn_49_mx1w1, FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm, {(and_956_nl)
      , (and_958_nl) , or_334_cse});
  assign FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_mx2 = MUX_v_50_2_2(FpAdd_8U_23U_asn_49_mx1w1,
      FpAdd_8U_23U_int_mant_p1_10_sva, reg_alu_loop_op_10_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse);
  assign nl_FpAdd_8U_23U_asn_46_mx1w1 = ({1'b1 , (~ FpAdd_8U_23U_addend_smaller_qr_11_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_11_lpi_1_dfm_mx0) + 50'b1;
  assign FpAdd_8U_23U_asn_46_mx1w1 = nl_FpAdd_8U_23U_asn_46_mx1w1[49:0];
  assign and_960_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & reg_alu_loop_op_11_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign and_962_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & (~ reg_alu_loop_op_11_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse)
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_mx1 = MUX1HOT_v_50_3_2(FpAdd_8U_23U_int_mant_p1_11_sva,
      FpAdd_8U_23U_asn_46_mx1w1, FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm, {(and_960_nl)
      , (and_962_nl) , or_334_cse});
  assign FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_mx2 = MUX_v_50_2_2(FpAdd_8U_23U_asn_46_mx1w1,
      FpAdd_8U_23U_int_mant_p1_11_sva, reg_alu_loop_op_11_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse);
  assign nl_FpAdd_8U_23U_asn_43_mx1w1 = ({1'b1 , (~ FpAdd_8U_23U_addend_smaller_qr_12_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_12_lpi_1_dfm_mx0) + 50'b1;
  assign FpAdd_8U_23U_asn_43_mx1w1 = nl_FpAdd_8U_23U_asn_43_mx1w1[49:0];
  assign and_964_nl = reg_alu_loop_op_12_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
      & (cfg_alu_algo_1_sva_st_204==2'b10);
  assign and_966_nl = (~ reg_alu_loop_op_12_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse)
      & (cfg_alu_algo_1_sva_st_204==2'b10);
  assign FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_mx1 = MUX1HOT_v_50_3_2(FpAdd_8U_23U_int_mant_p1_12_sva,
      FpAdd_8U_23U_asn_43_mx1w1, FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm, {(and_964_nl)
      , (and_966_nl) , or_334_cse});
  assign FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_mx2 = MUX_v_50_2_2(FpAdd_8U_23U_asn_43_mx1w1,
      FpAdd_8U_23U_int_mant_p1_12_sva, reg_alu_loop_op_12_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse);
  assign nl_FpAdd_8U_23U_asn_40_mx1w1 = ({1'b1 , (~ FpAdd_8U_23U_addend_smaller_qr_13_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_13_lpi_1_dfm_mx0) + 50'b1;
  assign FpAdd_8U_23U_asn_40_mx1w1 = nl_FpAdd_8U_23U_asn_40_mx1w1[49:0];
  assign and_979_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & reg_alu_loop_op_13_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign and_981_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & (~ reg_alu_loop_op_13_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse)
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_mx1 = MUX1HOT_v_50_3_2(FpAdd_8U_23U_int_mant_p1_13_sva,
      FpAdd_8U_23U_asn_40_mx1w1, FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm, {(and_979_nl)
      , (and_981_nl) , or_334_cse});
  assign FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_mx2 = MUX_v_50_2_2(FpAdd_8U_23U_asn_40_mx1w1,
      FpAdd_8U_23U_int_mant_p1_13_sva, reg_alu_loop_op_13_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse);
  assign nl_FpAdd_8U_23U_asn_37_mx1w1 = ({1'b1 , (~ FpAdd_8U_23U_addend_smaller_qr_14_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_14_lpi_1_dfm_mx0) + 50'b1;
  assign FpAdd_8U_23U_asn_37_mx1w1 = nl_FpAdd_8U_23U_asn_37_mx1w1[49:0];
  assign and_994_nl = reg_alu_loop_op_14_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
      & (cfg_alu_algo_1_sva_st_204==2'b10);
  assign and_996_nl = (~ reg_alu_loop_op_14_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse)
      & (cfg_alu_algo_1_sva_st_204==2'b10);
  assign FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_mx1 = MUX1HOT_v_50_3_2(FpAdd_8U_23U_int_mant_p1_14_sva,
      FpAdd_8U_23U_asn_37_mx1w1, FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm, {(and_994_nl)
      , (and_996_nl) , or_334_cse});
  assign FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_mx2 = MUX_v_50_2_2(FpAdd_8U_23U_asn_37_mx1w1,
      FpAdd_8U_23U_int_mant_p1_14_sva, reg_alu_loop_op_14_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse);
  assign nl_FpAdd_8U_23U_asn_34_mx1w1 = ({1'b1 , (~ FpAdd_8U_23U_addend_smaller_qr_15_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_15_lpi_1_dfm_mx0) + 50'b1;
  assign FpAdd_8U_23U_asn_34_mx1w1 = nl_FpAdd_8U_23U_asn_34_mx1w1[49:0];
  assign and_1009_nl = reg_alu_loop_op_15_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
      & (cfg_alu_algo_1_sva_st_204==2'b10);
  assign and_1011_nl = (~ reg_alu_loop_op_15_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse)
      & (cfg_alu_algo_1_sva_st_204==2'b10);
  assign FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_mx1 = MUX1HOT_v_50_3_2(FpAdd_8U_23U_int_mant_p1_15_sva,
      FpAdd_8U_23U_asn_34_mx1w1, FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm, {(and_1009_nl)
      , (and_1011_nl) , or_334_cse});
  assign FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_mx2 = MUX_v_50_2_2(FpAdd_8U_23U_asn_34_mx1w1,
      FpAdd_8U_23U_int_mant_p1_15_sva, reg_alu_loop_op_15_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse);
  assign nl_FpAdd_8U_23U_asn_mx1w1 = ({1'b1 , (~ FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_mx0) + 50'b1;
  assign FpAdd_8U_23U_asn_mx1w1 = nl_FpAdd_8U_23U_asn_mx1w1[49:0];
  assign and_1024_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & reg_alu_loop_op_16_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign and_1026_nl = (~ (cfg_alu_algo_1_sva_st_204[0])) & (~ reg_alu_loop_op_16_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse)
      & (cfg_alu_algo_1_sva_st_204[1]);
  assign FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_mx1 = MUX1HOT_v_50_3_2(FpAdd_8U_23U_int_mant_p1_sva,
      FpAdd_8U_23U_asn_mx1w1, FpAdd_8U_23U_int_mant_p1_lpi_1_dfm, {(and_1024_nl)
      , (and_1026_nl) , or_334_cse});
  assign FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_mx2 = MUX_v_50_2_2(FpAdd_8U_23U_asn_mx1w1,
      FpAdd_8U_23U_int_mant_p1_sva, reg_alu_loop_op_16_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse);
  assign alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0 = ~(alu_loop_op_4_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm_2
      & alu_loop_op_4_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm_2);
  assign alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0 = ~(alu_loop_op_6_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm_2
      & alu_loop_op_6_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm_2);
  assign alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0 = ~(alu_loop_op_13_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_itm_2
      & alu_loop_op_13_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_itm_2);
  assign alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0 = ~((~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_9_0_mx2!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_mx0w0!=4'b0000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0
      = ~((AluIn_data_sva_1[31]) ^ alu_nan_to_zero_op_sign_1_lpi_1_dfm_mx0w0);
  assign alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0 = ~((~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_9_0_mx2!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_mx0w0!=4'b0000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0
      = ~((AluIn_data_sva_1[63]) ^ alu_nan_to_zero_op_sign_2_lpi_1_dfm_mx0w0);
  assign alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0 = ~((~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_9_0_mx2!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_mx0w0!=4'b0000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0
      = ~((AluIn_data_sva_1[95]) ^ alu_nan_to_zero_op_sign_3_lpi_1_dfm_mx0w0);
  assign alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0
      = ~((AluIn_data_sva_1[127]) ^ alu_nan_to_zero_op_sign_4_lpi_1_dfm_mx0w0);
  assign alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0 = ~((~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_9_0_mx2!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_mx0w0!=4'b0000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign alu_loop_op_5_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0
      = ~((AluIn_data_sva_1[159]) ^ alu_nan_to_zero_op_sign_5_lpi_1_dfm_mx0w0);
  assign alu_loop_op_6_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0
      = ~((AluIn_data_sva_1[191]) ^ alu_nan_to_zero_op_sign_6_lpi_1_dfm_mx0w0);
  assign alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0 = ~((~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_9_0_mx2!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_mx0w0!=4'b0000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign alu_loop_op_7_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0
      = ~((AluIn_data_sva_1[223]) ^ alu_nan_to_zero_op_sign_7_lpi_1_dfm_mx0w0);
  assign alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0 = ~((~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_9_0_mx2!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_mx0w0!=4'b0000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign alu_loop_op_8_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0
      = ~((AluIn_data_sva_1[255]) ^ alu_nan_to_zero_op_sign_8_lpi_1_dfm_mx0w0);
  assign alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0 = ~((~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_9_0_mx2!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_mx0w0!=4'b0000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign alu_loop_op_9_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0
      = ~((AluIn_data_sva_1[287]) ^ alu_nan_to_zero_op_sign_9_lpi_1_dfm_mx0w0);
  assign alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0 = ~((~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_9_0_mx2!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_mx0w0!=4'b0000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign alu_loop_op_10_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0
      = ~((AluIn_data_sva_1[319]) ^ alu_nan_to_zero_op_sign_10_lpi_1_dfm_mx0w0);
  assign alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0 = ~((~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_9_0_mx2!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_mx0w0!=4'b0000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign alu_loop_op_11_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0
      = ~((AluIn_data_sva_1[351]) ^ alu_nan_to_zero_op_sign_11_lpi_1_dfm_mx0w0);
  assign alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0 = ~((~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_9_0_mx2!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_mx0w0!=4'b0000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign alu_loop_op_12_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0
      = ~((AluIn_data_sva_1[383]) ^ alu_nan_to_zero_op_sign_12_lpi_1_dfm_mx0w0);
  assign alu_loop_op_13_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0
      = ~((AluIn_data_sva_1[415]) ^ alu_nan_to_zero_op_sign_13_lpi_1_dfm_mx0w0);
  assign alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0 = ~((~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_9_0_mx2!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_mx0w0!=4'b0000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign alu_loop_op_14_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0
      = ~((AluIn_data_sva_1[447]) ^ alu_nan_to_zero_op_sign_14_lpi_1_dfm_mx0w0);
  assign alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0 = ~((~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_9_0_mx2!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_mx0w0!=4'b0000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign alu_loop_op_15_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0
      = ~((AluIn_data_sva_1[479]) ^ alu_nan_to_zero_op_sign_15_lpi_1_dfm_mx0w0);
  assign alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0 = ~((~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_12_10_mx0w0!=3'b000) |
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_9_0_mx2!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_mx0w0!=4'b0000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign alu_loop_op_16_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0
      = ~((AluIn_data_sva_1[511]) ^ alu_nan_to_zero_op_sign_lpi_1_dfm_mx0w0);
  assign alu_loop_op_4_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm_mx0w0
      = ~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_9_0_mx2!=10'b0000000000));
  assign alu_loop_op_4_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm_mx0w0 = ~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_mx0w0!=4'b0000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3_mx0w0!=4'b0000));
  assign alu_loop_op_6_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm_mx0w0
      = ~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_9_0_mx2!=10'b0000000000));
  assign alu_loop_op_6_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm_mx0w0 = ~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_mx0w0!=4'b0000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3_mx0w0!=4'b0000));
  assign alu_loop_op_13_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_itm_mx0w0 =
      ~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_9_0_mx2!=10'b0000000000));
  assign alu_loop_op_13_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_itm_mx0w0 = ~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_mx0w0!=4'b0000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3_mx0w0!=4'b0000));
  assign FpAlu_8U_23U_or_831_itm_mx0w0 = ((~ FpCmp_8U_23U_true_else_3_and_tmp) &
      FpAlu_8U_23U_and_66_m1c) | (FpCmp_8U_23U_false_else_3_or_tmp & FpAlu_8U_23U_and_68_m1c);
  assign FpAlu_8U_23U_or_752_itm_mx0w0 = (FpCmp_8U_23U_true_else_3_and_tmp & FpAlu_8U_23U_and_66_m1c)
      | FpAlu_8U_23U_and_67_cse | FpAlu_8U_23U_and_69_cse | ((~ FpCmp_8U_23U_false_else_3_or_tmp)
      & FpAlu_8U_23U_and_68_m1c);
  assign FpAlu_8U_23U_or_833_itm_mx0w0 = ((~ FpCmp_8U_23U_true_else_3_and_3_tmp)
      & FpAlu_8U_23U_and_80_m1c) | (FpCmp_8U_23U_false_else_3_or_3_tmp & FpAlu_8U_23U_and_82_m1c);
  assign FpAlu_8U_23U_or_755_itm_mx0w0 = (FpCmp_8U_23U_true_else_3_and_3_tmp & FpAlu_8U_23U_and_80_m1c)
      | FpAlu_8U_23U_and_81_cse | FpAlu_8U_23U_and_83_cse | ((~ FpCmp_8U_23U_false_else_3_or_3_tmp)
      & FpAlu_8U_23U_and_82_m1c);
  assign FpAlu_8U_23U_or_835_itm_mx0w0 = ((~ FpCmp_8U_23U_true_else_3_and_6_tmp)
      & FpAlu_8U_23U_and_94_m1c) | (FpCmp_8U_23U_false_else_3_or_6_tmp & FpAlu_8U_23U_and_96_m1c);
  assign FpAlu_8U_23U_or_758_itm_mx0w0 = (FpCmp_8U_23U_true_else_3_and_6_tmp & FpAlu_8U_23U_and_94_m1c)
      | FpAlu_8U_23U_and_95_cse | FpAlu_8U_23U_and_97_cse | ((~ FpCmp_8U_23U_false_else_3_or_6_tmp)
      & FpAlu_8U_23U_and_96_m1c);
  assign FpAlu_8U_23U_or_837_itm_mx0w0 = ((~ FpCmp_8U_23U_true_else_3_and_9_tmp)
      & FpAlu_8U_23U_and_108_m1c) | (FpCmp_8U_23U_false_else_3_or_9_tmp & FpAlu_8U_23U_and_110_m1c);
  assign FpAlu_8U_23U_or_761_itm_mx0w0 = (FpCmp_8U_23U_true_else_3_and_9_tmp & FpAlu_8U_23U_and_108_m1c)
      | FpAlu_8U_23U_and_109_cse | FpAlu_8U_23U_and_111_cse | ((~ FpCmp_8U_23U_false_else_3_or_9_tmp)
      & FpAlu_8U_23U_and_110_m1c);
  assign FpAlu_8U_23U_or_839_itm_mx0w0 = ((~ FpCmp_8U_23U_true_else_3_and_12_tmp)
      & FpAlu_8U_23U_and_122_m1c) | (FpCmp_8U_23U_false_else_3_or_12_tmp & FpAlu_8U_23U_and_124_m1c);
  assign FpAlu_8U_23U_or_764_itm_mx0w0 = (FpCmp_8U_23U_true_else_3_and_12_tmp & FpAlu_8U_23U_and_122_m1c)
      | FpAlu_8U_23U_and_123_cse | FpAlu_8U_23U_and_125_cse | ((~ FpCmp_8U_23U_false_else_3_or_12_tmp)
      & FpAlu_8U_23U_and_124_m1c);
  assign FpAlu_8U_23U_or_841_itm_mx0w0 = ((~ FpCmp_8U_23U_true_else_3_and_15_tmp)
      & FpAlu_8U_23U_and_136_m1c) | (FpCmp_8U_23U_false_else_3_or_15_tmp & FpAlu_8U_23U_and_138_m1c);
  assign FpAlu_8U_23U_or_767_itm_mx0w0 = (FpCmp_8U_23U_true_else_3_and_15_tmp & FpAlu_8U_23U_and_136_m1c)
      | FpAlu_8U_23U_and_137_cse | FpAlu_8U_23U_and_139_cse | ((~ FpCmp_8U_23U_false_else_3_or_15_tmp)
      & FpAlu_8U_23U_and_138_m1c);
  assign FpAlu_8U_23U_or_843_itm_mx0w0 = ((~ FpCmp_8U_23U_true_else_3_and_18_tmp)
      & FpAlu_8U_23U_and_150_m1c) | (FpCmp_8U_23U_false_else_3_or_18_tmp & FpAlu_8U_23U_and_152_m1c);
  assign FpAlu_8U_23U_or_770_itm_mx0w0 = (FpCmp_8U_23U_true_else_3_and_18_tmp & FpAlu_8U_23U_and_150_m1c)
      | FpAlu_8U_23U_and_151_cse | FpAlu_8U_23U_and_153_cse | ((~ FpCmp_8U_23U_false_else_3_or_18_tmp)
      & FpAlu_8U_23U_and_152_m1c);
  assign FpAlu_8U_23U_or_845_itm_mx0w0 = ((~ FpCmp_8U_23U_true_else_3_and_21_tmp)
      & FpAlu_8U_23U_and_164_m1c) | (FpCmp_8U_23U_false_else_3_or_21_tmp & FpAlu_8U_23U_and_166_m1c);
  assign FpAlu_8U_23U_or_773_itm_mx0w0 = (FpCmp_8U_23U_true_else_3_and_21_tmp & FpAlu_8U_23U_and_164_m1c)
      | FpAlu_8U_23U_and_165_cse | FpAlu_8U_23U_and_167_cse | ((~ FpCmp_8U_23U_false_else_3_or_21_tmp)
      & FpAlu_8U_23U_and_166_m1c);
  assign FpAlu_8U_23U_or_847_itm_mx0w0 = ((~ FpCmp_8U_23U_true_else_3_and_24_tmp)
      & FpAlu_8U_23U_and_178_m1c) | (FpCmp_8U_23U_false_else_3_or_24_tmp & FpAlu_8U_23U_and_180_m1c);
  assign FpAlu_8U_23U_or_776_itm_mx0w0 = (FpCmp_8U_23U_true_else_3_and_24_tmp & FpAlu_8U_23U_and_178_m1c)
      | FpAlu_8U_23U_and_179_cse | FpAlu_8U_23U_and_181_cse | ((~ FpCmp_8U_23U_false_else_3_or_24_tmp)
      & FpAlu_8U_23U_and_180_m1c);
  assign FpAlu_8U_23U_or_849_itm_mx0w0 = ((~ FpCmp_8U_23U_true_else_3_and_27_tmp)
      & FpAlu_8U_23U_and_192_m1c) | (FpCmp_8U_23U_false_else_3_or_27_tmp & FpAlu_8U_23U_and_194_m1c);
  assign FpAlu_8U_23U_or_779_itm_mx0w0 = (FpCmp_8U_23U_true_else_3_and_27_tmp & FpAlu_8U_23U_and_192_m1c)
      | FpAlu_8U_23U_and_193_cse | FpAlu_8U_23U_and_195_cse | ((~ FpCmp_8U_23U_false_else_3_or_27_tmp)
      & FpAlu_8U_23U_and_194_m1c);
  assign FpAlu_8U_23U_or_851_itm_mx0w0 = ((~ FpCmp_8U_23U_true_else_3_and_30_tmp)
      & FpAlu_8U_23U_and_206_m1c) | (FpCmp_8U_23U_false_else_3_or_30_tmp & FpAlu_8U_23U_and_208_m1c);
  assign FpAlu_8U_23U_or_782_itm_mx0w0 = (FpCmp_8U_23U_true_else_3_and_30_tmp & FpAlu_8U_23U_and_206_m1c)
      | FpAlu_8U_23U_and_207_cse | FpAlu_8U_23U_and_209_cse | ((~ FpCmp_8U_23U_false_else_3_or_30_tmp)
      & FpAlu_8U_23U_and_208_m1c);
  assign FpAlu_8U_23U_or_853_itm_mx0w0 = ((~ FpCmp_8U_23U_true_else_3_and_33_tmp)
      & FpAlu_8U_23U_and_220_m1c) | (FpCmp_8U_23U_false_else_3_or_33_tmp & FpAlu_8U_23U_and_222_m1c);
  assign FpAlu_8U_23U_or_785_itm_mx0w0 = (FpCmp_8U_23U_true_else_3_and_33_tmp & FpAlu_8U_23U_and_220_m1c)
      | FpAlu_8U_23U_and_221_cse | FpAlu_8U_23U_and_223_cse | ((~ FpCmp_8U_23U_false_else_3_or_33_tmp)
      & FpAlu_8U_23U_and_222_m1c);
  assign FpAlu_8U_23U_or_855_itm_mx0w0 = ((~ FpCmp_8U_23U_true_else_3_and_36_tmp)
      & FpAlu_8U_23U_and_234_m1c) | (FpCmp_8U_23U_false_else_3_or_36_tmp & FpAlu_8U_23U_and_236_m1c);
  assign FpAlu_8U_23U_or_788_itm_mx0w0 = (FpCmp_8U_23U_true_else_3_and_36_tmp & FpAlu_8U_23U_and_234_m1c)
      | FpAlu_8U_23U_and_235_cse | FpAlu_8U_23U_and_237_cse | ((~ FpCmp_8U_23U_false_else_3_or_36_tmp)
      & FpAlu_8U_23U_and_236_m1c);
  assign FpAlu_8U_23U_or_857_itm_mx0w0 = ((~ FpCmp_8U_23U_true_else_3_and_39_tmp)
      & FpAlu_8U_23U_and_248_m1c) | (FpCmp_8U_23U_false_else_3_or_39_tmp & FpAlu_8U_23U_and_250_m1c);
  assign FpAlu_8U_23U_or_791_itm_mx0w0 = (FpCmp_8U_23U_true_else_3_and_39_tmp & FpAlu_8U_23U_and_248_m1c)
      | FpAlu_8U_23U_and_249_cse | FpAlu_8U_23U_and_251_cse | ((~ FpCmp_8U_23U_false_else_3_or_39_tmp)
      & FpAlu_8U_23U_and_250_m1c);
  assign FpAlu_8U_23U_or_859_itm_mx0w0 = ((~ FpCmp_8U_23U_true_else_3_and_42_tmp)
      & FpAlu_8U_23U_and_262_m1c) | (FpCmp_8U_23U_false_else_3_or_42_tmp & FpAlu_8U_23U_and_264_m1c);
  assign FpAlu_8U_23U_or_794_itm_mx0w0 = (FpCmp_8U_23U_true_else_3_and_42_tmp & FpAlu_8U_23U_and_262_m1c)
      | FpAlu_8U_23U_and_263_cse | FpAlu_8U_23U_and_265_cse | ((~ FpCmp_8U_23U_false_else_3_or_42_tmp)
      & FpAlu_8U_23U_and_264_m1c);
  assign FpAlu_8U_23U_or_861_itm_mx0w0 = ((~ FpCmp_8U_23U_true_else_3_and_45_tmp)
      & FpAlu_8U_23U_and_276_m1c) | (FpCmp_8U_23U_false_else_3_or_45_tmp & FpAlu_8U_23U_and_278_m1c);
  assign FpAlu_8U_23U_or_797_itm_mx0w0 = (FpCmp_8U_23U_true_else_3_and_45_tmp & FpAlu_8U_23U_and_276_m1c)
      | FpAlu_8U_23U_and_277_cse | FpAlu_8U_23U_and_279_cse | ((~ FpCmp_8U_23U_false_else_3_or_45_tmp)
      & FpAlu_8U_23U_and_278_m1c);
  assign FpAlu_8U_23U_or_800_nl = (FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w4
      & (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_7) & (~ IsNaN_8U_23U_land_1_lpi_1_dfm_8)
      & FpAlu_8U_23U_nor_dfs_mx0w0) | (IsNaN_8U_23U_land_1_lpi_1_dfm_8 & FpAlu_8U_23U_nor_dfs_mx0w0)
      | (FpCmp_8U_23U_true_is_a_greater_1_lpi_1_dfm_2_mx0 & (~ IsNaN_8U_23U_3_land_1_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_66_m1c) | FpAlu_8U_23U_and_67_cse | FpAlu_8U_23U_and_69_cse
      | ((~ FpCmp_8U_23U_false_is_a_greater_1_lpi_1_dfm_2_mx0) & (~ IsNaN_8U_23U_3_land_1_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_68_m1c);
  assign FpAlu_8U_23U_FpAlu_8U_23U_mux_15_nl = MUX_s_1_2_2(alu_nan_to_zero_op_sign_1_lpi_1_dfm_4,
      (AluIn_data_sva_501[31]), FpAlu_8U_23U_or_800_nl);
  assign FpAlu_8U_23U_and_itm_mx0w0 = (FpAlu_8U_23U_FpAlu_8U_23U_mux_15_nl) & (~
      and_3689_cse);
  assign FpAlu_8U_23U_or_802_nl = (FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w4
      & (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_7) & (~ IsNaN_8U_23U_land_2_lpi_1_dfm_8)
      & FpAlu_8U_23U_nor_dfs_mx0w0) | (IsNaN_8U_23U_land_2_lpi_1_dfm_8 & FpAlu_8U_23U_nor_dfs_mx0w0)
      | (FpCmp_8U_23U_true_is_a_greater_2_lpi_1_dfm_2_mx0 & (~ IsNaN_8U_23U_3_land_2_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_80_m1c) | FpAlu_8U_23U_and_81_cse | FpAlu_8U_23U_and_83_cse
      | ((~ FpCmp_8U_23U_false_is_a_greater_2_lpi_1_dfm_2_mx0) & (~ IsNaN_8U_23U_3_land_2_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_82_m1c);
  assign FpAlu_8U_23U_FpAlu_8U_23U_mux_14_nl = MUX_s_1_2_2(alu_nan_to_zero_op_sign_2_lpi_1_dfm_4,
      (AluIn_data_sva_501[63]), FpAlu_8U_23U_or_802_nl);
  assign FpAlu_8U_23U_and_4_itm_mx0w0 = (FpAlu_8U_23U_FpAlu_8U_23U_mux_14_nl) & (~
      and_3689_cse);
  assign FpAlu_8U_23U_or_804_nl = (FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w4
      & (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_7) & (~ IsNaN_8U_23U_land_3_lpi_1_dfm_8)
      & FpAlu_8U_23U_nor_dfs_mx0w0) | (IsNaN_8U_23U_land_3_lpi_1_dfm_8 & FpAlu_8U_23U_nor_dfs_mx0w0)
      | (FpCmp_8U_23U_true_is_a_greater_3_lpi_1_dfm_2_mx0 & (~ IsNaN_8U_23U_3_land_3_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_94_m1c) | FpAlu_8U_23U_and_95_cse | FpAlu_8U_23U_and_97_cse
      | ((~ FpCmp_8U_23U_false_is_a_greater_3_lpi_1_dfm_2_mx0) & (~ IsNaN_8U_23U_3_land_3_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_96_m1c);
  assign FpAlu_8U_23U_FpAlu_8U_23U_mux_13_nl = MUX_s_1_2_2(alu_nan_to_zero_op_sign_3_lpi_1_dfm_4,
      (AluIn_data_sva_501[95]), FpAlu_8U_23U_or_804_nl);
  assign FpAlu_8U_23U_and_8_itm_mx0w0 = (FpAlu_8U_23U_FpAlu_8U_23U_mux_13_nl) & (~
      and_3689_cse);
  assign FpAlu_8U_23U_or_806_nl = (FpAdd_8U_23U_is_a_greater_lor_4_lpi_1_dfm_1_mx0w4
      & (~ IsNaN_8U_23U_1_land_4_lpi_1_dfm_7) & (~ IsNaN_8U_23U_land_4_lpi_1_dfm_8)
      & FpAlu_8U_23U_nor_dfs_mx0w0) | (IsNaN_8U_23U_land_4_lpi_1_dfm_8 & FpAlu_8U_23U_nor_dfs_mx0w0)
      | (FpCmp_8U_23U_true_is_a_greater_4_lpi_1_dfm_2_mx0 & (~ IsNaN_8U_23U_3_land_4_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_108_m1c) | FpAlu_8U_23U_and_109_cse | FpAlu_8U_23U_and_111_cse
      | ((~ FpCmp_8U_23U_false_is_a_greater_4_lpi_1_dfm_2_mx0) & (~ IsNaN_8U_23U_3_land_4_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_110_m1c);
  assign FpAlu_8U_23U_FpAlu_8U_23U_mux_12_nl = MUX_s_1_2_2(alu_nan_to_zero_op_sign_4_lpi_1_dfm_4,
      (AluIn_data_sva_501[127]), FpAlu_8U_23U_or_806_nl);
  assign FpAlu_8U_23U_and_12_itm_mx0w0 = (FpAlu_8U_23U_FpAlu_8U_23U_mux_12_nl) &
      (~ and_3689_cse);
  assign FpAlu_8U_23U_or_808_nl = (FpAdd_8U_23U_is_a_greater_lor_5_lpi_1_dfm_1_mx0w4
      & (~ IsNaN_8U_23U_1_land_5_lpi_1_dfm_7) & (~ IsNaN_8U_23U_land_5_lpi_1_dfm_8)
      & FpAlu_8U_23U_nor_dfs_mx0w0) | (IsNaN_8U_23U_land_5_lpi_1_dfm_8 & FpAlu_8U_23U_nor_dfs_mx0w0)
      | (FpCmp_8U_23U_true_is_a_greater_5_lpi_1_dfm_2_mx0 & (~ IsNaN_8U_23U_3_land_5_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_122_m1c) | FpAlu_8U_23U_and_123_cse | FpAlu_8U_23U_and_125_cse
      | ((~ FpCmp_8U_23U_false_is_a_greater_5_lpi_1_dfm_2_mx0) & (~ IsNaN_8U_23U_3_land_5_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_124_m1c);
  assign FpAlu_8U_23U_FpAlu_8U_23U_mux_11_nl = MUX_s_1_2_2(alu_nan_to_zero_op_sign_5_lpi_1_dfm_4,
      (AluIn_data_sva_501[159]), FpAlu_8U_23U_or_808_nl);
  assign FpAlu_8U_23U_and_16_itm_mx0w0 = (FpAlu_8U_23U_FpAlu_8U_23U_mux_11_nl) &
      (~ and_3689_cse);
  assign FpAlu_8U_23U_or_810_nl = (FpAdd_8U_23U_is_a_greater_lor_6_lpi_1_dfm_1_mx0w4
      & (~ IsNaN_8U_23U_1_land_6_lpi_1_dfm_7) & (~ IsNaN_8U_23U_land_6_lpi_1_dfm_8)
      & FpAlu_8U_23U_nor_dfs_mx0w0) | (IsNaN_8U_23U_land_6_lpi_1_dfm_8 & FpAlu_8U_23U_nor_dfs_mx0w0)
      | (FpCmp_8U_23U_true_is_a_greater_6_lpi_1_dfm_2_mx0 & (~ IsNaN_8U_23U_3_land_6_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_136_m1c) | FpAlu_8U_23U_and_137_cse | FpAlu_8U_23U_and_139_cse
      | ((~ FpCmp_8U_23U_false_is_a_greater_6_lpi_1_dfm_2_mx0) & (~ IsNaN_8U_23U_3_land_6_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_138_m1c);
  assign FpAlu_8U_23U_FpAlu_8U_23U_mux_10_nl = MUX_s_1_2_2(alu_nan_to_zero_op_sign_6_lpi_1_dfm_4,
      (AluIn_data_sva_501[191]), FpAlu_8U_23U_or_810_nl);
  assign FpAlu_8U_23U_and_20_itm_mx0w0 = (FpAlu_8U_23U_FpAlu_8U_23U_mux_10_nl) &
      (~ and_3689_cse);
  assign FpAlu_8U_23U_or_812_nl = (FpAdd_8U_23U_is_a_greater_lor_7_lpi_1_dfm_1_mx0w4
      & (~ IsNaN_8U_23U_1_land_7_lpi_1_dfm_7) & (~ IsNaN_8U_23U_land_7_lpi_1_dfm_8)
      & FpAlu_8U_23U_nor_dfs_mx0w0) | (IsNaN_8U_23U_land_7_lpi_1_dfm_8 & FpAlu_8U_23U_nor_dfs_mx0w0)
      | (FpCmp_8U_23U_true_is_a_greater_7_lpi_1_dfm_2_mx0 & (~ IsNaN_8U_23U_3_land_7_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_150_m1c) | FpAlu_8U_23U_and_151_cse | FpAlu_8U_23U_and_153_cse
      | ((~ FpCmp_8U_23U_false_is_a_greater_7_lpi_1_dfm_2_mx0) & (~ IsNaN_8U_23U_3_land_7_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_152_m1c);
  assign FpAlu_8U_23U_FpAlu_8U_23U_mux_9_nl = MUX_s_1_2_2(alu_nan_to_zero_op_sign_7_lpi_1_dfm_4,
      (AluIn_data_sva_501[223]), FpAlu_8U_23U_or_812_nl);
  assign FpAlu_8U_23U_and_24_itm_mx0w0 = (FpAlu_8U_23U_FpAlu_8U_23U_mux_9_nl) & (~
      and_3689_cse);
  assign FpAlu_8U_23U_or_814_nl = (FpAdd_8U_23U_is_a_greater_lor_8_lpi_1_dfm_1_mx0w4
      & (~ IsNaN_8U_23U_1_land_8_lpi_1_dfm_7) & (~ IsNaN_8U_23U_land_8_lpi_1_dfm_8)
      & FpAlu_8U_23U_nor_dfs_mx0w0) | (IsNaN_8U_23U_land_8_lpi_1_dfm_8 & FpAlu_8U_23U_nor_dfs_mx0w0)
      | (FpCmp_8U_23U_true_is_a_greater_8_lpi_1_dfm_2_mx0 & (~ IsNaN_8U_23U_3_land_8_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_164_m1c) | FpAlu_8U_23U_and_165_cse | FpAlu_8U_23U_and_167_cse
      | ((~ FpCmp_8U_23U_false_is_a_greater_8_lpi_1_dfm_2_mx0) & (~ IsNaN_8U_23U_3_land_8_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_166_m1c);
  assign FpAlu_8U_23U_FpAlu_8U_23U_mux_8_nl = MUX_s_1_2_2(alu_nan_to_zero_op_sign_8_lpi_1_dfm_3,
      (AluIn_data_sva_501[255]), FpAlu_8U_23U_or_814_nl);
  assign FpAlu_8U_23U_and_28_itm_mx0w0 = (FpAlu_8U_23U_FpAlu_8U_23U_mux_8_nl) & (~
      and_3689_cse);
  assign FpAlu_8U_23U_or_816_nl = (FpAdd_8U_23U_is_a_greater_lor_9_lpi_1_dfm_1_mx0w4
      & (~ IsNaN_8U_23U_1_land_9_lpi_1_dfm_7) & (~ IsNaN_8U_23U_land_9_lpi_1_dfm_8)
      & FpAlu_8U_23U_nor_dfs_mx0w0) | (IsNaN_8U_23U_land_9_lpi_1_dfm_8 & FpAlu_8U_23U_nor_dfs_mx0w0)
      | (FpCmp_8U_23U_true_is_a_greater_9_lpi_1_dfm_2_mx0 & (~ IsNaN_8U_23U_3_land_9_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_178_m1c) | FpAlu_8U_23U_and_179_cse | FpAlu_8U_23U_and_181_cse
      | ((~ FpCmp_8U_23U_false_is_a_greater_9_lpi_1_dfm_2_mx0) & (~ IsNaN_8U_23U_3_land_9_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_180_m1c);
  assign FpAlu_8U_23U_FpAlu_8U_23U_mux_7_nl = MUX_s_1_2_2(alu_nan_to_zero_op_sign_9_lpi_1_dfm_3,
      (AluIn_data_sva_501[287]), FpAlu_8U_23U_or_816_nl);
  assign FpAlu_8U_23U_and_32_itm_mx0w0 = (FpAlu_8U_23U_FpAlu_8U_23U_mux_7_nl) & (~
      and_3689_cse);
  assign FpAlu_8U_23U_or_818_nl = (FpAdd_8U_23U_is_a_greater_lor_10_lpi_1_dfm_1_mx0w4
      & (~ IsNaN_8U_23U_1_land_10_lpi_1_dfm_7) & (~ IsNaN_8U_23U_land_10_lpi_1_dfm_8)
      & FpAlu_8U_23U_nor_dfs_mx0w0) | (IsNaN_8U_23U_land_10_lpi_1_dfm_8 & FpAlu_8U_23U_nor_dfs_mx0w0)
      | (FpCmp_8U_23U_true_is_a_greater_10_lpi_1_dfm_2_mx0 & (~ IsNaN_8U_23U_3_land_10_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_192_m1c) | FpAlu_8U_23U_and_193_cse | FpAlu_8U_23U_and_195_cse
      | ((~ FpCmp_8U_23U_false_is_a_greater_10_lpi_1_dfm_2_mx0) & (~ IsNaN_8U_23U_3_land_10_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_194_m1c);
  assign FpAlu_8U_23U_FpAlu_8U_23U_mux_6_nl = MUX_s_1_2_2(alu_nan_to_zero_op_sign_10_lpi_1_dfm_3,
      (AluIn_data_sva_501[319]), FpAlu_8U_23U_or_818_nl);
  assign FpAlu_8U_23U_and_36_itm_mx0w0 = (FpAlu_8U_23U_FpAlu_8U_23U_mux_6_nl) & (~
      and_3689_cse);
  assign FpAlu_8U_23U_or_820_nl = (FpAdd_8U_23U_is_a_greater_lor_11_lpi_1_dfm_1_mx0w4
      & (~ IsNaN_8U_23U_1_land_11_lpi_1_dfm_7) & (~ IsNaN_8U_23U_land_11_lpi_1_dfm_8)
      & FpAlu_8U_23U_nor_dfs_mx0w0) | (IsNaN_8U_23U_land_11_lpi_1_dfm_8 & FpAlu_8U_23U_nor_dfs_mx0w0)
      | (FpCmp_8U_23U_true_is_a_greater_11_lpi_1_dfm_2_mx0 & (~ IsNaN_8U_23U_3_land_11_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_206_m1c) | FpAlu_8U_23U_and_207_cse | FpAlu_8U_23U_and_209_cse
      | ((~ FpCmp_8U_23U_false_is_a_greater_11_lpi_1_dfm_2_mx0) & (~ IsNaN_8U_23U_3_land_11_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_208_m1c);
  assign FpAlu_8U_23U_FpAlu_8U_23U_mux_5_nl = MUX_s_1_2_2(alu_nan_to_zero_op_sign_11_lpi_1_dfm_3,
      (AluIn_data_sva_501[351]), FpAlu_8U_23U_or_820_nl);
  assign FpAlu_8U_23U_and_40_itm_mx0w0 = (FpAlu_8U_23U_FpAlu_8U_23U_mux_5_nl) & (~
      and_3689_cse);
  assign FpAlu_8U_23U_or_822_nl = (FpAdd_8U_23U_is_a_greater_lor_12_lpi_1_dfm_1_mx0w4
      & (~ IsNaN_8U_23U_1_land_12_lpi_1_dfm_7) & (~ IsNaN_8U_23U_land_12_lpi_1_dfm_8)
      & FpAlu_8U_23U_nor_dfs_mx0w0) | (IsNaN_8U_23U_land_12_lpi_1_dfm_8 & FpAlu_8U_23U_nor_dfs_mx0w0)
      | (FpCmp_8U_23U_true_is_a_greater_12_lpi_1_dfm_2_mx0 & (~ IsNaN_8U_23U_3_land_12_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_220_m1c) | FpAlu_8U_23U_and_221_cse | FpAlu_8U_23U_and_223_cse
      | ((~ FpCmp_8U_23U_false_is_a_greater_12_lpi_1_dfm_2_mx0) & (~ IsNaN_8U_23U_3_land_12_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_222_m1c);
  assign FpAlu_8U_23U_FpAlu_8U_23U_mux_4_nl = MUX_s_1_2_2(alu_nan_to_zero_op_sign_12_lpi_1_dfm_3,
      (AluIn_data_sva_501[383]), FpAlu_8U_23U_or_822_nl);
  assign FpAlu_8U_23U_and_44_itm_mx0w0 = (FpAlu_8U_23U_FpAlu_8U_23U_mux_4_nl) & (~
      and_3689_cse);
  assign FpAlu_8U_23U_or_824_nl = (FpAdd_8U_23U_is_a_greater_lor_13_lpi_1_dfm_1_mx0w4
      & (~ IsNaN_8U_23U_1_land_13_lpi_1_dfm_7) & (~ IsNaN_8U_23U_land_13_lpi_1_dfm_8)
      & FpAlu_8U_23U_nor_dfs_mx0w0) | (IsNaN_8U_23U_land_13_lpi_1_dfm_8 & FpAlu_8U_23U_nor_dfs_mx0w0)
      | (FpCmp_8U_23U_true_is_a_greater_13_lpi_1_dfm_2_mx0 & (~ IsNaN_8U_23U_3_land_13_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_234_m1c) | FpAlu_8U_23U_and_235_cse | FpAlu_8U_23U_and_237_cse
      | ((~ FpCmp_8U_23U_false_is_a_greater_13_lpi_1_dfm_2_mx0) & (~ IsNaN_8U_23U_3_land_13_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_236_m1c);
  assign FpAlu_8U_23U_FpAlu_8U_23U_mux_3_nl = MUX_s_1_2_2(alu_nan_to_zero_op_sign_13_lpi_1_dfm_3,
      (AluIn_data_sva_501[415]), FpAlu_8U_23U_or_824_nl);
  assign FpAlu_8U_23U_and_48_itm_mx0w0 = (FpAlu_8U_23U_FpAlu_8U_23U_mux_3_nl) & (~
      and_3689_cse);
  assign FpAlu_8U_23U_or_826_nl = (FpAdd_8U_23U_is_a_greater_lor_14_lpi_1_dfm_1_mx0w4
      & (~ IsNaN_8U_23U_1_land_14_lpi_1_dfm_7) & (~ IsNaN_8U_23U_land_14_lpi_1_dfm_8)
      & FpAlu_8U_23U_nor_dfs_mx0w0) | (IsNaN_8U_23U_land_14_lpi_1_dfm_8 & FpAlu_8U_23U_nor_dfs_mx0w0)
      | (FpCmp_8U_23U_true_is_a_greater_14_lpi_1_dfm_2_mx0 & (~ IsNaN_8U_23U_3_land_14_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_248_m1c) | FpAlu_8U_23U_and_249_cse | FpAlu_8U_23U_and_251_cse
      | ((~ FpCmp_8U_23U_false_is_a_greater_14_lpi_1_dfm_2_mx0) & (~ IsNaN_8U_23U_3_land_14_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_250_m1c);
  assign FpAlu_8U_23U_FpAlu_8U_23U_mux_2_nl = MUX_s_1_2_2(alu_nan_to_zero_op_sign_14_lpi_1_dfm_3,
      (AluIn_data_sva_501[447]), FpAlu_8U_23U_or_826_nl);
  assign FpAlu_8U_23U_and_52_itm_mx0w0 = (FpAlu_8U_23U_FpAlu_8U_23U_mux_2_nl) & (~
      and_3689_cse);
  assign FpAlu_8U_23U_or_828_nl = (FpAdd_8U_23U_is_a_greater_lor_15_lpi_1_dfm_1_mx0w4
      & (~ IsNaN_8U_23U_1_land_15_lpi_1_dfm_7) & (~ IsNaN_8U_23U_land_15_lpi_1_dfm_8)
      & FpAlu_8U_23U_nor_dfs_mx0w0) | (IsNaN_8U_23U_land_15_lpi_1_dfm_8 & FpAlu_8U_23U_nor_dfs_mx0w0)
      | (FpCmp_8U_23U_true_is_a_greater_15_lpi_1_dfm_2_mx0 & (~ IsNaN_8U_23U_3_land_15_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_262_m1c) | FpAlu_8U_23U_and_263_cse | FpAlu_8U_23U_and_265_cse
      | ((~ FpCmp_8U_23U_false_is_a_greater_15_lpi_1_dfm_2_mx0) & (~ IsNaN_8U_23U_3_land_15_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_264_m1c);
  assign FpAlu_8U_23U_FpAlu_8U_23U_mux_1_nl = MUX_s_1_2_2(alu_nan_to_zero_op_sign_15_lpi_1_dfm_3,
      (AluIn_data_sva_501[479]), FpAlu_8U_23U_or_828_nl);
  assign FpAlu_8U_23U_and_56_itm_mx0w0 = (FpAlu_8U_23U_FpAlu_8U_23U_mux_1_nl) & (~
      and_3689_cse);
  assign FpAlu_8U_23U_or_830_nl = (FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w4
      & (~ IsNaN_8U_23U_1_land_lpi_1_dfm_7) & (~ IsNaN_8U_23U_land_lpi_1_dfm_8) &
      FpAlu_8U_23U_nor_dfs_mx0w0) | (IsNaN_8U_23U_land_lpi_1_dfm_8 & FpAlu_8U_23U_nor_dfs_mx0w0)
      | (FpCmp_8U_23U_true_is_a_greater_lpi_1_dfm_2_mx0 & (~ IsNaN_8U_23U_3_land_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_276_m1c) | FpAlu_8U_23U_and_277_cse | FpAlu_8U_23U_and_279_cse
      | ((~ FpCmp_8U_23U_false_is_a_greater_lpi_1_dfm_2_mx0) & (~ IsNaN_8U_23U_3_land_lpi_1_dfm_6)
      & FpAlu_8U_23U_and_278_m1c);
  assign FpAlu_8U_23U_FpAlu_8U_23U_mux_nl = MUX_s_1_2_2(alu_nan_to_zero_op_sign_lpi_1_dfm_3,
      (AluIn_data_sva_501[511]), FpAlu_8U_23U_or_830_nl);
  assign FpAlu_8U_23U_and_60_itm_mx0w0 = (FpAlu_8U_23U_FpAlu_8U_23U_mux_nl) & (~
      and_3689_cse);
  assign FpAlu_8U_23U_equal_tmp_mx0w0 = ~((cfg_alu_algo_1_sva_5!=2'b00));
  assign FpAlu_8U_23U_equal_tmp_2_mx0w0 = (cfg_alu_algo_1_sva_5==2'b01);
  assign FpAlu_8U_23U_nor_dfs_mx0w0 = ~(FpAlu_8U_23U_equal_tmp_mx0w0 | and_3689_cse
      | FpAlu_8U_23U_equal_tmp_2_mx0w0);
  assign FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_mx0w0 = (~ FpCmp_8U_23U_false_is_abs_a_greater_1_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_1_lpi_1_dfm_4;
  assign FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_mx0w1 = FpCmp_8U_23U_false_is_abs_a_greater_1_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_1_lpi_1_dfm_4;
  assign FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_mx0w2 = (~ FpCmp_8U_23U_true_is_abs_a_greater_1_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_1_lpi_1_dfm_4;
  assign FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_mx0w3 = FpCmp_8U_23U_true_is_abs_a_greater_1_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_1_lpi_1_dfm_4;
  assign FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w4 = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_itm_23_1)
      & alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2) | alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_1_mx0w0 = (~ FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_2_lpi_1_dfm_4;
  assign FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_1_mx0w1 = FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_2_lpi_1_dfm_4;
  assign FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_1_mx0w2 = (~ FpCmp_8U_23U_true_is_abs_a_greater_2_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_2_lpi_1_dfm_4;
  assign FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_1_mx0w3 = FpCmp_8U_23U_true_is_abs_a_greater_2_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_2_lpi_1_dfm_4;
  assign FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w4 = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_itm_23_1)
      & alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2) | alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_2_mx0w0 = (~ FpCmp_8U_23U_false_is_abs_a_greater_3_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_3_lpi_1_dfm_4;
  assign FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_2_mx0w1 = FpCmp_8U_23U_false_is_abs_a_greater_3_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_3_lpi_1_dfm_4;
  assign FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_2_mx0w2 = (~ FpCmp_8U_23U_true_is_abs_a_greater_3_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_3_lpi_1_dfm_4;
  assign FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_2_mx0w3 = FpCmp_8U_23U_true_is_abs_a_greater_3_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_3_lpi_1_dfm_4;
  assign FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w4 = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_itm_23_1)
      & alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2) | alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_3_mx0w0 = (~ FpCmp_8U_23U_false_is_abs_a_greater_4_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_4_lpi_1_dfm_4;
  assign FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_3_mx0w1 = FpCmp_8U_23U_false_is_abs_a_greater_4_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_4_lpi_1_dfm_4;
  assign FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_3_mx0w2 = (~ FpCmp_8U_23U_true_is_abs_a_greater_4_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_4_lpi_1_dfm_4;
  assign FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_3_mx0w3 = FpCmp_8U_23U_true_is_abs_a_greater_4_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_4_lpi_1_dfm_4;
  assign FpAdd_8U_23U_is_a_greater_lor_4_lpi_1_dfm_1_mx0w4 = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_itm_23_1)
      & alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2) | alu_loop_op_4_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_4_mx0w0 = (~ FpCmp_8U_23U_false_is_abs_a_greater_5_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_5_lpi_1_dfm_4;
  assign FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_4_mx0w1 = FpCmp_8U_23U_false_is_abs_a_greater_5_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_5_lpi_1_dfm_4;
  assign FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_4_mx0w2 = (~ FpCmp_8U_23U_true_is_abs_a_greater_5_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_5_lpi_1_dfm_4;
  assign FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_4_mx0w3 = FpCmp_8U_23U_true_is_abs_a_greater_5_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_5_lpi_1_dfm_4;
  assign FpAdd_8U_23U_is_a_greater_lor_5_lpi_1_dfm_1_mx0w4 = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_itm_23_1)
      & alu_loop_op_5_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2) | alu_loop_op_5_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_5_mx0w0 = (~ FpCmp_8U_23U_false_is_abs_a_greater_6_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_6_lpi_1_dfm_4;
  assign FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_5_mx0w1 = FpCmp_8U_23U_false_is_abs_a_greater_6_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_6_lpi_1_dfm_4;
  assign FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_5_mx0w2 = (~ FpCmp_8U_23U_true_is_abs_a_greater_6_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_6_lpi_1_dfm_4;
  assign FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_5_mx0w3 = FpCmp_8U_23U_true_is_abs_a_greater_6_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_6_lpi_1_dfm_4;
  assign FpAdd_8U_23U_is_a_greater_lor_6_lpi_1_dfm_1_mx0w4 = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_5_itm_23_1)
      & alu_loop_op_6_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2) | alu_loop_op_6_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_6_mx0w0 = (~ FpCmp_8U_23U_false_is_abs_a_greater_7_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_7_lpi_1_dfm_4;
  assign FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_6_mx0w1 = FpCmp_8U_23U_false_is_abs_a_greater_7_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_7_lpi_1_dfm_4;
  assign FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_6_mx0w2 = (~ FpCmp_8U_23U_true_is_abs_a_greater_7_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_7_lpi_1_dfm_4;
  assign FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_6_mx0w3 = FpCmp_8U_23U_true_is_abs_a_greater_7_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_7_lpi_1_dfm_4;
  assign FpAdd_8U_23U_is_a_greater_lor_7_lpi_1_dfm_1_mx0w4 = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_itm_23_1)
      & alu_loop_op_7_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2) | alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_7_mx0w0 = (~ FpCmp_8U_23U_false_is_abs_a_greater_8_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_8_lpi_1_dfm_3;
  assign FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_7_mx0w1 = FpCmp_8U_23U_false_is_abs_a_greater_8_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_8_lpi_1_dfm_3;
  assign FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_7_mx0w2 = (~ FpCmp_8U_23U_true_is_abs_a_greater_8_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_8_lpi_1_dfm_3;
  assign FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_7_mx0w3 = FpCmp_8U_23U_true_is_abs_a_greater_8_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_8_lpi_1_dfm_3;
  assign FpAdd_8U_23U_is_a_greater_lor_8_lpi_1_dfm_1_mx0w4 = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_7_itm_23_1)
      & alu_loop_op_8_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2) | alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_8_mx0w0 = (~ FpCmp_8U_23U_false_is_abs_a_greater_9_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_9_lpi_1_dfm_3;
  assign FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_8_mx0w1 = FpCmp_8U_23U_false_is_abs_a_greater_9_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_9_lpi_1_dfm_3;
  assign FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_8_mx0w2 = (~ FpCmp_8U_23U_true_is_abs_a_greater_9_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_9_lpi_1_dfm_3;
  assign FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_8_mx0w3 = FpCmp_8U_23U_true_is_abs_a_greater_9_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_9_lpi_1_dfm_3;
  assign FpAdd_8U_23U_is_a_greater_lor_9_lpi_1_dfm_1_mx0w4 = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_itm_23_1)
      & alu_loop_op_9_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2) | alu_loop_op_9_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_9_mx0w0 = (~ FpCmp_8U_23U_false_is_abs_a_greater_10_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_10_lpi_1_dfm_3;
  assign FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_9_mx0w1 = FpCmp_8U_23U_false_is_abs_a_greater_10_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_10_lpi_1_dfm_3;
  assign FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_9_mx0w2 = (~ FpCmp_8U_23U_true_is_abs_a_greater_10_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_10_lpi_1_dfm_3;
  assign FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_9_mx0w3 = FpCmp_8U_23U_true_is_abs_a_greater_10_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_10_lpi_1_dfm_3;
  assign FpAdd_8U_23U_is_a_greater_lor_10_lpi_1_dfm_1_mx0w4 = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_9_itm_23_1)
      & alu_loop_op_10_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2) | alu_loop_op_10_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_10_mx0w0 = (~ FpCmp_8U_23U_false_is_abs_a_greater_11_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_11_lpi_1_dfm_3;
  assign FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_10_mx0w1 = FpCmp_8U_23U_false_is_abs_a_greater_11_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_11_lpi_1_dfm_3;
  assign FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_10_mx0w2 = (~ FpCmp_8U_23U_true_is_abs_a_greater_11_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_11_lpi_1_dfm_3;
  assign FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_10_mx0w3 = FpCmp_8U_23U_true_is_abs_a_greater_11_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_11_lpi_1_dfm_3;
  assign FpAdd_8U_23U_is_a_greater_lor_11_lpi_1_dfm_1_mx0w4 = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_itm_23_1)
      & alu_loop_op_11_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2) | alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_11_mx0w0 = (~ FpCmp_8U_23U_false_is_abs_a_greater_12_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_12_lpi_1_dfm_3;
  assign FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_11_mx0w1 = FpCmp_8U_23U_false_is_abs_a_greater_12_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_12_lpi_1_dfm_3;
  assign FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_11_mx0w2 = (~ FpCmp_8U_23U_true_is_abs_a_greater_12_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_12_lpi_1_dfm_3;
  assign FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_11_mx0w3 = FpCmp_8U_23U_true_is_abs_a_greater_12_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_12_lpi_1_dfm_3;
  assign FpAdd_8U_23U_is_a_greater_lor_12_lpi_1_dfm_1_mx0w4 = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_11_itm_23_1)
      & alu_loop_op_12_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2) | alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_12_mx0w0 = (~ FpCmp_8U_23U_false_is_abs_a_greater_13_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_13_lpi_1_dfm_3;
  assign FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_12_mx0w1 = FpCmp_8U_23U_false_is_abs_a_greater_13_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_13_lpi_1_dfm_3;
  assign FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_12_mx0w2 = (~ FpCmp_8U_23U_true_is_abs_a_greater_13_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_13_lpi_1_dfm_3;
  assign FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_12_mx0w3 = FpCmp_8U_23U_true_is_abs_a_greater_13_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_13_lpi_1_dfm_3;
  assign FpAdd_8U_23U_is_a_greater_lor_13_lpi_1_dfm_1_mx0w4 = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_12_itm_23_1)
      & alu_loop_op_13_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2) | alu_loop_op_13_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_13_mx0w0 = (~ FpCmp_8U_23U_false_is_abs_a_greater_14_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_14_lpi_1_dfm_3;
  assign FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_13_mx0w1 = FpCmp_8U_23U_false_is_abs_a_greater_14_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_14_lpi_1_dfm_3;
  assign FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_13_mx0w2 = (~ FpCmp_8U_23U_true_is_abs_a_greater_14_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_14_lpi_1_dfm_3;
  assign FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_13_mx0w3 = FpCmp_8U_23U_true_is_abs_a_greater_14_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_14_lpi_1_dfm_3;
  assign FpAdd_8U_23U_is_a_greater_lor_14_lpi_1_dfm_1_mx0w4 = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_13_itm_23_1)
      & alu_loop_op_14_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2) | alu_loop_op_14_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_14_mx0w0 = (~ FpCmp_8U_23U_false_is_abs_a_greater_15_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_15_lpi_1_dfm_3;
  assign FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_14_mx0w1 = FpCmp_8U_23U_false_is_abs_a_greater_15_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_15_lpi_1_dfm_3;
  assign FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_14_mx0w2 = (~ FpCmp_8U_23U_true_is_abs_a_greater_15_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_15_lpi_1_dfm_3;
  assign FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_14_mx0w3 = FpCmp_8U_23U_true_is_abs_a_greater_15_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_15_lpi_1_dfm_3;
  assign FpAdd_8U_23U_is_a_greater_lor_15_lpi_1_dfm_1_mx0w4 = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_14_itm_23_1)
      & alu_loop_op_15_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2) | alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_15_mx0w0 = (~ FpCmp_8U_23U_false_is_abs_a_greater_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_lpi_1_dfm_3;
  assign FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_15_mx0w1 = FpCmp_8U_23U_false_is_abs_a_greater_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_lpi_1_dfm_3;
  assign FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_15_mx0w2 = (~ FpCmp_8U_23U_true_is_abs_a_greater_lpi_1_dfm_1)
      & alu_nan_to_zero_op_sign_lpi_1_dfm_3;
  assign FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_15_mx0w3 = FpCmp_8U_23U_true_is_abs_a_greater_lpi_1_dfm_1
      | alu_nan_to_zero_op_sign_lpi_1_dfm_3;
  assign FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w4 = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_15_itm_23_1)
      & alu_loop_op_16_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2) | alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_177_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_1_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_65_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_177_nl), 10'b1111111111,
      IsInf_5U_23U_land_1_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_22_13_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_1_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_65_mx0w1,
      or_dcpl_391);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_nl = MUX_v_3_2_2(3'b000,
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_sva_2[12:10]), (FpExpoWidthInc_5U_8U_23U_1U_1U_not_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_nl),
      3'b111, IsInf_5U_23U_land_1_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_nl),
      3'b111, IsNaN_5U_23U_land_1_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_179_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_1_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_64_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_179_nl), 10'b1111111111,
      IsInf_5U_23U_land_1_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_9_0_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_1_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_64_mx0w1,
      or_dcpl_391);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_181_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_2_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_67_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_181_nl), 10'b1111111111,
      IsInf_5U_23U_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_22_13_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_2_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_67_mx0w1,
      or_dcpl_411);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_1_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_65_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_1_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_1_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_65_nl),
      3'b111, IsInf_5U_23U_land_2_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_1_nl),
      3'b111, IsNaN_5U_23U_land_2_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_145_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_2_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_66_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_145_nl), 10'b1111111111,
      IsInf_5U_23U_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_9_0_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_2_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_66_mx0w1,
      or_dcpl_411);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_184_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_3_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_69_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_184_nl), 10'b1111111111,
      IsInf_5U_23U_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_22_13_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_3_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_69_mx0w1,
      or_dcpl_429);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_2_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_66_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_2_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_66_nl),
      3'b111, IsInf_5U_23U_land_3_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_nl),
      3'b111, IsNaN_5U_23U_land_3_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_147_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_3_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_68_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_147_nl), 10'b1111111111,
      IsInf_5U_23U_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_9_0_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_3_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_68_mx0w1,
      or_dcpl_429);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_187_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_4_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_71_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_187_nl), 10'b1111111111,
      IsInf_5U_23U_land_4_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_22_13_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_4_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_71_mx0w1,
      or_dcpl_447);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_3_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_67_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_3_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_3_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_67_nl),
      3'b111, IsInf_5U_23U_land_4_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_3_nl),
      3'b111, IsNaN_5U_23U_land_4_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_149_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_4_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_70_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_149_nl), 10'b1111111111,
      IsInf_5U_23U_land_4_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_9_0_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_4_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_70_mx0w1,
      or_dcpl_447);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_190_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_5_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_73_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_190_nl), 10'b1111111111,
      IsInf_5U_23U_land_5_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_22_13_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_5_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_73_mx0w1,
      or_dcpl_465);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_4_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_68_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_4_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_68_nl),
      3'b111, IsInf_5U_23U_land_5_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_nl),
      3'b111, IsNaN_5U_23U_land_5_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_151_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_5_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_72_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_151_nl), 10'b1111111111,
      IsInf_5U_23U_land_5_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_9_0_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_5_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_72_mx0w1,
      or_dcpl_465);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_193_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_6_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_75_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_193_nl), 10'b1111111111,
      IsInf_5U_23U_land_6_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_22_13_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_6_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_75_mx0w1,
      or_dcpl_483);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_5_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_69_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_5_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_5_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_69_nl),
      3'b111, IsInf_5U_23U_land_6_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_5_nl),
      3'b111, IsNaN_5U_23U_land_6_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_153_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_6_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_74_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_153_nl), 10'b1111111111,
      IsInf_5U_23U_land_6_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_9_0_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_6_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_74_mx0w1,
      or_dcpl_483);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_196_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_7_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_77_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_196_nl), 10'b1111111111,
      IsInf_5U_23U_land_7_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_22_13_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_7_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_77_mx0w1,
      or_dcpl_501);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_6_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_70_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_6_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_70_nl),
      3'b111, IsInf_5U_23U_land_7_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_nl),
      3'b111, IsNaN_5U_23U_land_7_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_155_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_7_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_76_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_155_nl), 10'b1111111111,
      IsInf_5U_23U_land_7_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_9_0_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_7_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_76_mx0w1,
      or_dcpl_501);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_199_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_8_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_79_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_199_nl), 10'b1111111111,
      IsInf_5U_23U_land_8_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_22_13_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_8_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_79_mx0w1,
      or_dcpl_519);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_7_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_71_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_7_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_7_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_71_nl),
      3'b111, IsInf_5U_23U_land_8_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_7_nl),
      3'b111, IsNaN_5U_23U_land_8_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_157_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_8_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_78_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_157_nl), 10'b1111111111,
      IsInf_5U_23U_land_8_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_9_0_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_8_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_78_mx0w1,
      or_dcpl_519);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_202_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_9_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_16_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_81_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_202_nl), 10'b1111111111,
      IsInf_5U_23U_land_9_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_22_13_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_9_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_81_mx0w1,
      or_dcpl_537);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_8_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_16_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_72_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_8_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_72_nl),
      3'b111, IsInf_5U_23U_land_9_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_nl),
      3'b111, IsNaN_5U_23U_land_9_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_159_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_9_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_16_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_80_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_159_nl), 10'b1111111111,
      IsInf_5U_23U_land_9_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_9_0_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_9_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_80_mx0w1,
      or_dcpl_537);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_205_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_10_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_18_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_83_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_205_nl), 10'b1111111111,
      IsInf_5U_23U_land_10_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_22_13_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_10_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_83_mx0w1,
      or_dcpl_555);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_9_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_18_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_73_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_9_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_9_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_73_nl),
      3'b111, IsInf_5U_23U_land_10_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_9_nl),
      3'b111, IsNaN_5U_23U_land_10_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_161_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_10_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_18_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_82_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_161_nl), 10'b1111111111,
      IsInf_5U_23U_land_10_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_9_0_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_10_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_82_mx0w1,
      or_dcpl_555);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_208_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_11_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_20_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_85_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_208_nl), 10'b1111111111,
      IsInf_5U_23U_land_11_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_22_13_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_11_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_85_mx0w1,
      or_dcpl_573);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_10_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_20_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_74_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_10_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_74_nl),
      3'b111, IsInf_5U_23U_land_11_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_nl),
      3'b111, IsNaN_5U_23U_land_11_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_163_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_11_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_20_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_84_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_163_nl), 10'b1111111111,
      IsInf_5U_23U_land_11_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_9_0_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_11_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_84_mx0w1,
      or_dcpl_573);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_211_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_12_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_22_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_87_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_211_nl), 10'b1111111111,
      IsInf_5U_23U_land_12_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_22_13_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_12_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_87_mx0w1,
      or_dcpl_591);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_11_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_22_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_75_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_11_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_11_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_75_nl),
      3'b111, IsInf_5U_23U_land_12_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_11_nl),
      3'b111, IsNaN_5U_23U_land_12_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_165_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_12_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_22_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_86_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_165_nl), 10'b1111111111,
      IsInf_5U_23U_land_12_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_9_0_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_12_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_86_mx0w1,
      or_dcpl_591);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_214_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_13_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_24_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_89_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_214_nl), 10'b1111111111,
      IsInf_5U_23U_land_13_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_22_13_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_13_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_89_mx0w1,
      or_dcpl_609);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_12_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_24_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_76_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_12_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_76_nl),
      3'b111, IsInf_5U_23U_land_13_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_nl),
      3'b111, IsNaN_5U_23U_land_13_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_167_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_13_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_24_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_88_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_167_nl), 10'b1111111111,
      IsInf_5U_23U_land_13_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_9_0_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_13_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_88_mx0w1,
      or_dcpl_609);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_217_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_14_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_26_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_91_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_217_nl), 10'b1111111111,
      IsInf_5U_23U_land_14_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_22_13_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_14_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_91_mx0w1,
      or_dcpl_627);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_13_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_26_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_77_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_13_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_13_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_77_nl),
      3'b111, IsInf_5U_23U_land_14_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_13_nl),
      3'b111, IsNaN_5U_23U_land_14_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_169_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_14_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_26_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_90_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_169_nl), 10'b1111111111,
      IsInf_5U_23U_land_14_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_9_0_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_14_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_90_mx0w1,
      or_dcpl_627);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_220_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_15_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_28_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_93_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_220_nl), 10'b1111111111,
      IsInf_5U_23U_land_15_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_22_13_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_15_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_93_mx0w1,
      or_dcpl_645);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_14_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_28_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_78_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_14_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_78_nl),
      3'b111, IsInf_5U_23U_land_15_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_nl),
      3'b111, IsNaN_5U_23U_land_15_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_171_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_15_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_28_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_92_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_171_nl), 10'b1111111111,
      IsInf_5U_23U_land_15_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_9_0_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_15_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_92_mx0w1,
      or_dcpl_645);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_223_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_30_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_95_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_223_nl), 10'b1111111111,
      IsInf_5U_23U_land_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_22_13_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_95_mx0w1,
      or_dcpl_663);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_15_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_30_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_79_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_15_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_15_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_79_nl),
      3'b111, IsInf_5U_23U_land_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_15_nl),
      3'b111, IsNaN_5U_23U_land_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_173_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_30_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_94_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_173_nl), 10'b1111111111,
      IsInf_5U_23U_land_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_9_0_mx2 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_94_mx0w1,
      or_dcpl_663);
  assign IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0 = ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_12_10_mx0w0!=3'b000) |
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_9_0_mx2!=10'b0000000000))
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_mx0w0==4'b1111) &
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_8U_23U_3_land_15_lpi_1_dfm_mx0w0 = ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_9_0_mx2!=10'b0000000000))
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_mx0w0==4'b1111)
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_8U_23U_3_land_14_lpi_1_dfm_mx0w0 = ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_9_0_mx2!=10'b0000000000))
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_mx0w0==4'b1111)
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_8U_23U_3_land_13_lpi_1_dfm_mx0w0 = ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_9_0_mx2!=10'b0000000000))
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_mx0w0==4'b1111)
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_8U_23U_3_land_12_lpi_1_dfm_mx0w0 = ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_9_0_mx2!=10'b0000000000))
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_mx0w0==4'b1111)
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_8U_23U_3_land_11_lpi_1_dfm_mx0w0 = ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_9_0_mx2!=10'b0000000000))
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_mx0w0==4'b1111)
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_8U_23U_3_land_10_lpi_1_dfm_mx0w0 = ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_9_0_mx2!=10'b0000000000))
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_mx0w0==4'b1111)
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_8U_23U_3_land_9_lpi_1_dfm_mx0w0 = ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_9_0_mx2!=10'b0000000000))
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_mx0w0==4'b1111)
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_8U_23U_3_land_8_lpi_1_dfm_mx0w0 = ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_9_0_mx2!=10'b0000000000))
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_mx0w0==4'b1111)
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_8U_23U_3_land_7_lpi_1_dfm_mx0w0 = ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_9_0_mx2!=10'b0000000000))
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_mx0w0==4'b1111)
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_8U_23U_3_land_6_lpi_1_dfm_mx0w0 = ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_9_0_mx2!=10'b0000000000))
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_mx0w0==4'b1111)
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_8U_23U_3_land_5_lpi_1_dfm_mx0w0 = ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_9_0_mx2!=10'b0000000000))
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_mx0w0==4'b1111)
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_8U_23U_3_land_4_lpi_1_dfm_mx0w0 = ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_9_0_mx2!=10'b0000000000))
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_mx0w0==4'b1111)
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_8U_23U_3_land_3_lpi_1_dfm_mx0w0 = ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_9_0_mx2!=10'b0000000000))
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_mx0w0==4'b1111)
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_8U_23U_3_land_2_lpi_1_dfm_mx0w0 = ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_9_0_mx2!=10'b0000000000))
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_mx0w0==4'b1111)
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_8U_23U_3_land_1_lpi_1_dfm_mx0w0 = ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_22_13_mx2!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_9_0_mx2!=10'b0000000000))
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_mx0w0==4'b1111)
      & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w0==4'b1111);
  assign alu_nan_to_zero_op_sign_1_lpi_1_dfm_mx0w0 = else_AluOp_data_0_15_lpi_1_dfm_mx0
      & (~ alu_nan_to_zero_land_1_lpi_1_dfm);
  assign alu_nan_to_zero_op_sign_2_lpi_1_dfm_mx0w0 = else_AluOp_data_1_15_lpi_1_dfm_mx0
      & (~ alu_nan_to_zero_land_2_lpi_1_dfm);
  assign alu_nan_to_zero_op_sign_3_lpi_1_dfm_mx0w0 = else_AluOp_data_2_15_lpi_1_dfm_mx0
      & (~ alu_nan_to_zero_land_3_lpi_1_dfm);
  assign alu_nan_to_zero_op_sign_4_lpi_1_dfm_mx0w0 = else_AluOp_data_3_15_lpi_1_dfm_mx0
      & (~ alu_nan_to_zero_land_4_lpi_1_dfm);
  assign alu_nan_to_zero_op_sign_5_lpi_1_dfm_mx0w0 = else_AluOp_data_4_15_lpi_1_dfm_mx0
      & (~ alu_nan_to_zero_land_5_lpi_1_dfm);
  assign alu_nan_to_zero_op_sign_6_lpi_1_dfm_mx0w0 = else_AluOp_data_5_15_lpi_1_dfm_mx0
      & (~ alu_nan_to_zero_land_6_lpi_1_dfm);
  assign alu_nan_to_zero_op_sign_7_lpi_1_dfm_mx0w0 = else_AluOp_data_6_15_lpi_1_dfm_mx0
      & (~ alu_nan_to_zero_land_7_lpi_1_dfm);
  assign alu_nan_to_zero_op_sign_8_lpi_1_dfm_mx0w0 = else_AluOp_data_7_15_lpi_1_dfm_mx0
      & (~ alu_nan_to_zero_land_8_lpi_1_dfm);
  assign alu_nan_to_zero_op_sign_9_lpi_1_dfm_mx0w0 = else_AluOp_data_8_15_lpi_1_dfm_mx0
      & (~ alu_nan_to_zero_land_9_lpi_1_dfm);
  assign alu_nan_to_zero_op_sign_10_lpi_1_dfm_mx0w0 = else_AluOp_data_9_15_lpi_1_dfm_mx0
      & (~ alu_nan_to_zero_land_10_lpi_1_dfm);
  assign alu_nan_to_zero_op_sign_11_lpi_1_dfm_mx0w0 = else_AluOp_data_10_15_lpi_1_dfm_mx0
      & (~ alu_nan_to_zero_land_11_lpi_1_dfm);
  assign alu_nan_to_zero_op_sign_12_lpi_1_dfm_mx0w0 = else_AluOp_data_11_15_lpi_1_dfm_mx0
      & (~ alu_nan_to_zero_land_12_lpi_1_dfm);
  assign alu_nan_to_zero_op_sign_13_lpi_1_dfm_mx0w0 = else_AluOp_data_12_15_lpi_1_dfm_mx0
      & (~ alu_nan_to_zero_land_13_lpi_1_dfm);
  assign alu_nan_to_zero_op_sign_14_lpi_1_dfm_mx0w0 = else_AluOp_data_13_15_lpi_1_dfm_mx0
      & (~ alu_nan_to_zero_land_14_lpi_1_dfm);
  assign alu_nan_to_zero_op_sign_15_lpi_1_dfm_mx0w0 = else_AluOp_data_14_15_lpi_1_dfm_mx0
      & (~ alu_nan_to_zero_land_15_lpi_1_dfm);
  assign alu_nan_to_zero_op_sign_lpi_1_dfm_mx0w0 = else_AluOp_data_15_15_lpi_1_dfm_mx0
      & (~ alu_nan_to_zero_land_lpi_1_dfm);
  assign IntShiftLeft_16U_6U_32U_return_0_1_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_1_sva[0])
      | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_1_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_1_sva);
  assign alu_loop_op_1_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftLeft_16U_6U_32U_mbits_fixed_1_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_1_sva));
  assign IntShiftLeft_16U_6U_32U_return_30_1_1_sva_mx0w0 = ~(MUX_v_30_2_2((alu_loop_op_1_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_1_sva));
  assign IntShiftLeft_16U_6U_32U_return_31_1_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_1_sva[31])
      | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_1_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_1_sva);
  assign IntShiftLeft_16U_6U_32U_return_0_2_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_2_sva[0])
      | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_2_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_2_sva);
  assign alu_loop_op_2_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl = ~(MUX_v_30_2_2((IntShiftLeft_16U_6U_32U_mbits_fixed_2_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_2_sva));
  assign IntShiftLeft_16U_6U_32U_return_30_1_2_sva_mx0w0 = ~(MUX_v_30_2_2((alu_loop_op_2_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_2_sva));
  assign IntShiftLeft_16U_6U_32U_return_31_2_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_2_sva[31])
      | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_2_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_2_sva);
  assign IntShiftLeft_16U_6U_32U_return_0_3_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_3_sva[0])
      | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_3_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_3_sva);
  assign alu_loop_op_3_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftLeft_16U_6U_32U_mbits_fixed_3_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_3_sva));
  assign IntShiftLeft_16U_6U_32U_return_30_1_3_sva_mx0w0 = ~(MUX_v_30_2_2((alu_loop_op_3_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_3_sva));
  assign IntShiftLeft_16U_6U_32U_return_31_3_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_3_sva[31])
      | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_3_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_3_sva);
  assign IntShiftLeft_16U_6U_32U_return_0_4_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_4_sva[0])
      | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_4_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_4_sva);
  assign alu_loop_op_4_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl = ~(MUX_v_30_2_2((IntShiftLeft_16U_6U_32U_mbits_fixed_4_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_4_sva));
  assign IntShiftLeft_16U_6U_32U_return_30_1_4_sva_mx0w0 = ~(MUX_v_30_2_2((alu_loop_op_4_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_4_sva));
  assign IntShiftLeft_16U_6U_32U_return_31_4_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_4_sva[31])
      | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_4_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_4_sva);
  assign IntShiftLeft_16U_6U_32U_return_0_5_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_5_sva[0])
      | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_5_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_5_sva);
  assign alu_loop_op_5_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftLeft_16U_6U_32U_mbits_fixed_5_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_5_sva));
  assign IntShiftLeft_16U_6U_32U_return_30_1_5_sva_mx0w0 = ~(MUX_v_30_2_2((alu_loop_op_5_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_5_sva));
  assign IntShiftLeft_16U_6U_32U_return_31_5_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_5_sva[31])
      | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_5_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_5_sva);
  assign IntShiftLeft_16U_6U_32U_return_0_6_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_6_sva[0])
      | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_6_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_6_sva);
  assign alu_loop_op_6_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl = ~(MUX_v_30_2_2((IntShiftLeft_16U_6U_32U_mbits_fixed_6_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_6_sva));
  assign IntShiftLeft_16U_6U_32U_return_30_1_6_sva_mx0w0 = ~(MUX_v_30_2_2((alu_loop_op_6_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_6_sva));
  assign IntShiftLeft_16U_6U_32U_return_31_6_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_6_sva[31])
      | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_6_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_6_sva);
  assign IntShiftLeft_16U_6U_32U_return_0_7_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_7_sva[0])
      | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_7_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_7_sva);
  assign alu_loop_op_7_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftLeft_16U_6U_32U_mbits_fixed_7_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_7_sva));
  assign IntShiftLeft_16U_6U_32U_return_30_1_7_sva_mx0w0 = ~(MUX_v_30_2_2((alu_loop_op_7_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_7_sva));
  assign IntShiftLeft_16U_6U_32U_return_31_7_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_7_sva[31])
      | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_7_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_7_sva);
  assign IntShiftLeft_16U_6U_32U_return_0_8_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_8_sva[0])
      | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_8_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_8_sva);
  assign alu_loop_op_8_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl = ~(MUX_v_30_2_2((IntShiftLeft_16U_6U_32U_mbits_fixed_8_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_8_sva));
  assign IntShiftLeft_16U_6U_32U_return_30_1_8_sva_mx0w0 = ~(MUX_v_30_2_2((alu_loop_op_8_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_8_sva));
  assign IntShiftLeft_16U_6U_32U_return_31_8_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_8_sva[31])
      | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_8_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_8_sva);
  assign IntShiftLeft_16U_6U_32U_return_0_9_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_9_sva[0])
      | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_9_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_9_sva);
  assign alu_loop_op_9_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftLeft_16U_6U_32U_mbits_fixed_9_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_9_sva));
  assign IntShiftLeft_16U_6U_32U_return_30_1_9_sva_mx0w0 = ~(MUX_v_30_2_2((alu_loop_op_9_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_9_sva));
  assign IntShiftLeft_16U_6U_32U_return_31_9_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_9_sva[31])
      | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_9_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_9_sva);
  assign IntShiftLeft_16U_6U_32U_return_0_10_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_10_sva[0])
      | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_10_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_10_sva);
  assign alu_loop_op_10_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl = ~(MUX_v_30_2_2((IntShiftLeft_16U_6U_32U_mbits_fixed_10_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_10_sva));
  assign IntShiftLeft_16U_6U_32U_return_30_1_10_sva_mx0w0 = ~(MUX_v_30_2_2((alu_loop_op_10_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_10_sva));
  assign IntShiftLeft_16U_6U_32U_return_31_10_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_10_sva[31])
      | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_10_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_10_sva);
  assign IntShiftLeft_16U_6U_32U_return_0_11_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_11_sva[0])
      | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_11_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_11_sva);
  assign alu_loop_op_11_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftLeft_16U_6U_32U_mbits_fixed_11_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_11_sva));
  assign IntShiftLeft_16U_6U_32U_return_30_1_11_sva_mx0w0 = ~(MUX_v_30_2_2((alu_loop_op_11_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_11_sva));
  assign IntShiftLeft_16U_6U_32U_return_31_11_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_11_sva[31])
      | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_11_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_11_sva);
  assign IntShiftLeft_16U_6U_32U_return_0_12_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_12_sva[0])
      | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_12_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_12_sva);
  assign alu_loop_op_12_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl = ~(MUX_v_30_2_2((IntShiftLeft_16U_6U_32U_mbits_fixed_12_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_12_sva));
  assign IntShiftLeft_16U_6U_32U_return_30_1_12_sva_mx0w0 = ~(MUX_v_30_2_2((alu_loop_op_12_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_12_sva));
  assign IntShiftLeft_16U_6U_32U_return_31_12_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_12_sva[31])
      | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_12_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_12_sva);
  assign IntShiftLeft_16U_6U_32U_return_0_13_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_13_sva[0])
      | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_13_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_13_sva);
  assign alu_loop_op_13_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftLeft_16U_6U_32U_mbits_fixed_13_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_13_sva));
  assign IntShiftLeft_16U_6U_32U_return_30_1_13_sva_mx0w0 = ~(MUX_v_30_2_2((alu_loop_op_13_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_13_sva));
  assign IntShiftLeft_16U_6U_32U_return_31_13_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_13_sva[31])
      | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_13_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_13_sva);
  assign IntShiftLeft_16U_6U_32U_return_0_14_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_14_sva[0])
      | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_14_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_14_sva);
  assign alu_loop_op_14_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl = ~(MUX_v_30_2_2((IntShiftLeft_16U_6U_32U_mbits_fixed_14_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_14_sva));
  assign IntShiftLeft_16U_6U_32U_return_30_1_14_sva_mx0w0 = ~(MUX_v_30_2_2((alu_loop_op_14_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_14_sva));
  assign IntShiftLeft_16U_6U_32U_return_31_14_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_14_sva[31])
      | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_14_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_14_sva);
  assign IntShiftLeft_16U_6U_32U_return_0_15_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_15_sva[0])
      | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_15_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_15_sva);
  assign alu_loop_op_15_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftLeft_16U_6U_32U_mbits_fixed_15_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_15_sva));
  assign IntShiftLeft_16U_6U_32U_return_30_1_15_sva_mx0w0 = ~(MUX_v_30_2_2((alu_loop_op_15_IntShiftLeft_16U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_15_sva));
  assign IntShiftLeft_16U_6U_32U_return_31_15_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_15_sva[31])
      | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_15_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_15_sva);
  assign IntShiftLeft_16U_6U_32U_return_0_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_sva[0])
      | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_sva);
  assign alu_loop_op_16_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl = ~(MUX_v_30_2_2((IntShiftLeft_16U_6U_32U_mbits_fixed_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_sva));
  assign IntShiftLeft_16U_6U_32U_return_30_1_sva_mx0w0 = ~(MUX_v_30_2_2((alu_loop_op_16_IntShiftLeft_16U_6U_32U_obits_fixed_nor_7_nl),
      30'b111111111111111111111111111111, IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_sva));
  assign IntShiftLeft_16U_6U_32U_return_31_sva_mx0w0 = ~((~((IntShiftLeft_16U_6U_32U_mbits_fixed_sva[31])
      | IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_sva)) | IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_sva);
  assign alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = (chn_alu_in_rsci_d_mxwt[30:0]!=31'b0000000000000000000000000000000);
  assign alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = (chn_alu_in_rsci_d_mxwt[62:32]!=31'b0000000000000000000000000000000);
  assign alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = (chn_alu_in_rsci_d_mxwt[94:64]!=31'b0000000000000000000000000000000);
  assign alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = (chn_alu_in_rsci_d_mxwt[126:96]!=31'b0000000000000000000000000000000);
  assign alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = (chn_alu_in_rsci_d_mxwt[158:128]!=31'b0000000000000000000000000000000);
  assign alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = (chn_alu_in_rsci_d_mxwt[190:160]!=31'b0000000000000000000000000000000);
  assign alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = (chn_alu_in_rsci_d_mxwt[222:192]!=31'b0000000000000000000000000000000);
  assign alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = (chn_alu_in_rsci_d_mxwt[254:224]!=31'b0000000000000000000000000000000);
  assign alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = (chn_alu_in_rsci_d_mxwt[286:256]!=31'b0000000000000000000000000000000);
  assign alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = (chn_alu_in_rsci_d_mxwt[318:288]!=31'b0000000000000000000000000000000);
  assign alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = (chn_alu_in_rsci_d_mxwt[350:320]!=31'b0000000000000000000000000000000);
  assign alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = (chn_alu_in_rsci_d_mxwt[414:384]!=31'b0000000000000000000000000000000);
  assign alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = (chn_alu_in_rsci_d_mxwt[446:416]!=31'b0000000000000000000000000000000);
  assign alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = (chn_alu_in_rsci_d_mxwt[478:448]!=31'b0000000000000000000000000000000);
  assign alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = (chn_alu_in_rsci_d_mxwt[510:480]!=31'b0000000000000000000000000000000);
  assign alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = (chn_alu_in_rsci_d_mxwt[382:352]!=31'b0000000000000000000000000000000);
  assign IsNaN_8U_23U_2_land_lpi_1_dfm_mx1w0 = ~((~((chn_alu_in_rsci_d_mxwt[502:480]!=23'b00000000000000000000000)))
      | (chn_alu_in_rsci_d_mxwt[510:503]!=8'b11111111));
  assign IsNaN_8U_23U_2_land_15_lpi_1_dfm_mx1w0 = ~((~((chn_alu_in_rsci_d_mxwt[470:448]!=23'b00000000000000000000000)))
      | (chn_alu_in_rsci_d_mxwt[478:471]!=8'b11111111));
  assign IsNaN_8U_23U_2_land_14_lpi_1_dfm_mx1w0 = ~((~((chn_alu_in_rsci_d_mxwt[438:416]!=23'b00000000000000000000000)))
      | (chn_alu_in_rsci_d_mxwt[446:439]!=8'b11111111));
  assign IsNaN_8U_23U_2_land_13_lpi_1_dfm_mx1w0 = ~((~((chn_alu_in_rsci_d_mxwt[406:384]!=23'b00000000000000000000000)))
      | (chn_alu_in_rsci_d_mxwt[414:407]!=8'b11111111));
  assign IsNaN_8U_23U_2_land_12_lpi_1_dfm_mx1w0 = ~((~((chn_alu_in_rsci_d_mxwt[374:352]!=23'b00000000000000000000000)))
      | (chn_alu_in_rsci_d_mxwt[382:375]!=8'b11111111));
  assign IsNaN_8U_23U_2_land_11_lpi_1_dfm_mx1w0 = ~((~((chn_alu_in_rsci_d_mxwt[342:320]!=23'b00000000000000000000000)))
      | (chn_alu_in_rsci_d_mxwt[350:343]!=8'b11111111));
  assign IsNaN_8U_23U_2_land_10_lpi_1_dfm_mx1w0 = ~((~((chn_alu_in_rsci_d_mxwt[310:288]!=23'b00000000000000000000000)))
      | (chn_alu_in_rsci_d_mxwt[318:311]!=8'b11111111));
  assign IsNaN_8U_23U_2_land_9_lpi_1_dfm_mx1w0 = ~((~((chn_alu_in_rsci_d_mxwt[278:256]!=23'b00000000000000000000000)))
      | (chn_alu_in_rsci_d_mxwt[286:279]!=8'b11111111));
  assign IsNaN_8U_23U_2_land_8_lpi_1_dfm_mx1w0 = ~((~((chn_alu_in_rsci_d_mxwt[246:224]!=23'b00000000000000000000000)))
      | (chn_alu_in_rsci_d_mxwt[254:247]!=8'b11111111));
  assign IsNaN_8U_23U_2_land_7_lpi_1_dfm_mx1w0 = ~((~((chn_alu_in_rsci_d_mxwt[214:192]!=23'b00000000000000000000000)))
      | (chn_alu_in_rsci_d_mxwt[222:215]!=8'b11111111));
  assign IsNaN_8U_23U_2_land_6_lpi_1_dfm_mx1w0 = ~((~((chn_alu_in_rsci_d_mxwt[182:160]!=23'b00000000000000000000000)))
      | (chn_alu_in_rsci_d_mxwt[190:183]!=8'b11111111));
  assign IsNaN_8U_23U_2_land_5_lpi_1_dfm_mx1w0 = ~((~((chn_alu_in_rsci_d_mxwt[150:128]!=23'b00000000000000000000000)))
      | (chn_alu_in_rsci_d_mxwt[158:151]!=8'b11111111));
  assign IsNaN_8U_23U_2_land_4_lpi_1_dfm_mx1w0 = ~((~((chn_alu_in_rsci_d_mxwt[118:96]!=23'b00000000000000000000000)))
      | (chn_alu_in_rsci_d_mxwt[126:119]!=8'b11111111));
  assign IsNaN_8U_23U_2_land_3_lpi_1_dfm_mx1w0 = ~((~((chn_alu_in_rsci_d_mxwt[86:64]!=23'b00000000000000000000000)))
      | (chn_alu_in_rsci_d_mxwt[94:87]!=8'b11111111));
  assign IsNaN_8U_23U_2_land_2_lpi_1_dfm_mx1w0 = ~((~((chn_alu_in_rsci_d_mxwt[54:32]!=23'b00000000000000000000000)))
      | (chn_alu_in_rsci_d_mxwt[62:55]!=8'b11111111));
  assign IsNaN_8U_23U_2_land_1_lpi_1_dfm_mx1w0 = ~((~((chn_alu_in_rsci_d_mxwt[22:0]!=23'b00000000000000000000000)))
      | (chn_alu_in_rsci_d_mxwt[30:23]!=8'b11111111));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl = ({1'b1 , (AluIn_data_sva_501[22:0])})
      + conv_u2u_23_24({(~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp)
      , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp_1) , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp_2)})
      + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl = ({1'b1 , (AluIn_data_sva_501[54:32])})
      + conv_u2u_23_24({(~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp)
      , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp_1) , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp_2)})
      + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl = ({1'b1 , (AluIn_data_sva_501[86:64])})
      + conv_u2u_23_24({(~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp)
      , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp_1) , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp_2)})
      + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl = ({1'b1 , (AluIn_data_sva_501[118:96])})
      + conv_u2u_23_24({(~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp)
      , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp_1) , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp_2)})
      + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_nl = ({1'b1 , (AluIn_data_sva_501[150:128])})
      + conv_u2u_23_24({(~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp)
      , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp_1) , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp_2)})
      + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_5_nl = ({1'b1 , (AluIn_data_sva_501[182:160])})
      + conv_u2u_23_24({(~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp)
      , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp_1) , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp_2)})
      + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_5_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_5_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_5_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_5_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_nl = ({1'b1 , (AluIn_data_sva_501[214:192])})
      + conv_u2u_23_24({(~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp)
      , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp_1) , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp_2)})
      + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_7_nl = ({1'b1 , (AluIn_data_sva_501[246:224])})
      + conv_u2u_23_24({(~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp)
      , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp_1) , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp_2)})
      + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_7_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_7_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_7_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_7_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_nl = ({1'b1 , (AluIn_data_sva_501[278:256])})
      + conv_u2u_23_24({(~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp)
      , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp_1) , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp_2)})
      + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_9_nl = ({1'b1 , (AluIn_data_sva_501[310:288])})
      + conv_u2u_23_24({(~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp)
      , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp_1) , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp_2)})
      + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_9_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_9_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_9_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_9_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_nl = ({1'b1 , (AluIn_data_sva_501[342:320])})
      + conv_u2u_23_24({(~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp)
      , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp_1) , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp_2)})
      + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_11_nl = ({1'b1 , (AluIn_data_sva_501[374:352])})
      + conv_u2u_23_24({(~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp)
      , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp_1) , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp_2)})
      + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_11_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_11_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_11_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_11_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_12_nl = ({1'b1 , (AluIn_data_sva_501[406:384])})
      + conv_u2u_23_24({(~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp)
      , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp_1) , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp_2)})
      + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_12_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_12_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_12_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_12_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_13_nl = ({1'b1 , (AluIn_data_sva_501[438:416])})
      + conv_u2u_23_24({(~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp)
      , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp_1) , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp_2)})
      + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_13_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_13_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_13_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_13_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_14_nl = ({1'b1 , (AluIn_data_sva_501[470:448])})
      + conv_u2u_23_24({(~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp)
      , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp_1) , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp_2)})
      + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_14_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_14_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_14_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_14_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_15_nl = ({1'b1 , (AluIn_data_sva_501[502:480])})
      + conv_u2u_23_24({(~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp)
      , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp_1) , (~ reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp_2)})
      + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_15_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_15_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_15_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_15_nl));
  assign nl_FpAdd_8U_23U_int_mant_p1_1_sva = conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_mx0);
  assign FpAdd_8U_23U_int_mant_p1_1_sva = nl_FpAdd_8U_23U_int_mant_p1_1_sva[49:0];
  assign FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_91_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_1_sva, FpCmp_8U_23U_false_is_a_greater_1_lpi_1_dfm_7);
  assign FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_1_sva,
      FpAdd_8U_23U_addend_larger_asn_91_mx0w1, FpCmp_8U_23U_false_is_a_greater_1_lpi_1_dfm_7);
  assign nl_FpAdd_8U_23U_int_mant_p1_2_sva = conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_mx0);
  assign FpAdd_8U_23U_int_mant_p1_2_sva = nl_FpAdd_8U_23U_int_mant_p1_2_sva[49:0];
  assign FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_85_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_2_sva, FpCmp_8U_23U_false_is_a_greater_2_lpi_1_dfm_7);
  assign FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_2_sva,
      FpAdd_8U_23U_addend_larger_asn_85_mx0w1, FpCmp_8U_23U_false_is_a_greater_2_lpi_1_dfm_7);
  assign nl_FpAdd_8U_23U_int_mant_p1_3_sva = conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_mx0);
  assign FpAdd_8U_23U_int_mant_p1_3_sva = nl_FpAdd_8U_23U_int_mant_p1_3_sva[49:0];
  assign FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_79_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_3_sva, FpCmp_8U_23U_false_is_a_greater_3_lpi_1_dfm_7);
  assign FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_3_sva,
      FpAdd_8U_23U_addend_larger_asn_79_mx0w1, FpCmp_8U_23U_false_is_a_greater_3_lpi_1_dfm_7);
  assign nl_FpAdd_8U_23U_int_mant_p1_4_sva = conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_4_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_addend_smaller_qr_4_lpi_1_dfm_mx0);
  assign FpAdd_8U_23U_int_mant_p1_4_sva = nl_FpAdd_8U_23U_int_mant_p1_4_sva[49:0];
  assign FpAdd_8U_23U_addend_larger_qr_4_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_73_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_4_sva, FpCmp_8U_23U_false_is_a_greater_4_lpi_1_dfm_7);
  assign FpAdd_8U_23U_addend_smaller_qr_4_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_4_sva,
      FpAdd_8U_23U_addend_larger_asn_73_mx0w1, FpCmp_8U_23U_false_is_a_greater_4_lpi_1_dfm_7);
  assign nl_FpAdd_8U_23U_int_mant_p1_5_sva = conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_5_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_addend_smaller_qr_5_lpi_1_dfm_mx0);
  assign FpAdd_8U_23U_int_mant_p1_5_sva = nl_FpAdd_8U_23U_int_mant_p1_5_sva[49:0];
  assign FpAdd_8U_23U_addend_larger_qr_5_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_67_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_5_sva, FpCmp_8U_23U_false_is_a_greater_5_lpi_1_dfm_7);
  assign FpAdd_8U_23U_addend_smaller_qr_5_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_5_sva,
      FpAdd_8U_23U_addend_larger_asn_67_mx0w1, FpCmp_8U_23U_false_is_a_greater_5_lpi_1_dfm_7);
  assign nl_FpAdd_8U_23U_int_mant_p1_6_sva = conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_6_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_addend_smaller_qr_6_lpi_1_dfm_mx0);
  assign FpAdd_8U_23U_int_mant_p1_6_sva = nl_FpAdd_8U_23U_int_mant_p1_6_sva[49:0];
  assign FpAdd_8U_23U_addend_larger_qr_6_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_61_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_6_sva, FpCmp_8U_23U_false_is_a_greater_6_lpi_1_dfm_7);
  assign FpAdd_8U_23U_addend_smaller_qr_6_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_6_sva,
      FpAdd_8U_23U_addend_larger_asn_61_mx0w1, FpCmp_8U_23U_false_is_a_greater_6_lpi_1_dfm_7);
  assign nl_FpAdd_8U_23U_int_mant_p1_7_sva = conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_7_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_addend_smaller_qr_7_lpi_1_dfm_mx0);
  assign FpAdd_8U_23U_int_mant_p1_7_sva = nl_FpAdd_8U_23U_int_mant_p1_7_sva[49:0];
  assign FpAdd_8U_23U_addend_larger_qr_7_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_55_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_7_sva, FpCmp_8U_23U_false_is_a_greater_7_lpi_1_dfm_7);
  assign FpAdd_8U_23U_addend_smaller_qr_7_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_7_sva,
      FpAdd_8U_23U_addend_larger_asn_55_mx0w1, FpCmp_8U_23U_false_is_a_greater_7_lpi_1_dfm_7);
  assign nl_FpAdd_8U_23U_int_mant_p1_8_sva = conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_8_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_addend_smaller_qr_8_lpi_1_dfm_mx0);
  assign FpAdd_8U_23U_int_mant_p1_8_sva = nl_FpAdd_8U_23U_int_mant_p1_8_sva[49:0];
  assign FpAdd_8U_23U_addend_larger_qr_8_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_49_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_8_sva, FpCmp_8U_23U_false_is_a_greater_8_lpi_1_dfm_7);
  assign FpAdd_8U_23U_addend_smaller_qr_8_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_8_sva,
      FpAdd_8U_23U_addend_larger_asn_49_mx0w1, FpCmp_8U_23U_false_is_a_greater_8_lpi_1_dfm_7);
  assign nl_FpAdd_8U_23U_int_mant_p1_9_sva = conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_9_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_addend_smaller_qr_9_lpi_1_dfm_mx0);
  assign FpAdd_8U_23U_int_mant_p1_9_sva = nl_FpAdd_8U_23U_int_mant_p1_9_sva[49:0];
  assign FpAdd_8U_23U_addend_larger_qr_9_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_43_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_9_sva, FpCmp_8U_23U_false_is_a_greater_9_lpi_1_dfm_7);
  assign FpAdd_8U_23U_addend_smaller_qr_9_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_9_sva,
      FpAdd_8U_23U_addend_larger_asn_43_mx0w1, FpCmp_8U_23U_false_is_a_greater_9_lpi_1_dfm_7);
  assign nl_FpAdd_8U_23U_int_mant_p1_10_sva = conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_10_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_addend_smaller_qr_10_lpi_1_dfm_mx0);
  assign FpAdd_8U_23U_int_mant_p1_10_sva = nl_FpAdd_8U_23U_int_mant_p1_10_sva[49:0];
  assign FpAdd_8U_23U_addend_larger_qr_10_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_37_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_10_sva, FpCmp_8U_23U_false_is_a_greater_10_lpi_1_dfm_7);
  assign FpAdd_8U_23U_addend_smaller_qr_10_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_10_sva,
      FpAdd_8U_23U_addend_larger_asn_37_mx0w1, FpCmp_8U_23U_false_is_a_greater_10_lpi_1_dfm_7);
  assign nl_FpAdd_8U_23U_int_mant_p1_11_sva = conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_11_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_addend_smaller_qr_11_lpi_1_dfm_mx0);
  assign FpAdd_8U_23U_int_mant_p1_11_sva = nl_FpAdd_8U_23U_int_mant_p1_11_sva[49:0];
  assign FpAdd_8U_23U_addend_larger_qr_11_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_31_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_11_sva, FpCmp_8U_23U_false_is_a_greater_11_lpi_1_dfm_7);
  assign FpAdd_8U_23U_addend_smaller_qr_11_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_11_sva,
      FpAdd_8U_23U_addend_larger_asn_31_mx0w1, FpCmp_8U_23U_false_is_a_greater_11_lpi_1_dfm_7);
  assign nl_FpAdd_8U_23U_int_mant_p1_12_sva = conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_12_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_addend_smaller_qr_12_lpi_1_dfm_mx0);
  assign FpAdd_8U_23U_int_mant_p1_12_sva = nl_FpAdd_8U_23U_int_mant_p1_12_sva[49:0];
  assign FpAdd_8U_23U_addend_larger_qr_12_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_25_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_12_sva, FpCmp_8U_23U_false_is_a_greater_12_lpi_1_dfm_7);
  assign FpAdd_8U_23U_addend_smaller_qr_12_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_12_sva,
      FpAdd_8U_23U_addend_larger_asn_25_mx0w1, FpCmp_8U_23U_false_is_a_greater_12_lpi_1_dfm_7);
  assign nl_FpAdd_8U_23U_int_mant_p1_13_sva = conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_13_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_addend_smaller_qr_13_lpi_1_dfm_mx0);
  assign FpAdd_8U_23U_int_mant_p1_13_sva = nl_FpAdd_8U_23U_int_mant_p1_13_sva[49:0];
  assign FpAdd_8U_23U_addend_larger_qr_13_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_19_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_13_sva, FpCmp_8U_23U_false_is_a_greater_13_lpi_1_dfm_7);
  assign FpAdd_8U_23U_addend_smaller_qr_13_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_13_sva,
      FpAdd_8U_23U_addend_larger_asn_19_mx0w1, FpCmp_8U_23U_false_is_a_greater_13_lpi_1_dfm_7);
  assign nl_FpAdd_8U_23U_int_mant_p1_14_sva = conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_14_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_addend_smaller_qr_14_lpi_1_dfm_mx0);
  assign FpAdd_8U_23U_int_mant_p1_14_sva = nl_FpAdd_8U_23U_int_mant_p1_14_sva[49:0];
  assign FpAdd_8U_23U_addend_larger_qr_14_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_13_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_14_sva, FpCmp_8U_23U_false_is_a_greater_14_lpi_1_dfm_7);
  assign FpAdd_8U_23U_addend_smaller_qr_14_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_14_sva,
      FpAdd_8U_23U_addend_larger_asn_13_mx0w1, FpCmp_8U_23U_false_is_a_greater_14_lpi_1_dfm_7);
  assign nl_FpAdd_8U_23U_int_mant_p1_15_sva = conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_15_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_addend_smaller_qr_15_lpi_1_dfm_mx0);
  assign FpAdd_8U_23U_int_mant_p1_15_sva = nl_FpAdd_8U_23U_int_mant_p1_15_sva[49:0];
  assign FpAdd_8U_23U_addend_larger_qr_15_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_7_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_15_sva, FpCmp_8U_23U_false_is_a_greater_15_lpi_1_dfm_7);
  assign FpAdd_8U_23U_addend_smaller_qr_15_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_15_sva,
      FpAdd_8U_23U_addend_larger_asn_7_mx0w1, FpCmp_8U_23U_false_is_a_greater_15_lpi_1_dfm_7);
  assign nl_FpAdd_8U_23U_int_mant_p1_sva = conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_mx0);
  assign FpAdd_8U_23U_int_mant_p1_sva = nl_FpAdd_8U_23U_int_mant_p1_sva[49:0];
  assign FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_1_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_sva, FpCmp_8U_23U_false_is_a_greater_lpi_1_dfm_7);
  assign FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_sva,
      FpAdd_8U_23U_addend_larger_asn_1_mx0w1, FpCmp_8U_23U_false_is_a_greater_lpi_1_dfm_7);
  assign alu_loop_op_if_alu_loop_op_if_nor_cse = ~(IsNaN_8U_23U_1_land_1_lpi_1_dfm_9
      | IsNaN_8U_23U_land_1_lpi_1_dfm_10);
  assign nl_alu_loop_op_1_FpMantRNE_49U_24U_else_acc_nl = (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_1_sva);
  assign alu_loop_op_1_FpMantRNE_49U_24U_else_acc_nl = nl_alu_loop_op_1_FpMantRNE_49U_24U_else_acc_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_16_nl = MUX_v_23_2_2((alu_loop_op_1_FpMantRNE_49U_24U_else_acc_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_o_mant_1_lpi_1_dfm_2_mx0 = MUX1HOT_v_23_3_2((FpAdd_8U_23U_FpAdd_8U_23U_or_16_nl),
      ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_tmp_2}), (AluIn_data_sva_503[22:0]),
      {alu_loop_op_if_alu_loop_op_if_nor_cse , FpAdd_8U_23U_and_ssc , IsNaN_8U_23U_land_1_lpi_1_dfm_10});
  assign alu_loop_op_if_alu_loop_op_if_nor_1_cse = ~(IsNaN_8U_23U_1_land_2_lpi_1_dfm_9
      | IsNaN_8U_23U_land_2_lpi_1_dfm_10);
  assign nl_alu_loop_op_2_FpMantRNE_49U_24U_else_acc_1_nl = (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_2_sva);
  assign alu_loop_op_2_FpMantRNE_49U_24U_else_acc_1_nl = nl_alu_loop_op_2_FpMantRNE_49U_24U_else_acc_1_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_17_nl = MUX_v_23_2_2((alu_loop_op_2_FpMantRNE_49U_24U_else_acc_1_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_o_mant_2_lpi_1_dfm_2_mx0 = MUX1HOT_v_23_3_2((FpAdd_8U_23U_FpAdd_8U_23U_or_17_nl),
      ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_tmp_2}), (AluIn_data_sva_503[54:32]),
      {alu_loop_op_if_alu_loop_op_if_nor_1_cse , FpAdd_8U_23U_and_2_ssc , IsNaN_8U_23U_land_2_lpi_1_dfm_10});
  assign alu_loop_op_if_alu_loop_op_if_nor_2_cse = ~(IsNaN_8U_23U_1_land_3_lpi_1_dfm_9
      | IsNaN_8U_23U_land_3_lpi_1_dfm_10);
  assign nl_alu_loop_op_3_FpMantRNE_49U_24U_else_acc_nl = (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_3_sva);
  assign alu_loop_op_3_FpMantRNE_49U_24U_else_acc_nl = nl_alu_loop_op_3_FpMantRNE_49U_24U_else_acc_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_18_nl = MUX_v_23_2_2((alu_loop_op_3_FpMantRNE_49U_24U_else_acc_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_o_mant_3_lpi_1_dfm_2_mx0 = MUX1HOT_v_23_3_2((FpAdd_8U_23U_FpAdd_8U_23U_or_18_nl),
      ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_tmp_2}), (AluIn_data_sva_503[86:64]),
      {alu_loop_op_if_alu_loop_op_if_nor_2_cse , FpAdd_8U_23U_and_4_ssc , IsNaN_8U_23U_land_3_lpi_1_dfm_10});
  assign alu_loop_op_if_alu_loop_op_if_nor_3_cse = ~(IsNaN_8U_23U_1_land_4_lpi_1_dfm_9
      | IsNaN_8U_23U_land_4_lpi_1_dfm_10);
  assign nl_alu_loop_op_4_FpMantRNE_49U_24U_else_acc_1_nl = (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_4_sva);
  assign alu_loop_op_4_FpMantRNE_49U_24U_else_acc_1_nl = nl_alu_loop_op_4_FpMantRNE_49U_24U_else_acc_1_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_19_nl = MUX_v_23_2_2((alu_loop_op_4_FpMantRNE_49U_24U_else_acc_1_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_4_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_o_mant_4_lpi_1_dfm_2_mx0 = MUX1HOT_v_23_3_2((FpAdd_8U_23U_FpAdd_8U_23U_or_19_nl),
      ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_tmp_2}), (AluIn_data_sva_503[118:96]),
      {alu_loop_op_if_alu_loop_op_if_nor_3_cse , FpAdd_8U_23U_and_6_ssc , IsNaN_8U_23U_land_4_lpi_1_dfm_10});
  assign alu_loop_op_if_alu_loop_op_if_nor_4_cse = ~(IsNaN_8U_23U_1_land_5_lpi_1_dfm_9
      | IsNaN_8U_23U_land_5_lpi_1_dfm_10);
  assign nl_alu_loop_op_5_FpMantRNE_49U_24U_else_acc_nl = (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_5_sva);
  assign alu_loop_op_5_FpMantRNE_49U_24U_else_acc_nl = nl_alu_loop_op_5_FpMantRNE_49U_24U_else_acc_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_20_nl = MUX_v_23_2_2((alu_loop_op_5_FpMantRNE_49U_24U_else_acc_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_5_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_o_mant_5_lpi_1_dfm_2_mx0 = MUX1HOT_v_23_3_2((FpAdd_8U_23U_FpAdd_8U_23U_or_20_nl),
      ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_tmp_2}), (AluIn_data_sva_503[150:128]),
      {alu_loop_op_if_alu_loop_op_if_nor_4_cse , FpAdd_8U_23U_and_8_ssc , IsNaN_8U_23U_land_5_lpi_1_dfm_10});
  assign alu_loop_op_if_alu_loop_op_if_nor_5_cse = ~(IsNaN_8U_23U_1_land_6_lpi_1_dfm_9
      | IsNaN_8U_23U_land_6_lpi_1_dfm_10);
  assign nl_alu_loop_op_6_FpMantRNE_49U_24U_else_acc_1_nl = (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_6_sva);
  assign alu_loop_op_6_FpMantRNE_49U_24U_else_acc_1_nl = nl_alu_loop_op_6_FpMantRNE_49U_24U_else_acc_1_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_21_nl = MUX_v_23_2_2((alu_loop_op_6_FpMantRNE_49U_24U_else_acc_1_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_6_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_o_mant_6_lpi_1_dfm_2_mx0 = MUX1HOT_v_23_3_2((FpAdd_8U_23U_FpAdd_8U_23U_or_21_nl),
      ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_tmp_2}), (AluIn_data_sva_503[182:160]),
      {alu_loop_op_if_alu_loop_op_if_nor_5_cse , FpAdd_8U_23U_and_10_ssc , IsNaN_8U_23U_land_6_lpi_1_dfm_10});
  assign alu_loop_op_if_alu_loop_op_if_nor_6_cse = ~(IsNaN_8U_23U_1_land_7_lpi_1_dfm_9
      | IsNaN_8U_23U_land_7_lpi_1_dfm_10);
  assign nl_alu_loop_op_7_FpMantRNE_49U_24U_else_acc_nl = (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_7_sva);
  assign alu_loop_op_7_FpMantRNE_49U_24U_else_acc_nl = nl_alu_loop_op_7_FpMantRNE_49U_24U_else_acc_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_22_nl = MUX_v_23_2_2((alu_loop_op_7_FpMantRNE_49U_24U_else_acc_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_7_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_o_mant_7_lpi_1_dfm_2_mx0 = MUX1HOT_v_23_3_2((FpAdd_8U_23U_FpAdd_8U_23U_or_22_nl),
      ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_tmp_2}), (AluIn_data_sva_503[214:192]),
      {alu_loop_op_if_alu_loop_op_if_nor_6_cse , FpAdd_8U_23U_and_12_ssc , IsNaN_8U_23U_land_7_lpi_1_dfm_10});
  assign alu_loop_op_if_alu_loop_op_if_nor_7_cse = ~(IsNaN_8U_23U_1_land_8_lpi_1_dfm_9
      | IsNaN_8U_23U_land_8_lpi_1_dfm_10);
  assign nl_alu_loop_op_8_FpMantRNE_49U_24U_else_acc_1_nl = (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_8_sva);
  assign alu_loop_op_8_FpMantRNE_49U_24U_else_acc_1_nl = nl_alu_loop_op_8_FpMantRNE_49U_24U_else_acc_1_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_23_nl = MUX_v_23_2_2((alu_loop_op_8_FpMantRNE_49U_24U_else_acc_1_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_8_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_o_mant_8_lpi_1_dfm_2_mx0 = MUX1HOT_v_23_3_2((FpAdd_8U_23U_FpAdd_8U_23U_or_23_nl),
      ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_tmp_2}), (AluIn_data_sva_503[246:224]),
      {alu_loop_op_if_alu_loop_op_if_nor_7_cse , FpAdd_8U_23U_and_14_ssc , IsNaN_8U_23U_land_8_lpi_1_dfm_10});
  assign alu_loop_op_if_alu_loop_op_if_nor_8_cse = ~(IsNaN_8U_23U_1_land_9_lpi_1_dfm_9
      | IsNaN_8U_23U_land_9_lpi_1_dfm_10);
  assign nl_alu_loop_op_9_FpMantRNE_49U_24U_else_acc_nl = (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_9_sva);
  assign alu_loop_op_9_FpMantRNE_49U_24U_else_acc_nl = nl_alu_loop_op_9_FpMantRNE_49U_24U_else_acc_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_24_nl = MUX_v_23_2_2((alu_loop_op_9_FpMantRNE_49U_24U_else_acc_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_9_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_o_mant_9_lpi_1_dfm_2_mx0 = MUX1HOT_v_23_3_2((FpAdd_8U_23U_FpAdd_8U_23U_or_24_nl),
      ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_tmp_2}), (AluIn_data_sva_503[278:256]),
      {alu_loop_op_if_alu_loop_op_if_nor_8_cse , FpAdd_8U_23U_and_16_ssc , IsNaN_8U_23U_land_9_lpi_1_dfm_10});
  assign alu_loop_op_if_alu_loop_op_if_nor_9_cse = ~(IsNaN_8U_23U_1_land_10_lpi_1_dfm_9
      | IsNaN_8U_23U_land_10_lpi_1_dfm_10);
  assign nl_alu_loop_op_10_FpMantRNE_49U_24U_else_acc_1_nl = (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_10_sva);
  assign alu_loop_op_10_FpMantRNE_49U_24U_else_acc_1_nl = nl_alu_loop_op_10_FpMantRNE_49U_24U_else_acc_1_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_25_nl = MUX_v_23_2_2((alu_loop_op_10_FpMantRNE_49U_24U_else_acc_1_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_10_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_o_mant_10_lpi_1_dfm_2_mx0 = MUX1HOT_v_23_3_2((FpAdd_8U_23U_FpAdd_8U_23U_or_25_nl),
      ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_tmp_2}), (AluIn_data_sva_503[310:288]),
      {alu_loop_op_if_alu_loop_op_if_nor_9_cse , FpAdd_8U_23U_and_18_ssc , IsNaN_8U_23U_land_10_lpi_1_dfm_10});
  assign alu_loop_op_if_alu_loop_op_if_nor_10_cse = ~(IsNaN_8U_23U_1_land_11_lpi_1_dfm_9
      | IsNaN_8U_23U_land_11_lpi_1_dfm_10);
  assign nl_alu_loop_op_11_FpMantRNE_49U_24U_else_acc_nl = (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_11_sva);
  assign alu_loop_op_11_FpMantRNE_49U_24U_else_acc_nl = nl_alu_loop_op_11_FpMantRNE_49U_24U_else_acc_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_26_nl = MUX_v_23_2_2((alu_loop_op_11_FpMantRNE_49U_24U_else_acc_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_11_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_o_mant_11_lpi_1_dfm_2_mx0 = MUX1HOT_v_23_3_2((FpAdd_8U_23U_FpAdd_8U_23U_or_26_nl),
      ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_tmp_2}), (AluIn_data_sva_503[342:320]),
      {alu_loop_op_if_alu_loop_op_if_nor_10_cse , FpAdd_8U_23U_and_20_ssc , IsNaN_8U_23U_land_11_lpi_1_dfm_10});
  assign alu_loop_op_if_alu_loop_op_if_nor_11_cse = ~(IsNaN_8U_23U_1_land_12_lpi_1_dfm_9
      | IsNaN_8U_23U_land_12_lpi_1_dfm_10);
  assign nl_alu_loop_op_12_FpMantRNE_49U_24U_else_acc_1_nl = (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_12_sva);
  assign alu_loop_op_12_FpMantRNE_49U_24U_else_acc_1_nl = nl_alu_loop_op_12_FpMantRNE_49U_24U_else_acc_1_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_27_nl = MUX_v_23_2_2((alu_loop_op_12_FpMantRNE_49U_24U_else_acc_1_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_12_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_o_mant_12_lpi_1_dfm_2_mx0 = MUX1HOT_v_23_3_2((FpAdd_8U_23U_FpAdd_8U_23U_or_27_nl),
      ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_tmp_2}), (AluIn_data_sva_503[374:352]),
      {alu_loop_op_if_alu_loop_op_if_nor_11_cse , FpAdd_8U_23U_and_22_ssc , IsNaN_8U_23U_land_12_lpi_1_dfm_10});
  assign alu_loop_op_if_alu_loop_op_if_nor_12_cse = ~(IsNaN_8U_23U_1_land_13_lpi_1_dfm_9
      | IsNaN_8U_23U_land_13_lpi_1_dfm_10);
  assign nl_alu_loop_op_13_FpMantRNE_49U_24U_else_acc_nl = (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_13_sva);
  assign alu_loop_op_13_FpMantRNE_49U_24U_else_acc_nl = nl_alu_loop_op_13_FpMantRNE_49U_24U_else_acc_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_28_nl = MUX_v_23_2_2((alu_loop_op_13_FpMantRNE_49U_24U_else_acc_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_13_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_o_mant_13_lpi_1_dfm_2_mx0 = MUX1HOT_v_23_3_2((FpAdd_8U_23U_FpAdd_8U_23U_or_28_nl),
      ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_tmp_2}), (AluIn_data_sva_503[406:384]),
      {alu_loop_op_if_alu_loop_op_if_nor_12_cse , FpAdd_8U_23U_and_24_ssc , IsNaN_8U_23U_land_13_lpi_1_dfm_10});
  assign alu_loop_op_if_alu_loop_op_if_nor_13_cse = ~(IsNaN_8U_23U_1_land_14_lpi_1_dfm_9
      | IsNaN_8U_23U_land_14_lpi_1_dfm_10);
  assign nl_alu_loop_op_14_FpMantRNE_49U_24U_else_acc_1_nl = (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_14_sva);
  assign alu_loop_op_14_FpMantRNE_49U_24U_else_acc_1_nl = nl_alu_loop_op_14_FpMantRNE_49U_24U_else_acc_1_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_29_nl = MUX_v_23_2_2((alu_loop_op_14_FpMantRNE_49U_24U_else_acc_1_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_14_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_o_mant_14_lpi_1_dfm_2_mx0 = MUX1HOT_v_23_3_2((FpAdd_8U_23U_FpAdd_8U_23U_or_29_nl),
      ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_tmp_2}), (AluIn_data_sva_503[438:416]),
      {alu_loop_op_if_alu_loop_op_if_nor_13_cse , FpAdd_8U_23U_and_26_ssc , IsNaN_8U_23U_land_14_lpi_1_dfm_10});
  assign alu_loop_op_if_alu_loop_op_if_nor_14_cse = ~(IsNaN_8U_23U_1_land_15_lpi_1_dfm_9
      | IsNaN_8U_23U_land_15_lpi_1_dfm_10);
  assign nl_alu_loop_op_15_FpMantRNE_49U_24U_else_acc_nl = (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_15_sva);
  assign alu_loop_op_15_FpMantRNE_49U_24U_else_acc_nl = nl_alu_loop_op_15_FpMantRNE_49U_24U_else_acc_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_30_nl = MUX_v_23_2_2((alu_loop_op_15_FpMantRNE_49U_24U_else_acc_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_15_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_o_mant_15_lpi_1_dfm_2_mx0 = MUX1HOT_v_23_3_2((FpAdd_8U_23U_FpAdd_8U_23U_or_30_nl),
      ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_tmp_2}), (AluIn_data_sva_503[470:448]),
      {alu_loop_op_if_alu_loop_op_if_nor_14_cse , FpAdd_8U_23U_and_28_ssc , IsNaN_8U_23U_land_15_lpi_1_dfm_10});
  assign alu_loop_op_if_alu_loop_op_if_nor_15_cse = ~(IsNaN_8U_23U_1_land_lpi_1_dfm_9
      | IsNaN_8U_23U_land_lpi_1_dfm_10);
  assign nl_alu_loop_op_16_FpMantRNE_49U_24U_else_acc_1_nl = (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_sva);
  assign alu_loop_op_16_FpMantRNE_49U_24U_else_acc_1_nl = nl_alu_loop_op_16_FpMantRNE_49U_24U_else_acc_1_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_31_nl = MUX_v_23_2_2((alu_loop_op_16_FpMantRNE_49U_24U_else_acc_1_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_o_mant_lpi_1_dfm_2_mx0 = MUX1HOT_v_23_3_2((FpAdd_8U_23U_FpAdd_8U_23U_or_31_nl),
      ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_tmp_1
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_tmp_2}), (AluIn_data_sva_503[502:480]),
      {alu_loop_op_if_alu_loop_op_if_nor_15_cse , FpAdd_8U_23U_and_30_ssc , IsNaN_8U_23U_land_lpi_1_dfm_10});
  assign alu_loop_op_else_equal_tmp = (cfg_alu_algo_1_sva_7==2'b01);
  assign else_unequal_tmp = ~((cfg_precision==2'b10));
  assign nl_FpAdd_8U_23U_o_expo_1_sva_4 = ({FpAdd_8U_23U_o_expo_1_lpi_1_dfm_2_7_4
      , FpAdd_8U_23U_o_expo_1_lpi_1_dfm_2_3_0}) + 8'b1;
  assign FpAdd_8U_23U_o_expo_1_sva_4 = nl_FpAdd_8U_23U_o_expo_1_sva_4[7:0];
  assign FpAdd_8U_23U_o_expo_1_lpi_1_dfm_1 = MUX_v_8_2_2(8'b00000000, z_out, FpNormalize_8U_49U_oelse_not_33);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_1_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      alu_loop_op_1_FpNormalize_8U_49U_else_lshift_itm, FpNormalize_8U_49U_oelse_not_33);
  assign FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_1_nl),
      (FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49:1]), FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49]);
  assign FpMantRNE_49U_24U_else_carry_1_sva = (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[25]));
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_nl = FpAdd_8U_23U_is_inf_1_lpi_1_dfm
      | (~ alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1);
  assign FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_is_inf_1_lpi_1_dfm,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_nl), alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp);
  assign nl_alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl = ({1'b1 , FpAdd_8U_23U_o_expo_1_lpi_1_dfm_2_7_4
      , (FpAdd_8U_23U_o_expo_1_lpi_1_dfm_2_3_0[3:1])}) + 8'b1;
  assign alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl = nl_alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl[7:0];
  assign alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1 = readslicef_8_1_7((alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl));
  assign FpAdd_8U_23U_o_expo_1_lpi_1_dfm_2_7_4 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_1_lpi_1_dfm_1[7:4]),
      FpAdd_8U_23U_qr_2_lpi_1_dfm_5_7_4_1, (z_out[7:4]), {(~ (FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_256 , FpAdd_8U_23U_asn_258});
  assign FpAdd_8U_23U_is_inf_1_lpi_1_dfm = ~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_2
      | (~ (FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49])));
  assign FpAdd_8U_23U_and_32_tmp = alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1
      & alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp;
  assign alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_else_carry_1_sva
      & (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign nl_FpAdd_8U_23U_o_expo_2_sva_4 = ({FpAdd_8U_23U_o_expo_2_lpi_1_dfm_2_7_4
      , FpAdd_8U_23U_o_expo_2_lpi_1_dfm_2_3_0}) + 8'b1;
  assign FpAdd_8U_23U_o_expo_2_sva_4 = nl_FpAdd_8U_23U_o_expo_2_sva_4[7:0];
  assign FpAdd_8U_23U_o_expo_2_lpi_1_dfm_1 = MUX_v_8_2_2(8'b00000000, z_out_1, FpNormalize_8U_49U_oelse_not_35);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_3_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      alu_loop_op_2_FpNormalize_8U_49U_else_lshift_1_itm, FpNormalize_8U_49U_oelse_not_35);
  assign FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_3_nl),
      (FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49:1]), FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49]);
  assign FpMantRNE_49U_24U_else_carry_2_sva = (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[25]));
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_1_nl = FpAdd_8U_23U_is_inf_2_lpi_1_dfm
      | (~ alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1);
  assign FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_is_inf_2_lpi_1_dfm,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_1_nl), alu_loop_op_2_FpMantRNE_49U_24U_else_and_1_tmp);
  assign nl_alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_2_nl = ({1'b1 , FpAdd_8U_23U_o_expo_2_lpi_1_dfm_2_7_4
      , (FpAdd_8U_23U_o_expo_2_lpi_1_dfm_2_3_0[3:1])}) + 8'b1;
  assign alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_2_nl = nl_alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_2_nl[7:0];
  assign alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1 = readslicef_8_1_7((alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_2_nl));
  assign FpAdd_8U_23U_o_expo_2_lpi_1_dfm_2_7_4 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_2_lpi_1_dfm_1[7:4]),
      FpAdd_8U_23U_qr_3_lpi_1_dfm_5_7_4_1, (z_out_1[7:4]), {(~ (FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_260 , FpAdd_8U_23U_asn_262});
  assign FpAdd_8U_23U_is_inf_2_lpi_1_dfm = ~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_2
      | (~ (FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49])));
  assign FpAdd_8U_23U_and_33_tmp = alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1
      & alu_loop_op_2_FpMantRNE_49U_24U_else_and_1_tmp;
  assign alu_loop_op_2_FpMantRNE_49U_24U_else_and_1_tmp = FpMantRNE_49U_24U_else_carry_2_sva
      & (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign nl_FpAdd_8U_23U_o_expo_3_sva_4 = ({FpAdd_8U_23U_o_expo_3_lpi_1_dfm_2_7_4
      , FpAdd_8U_23U_o_expo_3_lpi_1_dfm_2_3_0}) + 8'b1;
  assign FpAdd_8U_23U_o_expo_3_sva_4 = nl_FpAdd_8U_23U_o_expo_3_sva_4[7:0];
  assign FpAdd_8U_23U_o_expo_3_lpi_1_dfm_1 = MUX_v_8_2_2(8'b00000000, z_out_2, FpNormalize_8U_49U_oelse_not_37);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_5_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      alu_loop_op_3_FpNormalize_8U_49U_else_lshift_itm, FpNormalize_8U_49U_oelse_not_37);
  assign FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_5_nl),
      (FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49:1]), FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49]);
  assign FpMantRNE_49U_24U_else_carry_3_sva = (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[25]));
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_2_nl = FpAdd_8U_23U_is_inf_3_lpi_1_dfm
      | (~ alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1);
  assign FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_is_inf_3_lpi_1_dfm,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_2_nl), alu_loop_op_3_FpMantRNE_49U_24U_else_and_tmp);
  assign nl_alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_1_nl = ({1'b1 , FpAdd_8U_23U_o_expo_3_lpi_1_dfm_2_7_4
      , (FpAdd_8U_23U_o_expo_3_lpi_1_dfm_2_3_0[3:1])}) + 8'b1;
  assign alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_1_nl = nl_alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_1_nl[7:0];
  assign alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1 = readslicef_8_1_7((alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_1_nl));
  assign FpAdd_8U_23U_o_expo_3_lpi_1_dfm_2_7_4 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_3_lpi_1_dfm_1[7:4]),
      FpAdd_8U_23U_qr_4_lpi_1_dfm_5_7_4_1, (z_out_2[7:4]), {(~ (FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_264 , FpAdd_8U_23U_asn_266});
  assign FpAdd_8U_23U_is_inf_3_lpi_1_dfm = ~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_2
      | (~ (FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49])));
  assign FpAdd_8U_23U_and_34_tmp = alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1
      & alu_loop_op_3_FpMantRNE_49U_24U_else_and_tmp;
  assign alu_loop_op_3_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_else_carry_3_sva
      & (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign nl_FpAdd_8U_23U_o_expo_4_sva_4 = ({FpAdd_8U_23U_o_expo_4_lpi_1_dfm_2_7_4
      , FpAdd_8U_23U_o_expo_4_lpi_1_dfm_2_3_0}) + 8'b1;
  assign FpAdd_8U_23U_o_expo_4_sva_4 = nl_FpAdd_8U_23U_o_expo_4_sva_4[7:0];
  assign FpAdd_8U_23U_o_expo_4_lpi_1_dfm_1 = MUX_v_8_2_2(8'b00000000, z_out_3, FpNormalize_8U_49U_oelse_not_39);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_7_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      alu_loop_op_4_FpNormalize_8U_49U_else_lshift_1_itm, FpNormalize_8U_49U_oelse_not_39);
  assign FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_7_nl),
      (FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_5[49:1]), FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_5[49]);
  assign FpMantRNE_49U_24U_else_carry_4_sva = (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[25]));
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_3_nl = FpAdd_8U_23U_is_inf_4_lpi_1_dfm
      | (~ alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1);
  assign FpAdd_8U_23U_is_inf_4_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_is_inf_4_lpi_1_dfm,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_3_nl), alu_loop_op_4_FpMantRNE_49U_24U_else_and_1_tmp);
  assign nl_alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_2_nl = ({1'b1 , FpAdd_8U_23U_o_expo_4_lpi_1_dfm_2_7_4
      , (FpAdd_8U_23U_o_expo_4_lpi_1_dfm_2_3_0[3:1])}) + 8'b1;
  assign alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_2_nl = nl_alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_2_nl[7:0];
  assign alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1 = readslicef_8_1_7((alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_2_nl));
  assign FpAdd_8U_23U_o_expo_4_lpi_1_dfm_2_7_4 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_4_lpi_1_dfm_1[7:4]),
      FpAdd_8U_23U_qr_5_lpi_1_dfm_5_7_4_1, (z_out_3[7:4]), {(~ (FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_268 , FpAdd_8U_23U_asn_270});
  assign FpAdd_8U_23U_is_inf_4_lpi_1_dfm = ~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_4_sva_2
      | (~ (FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_5[49])));
  assign FpAdd_8U_23U_and_35_tmp = alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1
      & alu_loop_op_4_FpMantRNE_49U_24U_else_and_1_tmp;
  assign alu_loop_op_4_FpMantRNE_49U_24U_else_and_1_tmp = FpMantRNE_49U_24U_else_carry_4_sva
      & (FpAdd_8U_23U_int_mant_5_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign nl_FpAdd_8U_23U_o_expo_5_sva_4 = ({FpAdd_8U_23U_o_expo_5_lpi_1_dfm_2_7_4
      , FpAdd_8U_23U_o_expo_5_lpi_1_dfm_2_3_0}) + 8'b1;
  assign FpAdd_8U_23U_o_expo_5_sva_4 = nl_FpAdd_8U_23U_o_expo_5_sva_4[7:0];
  assign FpAdd_8U_23U_o_expo_5_lpi_1_dfm_1 = MUX_v_8_2_2(8'b00000000, z_out_4, FpNormalize_8U_49U_oelse_not_41);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_9_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      alu_loop_op_5_FpNormalize_8U_49U_else_lshift_itm, FpNormalize_8U_49U_oelse_not_41);
  assign FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_9_nl),
      (FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_5[49:1]), FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_5[49]);
  assign FpMantRNE_49U_24U_else_carry_5_sva = (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[25]));
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_4_nl = FpAdd_8U_23U_is_inf_5_lpi_1_dfm
      | (~ alu_loop_op_5_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1);
  assign FpAdd_8U_23U_is_inf_5_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_is_inf_5_lpi_1_dfm,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_4_nl), alu_loop_op_5_FpMantRNE_49U_24U_else_and_tmp);
  assign nl_alu_loop_op_5_FpAdd_8U_23U_if_4_if_acc_1_nl = ({1'b1 , FpAdd_8U_23U_o_expo_5_lpi_1_dfm_2_7_4
      , (FpAdd_8U_23U_o_expo_5_lpi_1_dfm_2_3_0[3:1])}) + 8'b1;
  assign alu_loop_op_5_FpAdd_8U_23U_if_4_if_acc_1_nl = nl_alu_loop_op_5_FpAdd_8U_23U_if_4_if_acc_1_nl[7:0];
  assign alu_loop_op_5_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1 = readslicef_8_1_7((alu_loop_op_5_FpAdd_8U_23U_if_4_if_acc_1_nl));
  assign FpAdd_8U_23U_o_expo_5_lpi_1_dfm_2_7_4 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_5_lpi_1_dfm_1[7:4]),
      FpAdd_8U_23U_qr_6_lpi_1_dfm_5_7_4_1, (z_out_4[7:4]), {(~ (FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_272 , FpAdd_8U_23U_asn_274});
  assign FpAdd_8U_23U_is_inf_5_lpi_1_dfm = ~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_5_sva_2
      | (~ (FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_5[49])));
  assign FpAdd_8U_23U_and_36_tmp = alu_loop_op_5_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1
      & alu_loop_op_5_FpMantRNE_49U_24U_else_and_tmp;
  assign alu_loop_op_5_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_else_carry_5_sva
      & (FpAdd_8U_23U_int_mant_6_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign nl_FpAdd_8U_23U_o_expo_6_sva_4 = ({FpAdd_8U_23U_o_expo_6_lpi_1_dfm_2_7_4
      , FpAdd_8U_23U_o_expo_6_lpi_1_dfm_2_3_0}) + 8'b1;
  assign FpAdd_8U_23U_o_expo_6_sva_4 = nl_FpAdd_8U_23U_o_expo_6_sva_4[7:0];
  assign FpAdd_8U_23U_o_expo_6_lpi_1_dfm_1 = MUX_v_8_2_2(8'b00000000, z_out_5, FpNormalize_8U_49U_oelse_not_43);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_11_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      alu_loop_op_6_FpNormalize_8U_49U_else_lshift_1_itm, FpNormalize_8U_49U_oelse_not_43);
  assign FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_11_nl),
      (FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_5[49:1]), FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_5[49]);
  assign FpMantRNE_49U_24U_else_carry_6_sva = (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[25]));
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_5_nl = FpAdd_8U_23U_is_inf_6_lpi_1_dfm
      | (~ alu_loop_op_6_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1);
  assign FpAdd_8U_23U_is_inf_6_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_is_inf_6_lpi_1_dfm,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_5_nl), alu_loop_op_6_FpMantRNE_49U_24U_else_and_1_tmp);
  assign nl_alu_loop_op_6_FpAdd_8U_23U_if_4_if_acc_2_nl = ({1'b1 , FpAdd_8U_23U_o_expo_6_lpi_1_dfm_2_7_4
      , (FpAdd_8U_23U_o_expo_6_lpi_1_dfm_2_3_0[3:1])}) + 8'b1;
  assign alu_loop_op_6_FpAdd_8U_23U_if_4_if_acc_2_nl = nl_alu_loop_op_6_FpAdd_8U_23U_if_4_if_acc_2_nl[7:0];
  assign alu_loop_op_6_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1 = readslicef_8_1_7((alu_loop_op_6_FpAdd_8U_23U_if_4_if_acc_2_nl));
  assign FpAdd_8U_23U_o_expo_6_lpi_1_dfm_2_7_4 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_6_lpi_1_dfm_1[7:4]),
      FpAdd_8U_23U_qr_7_lpi_1_dfm_5_7_4_1, (z_out_5[7:4]), {(~ (FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_276 , FpAdd_8U_23U_asn_278});
  assign FpAdd_8U_23U_is_inf_6_lpi_1_dfm = ~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_6_sva_2
      | (~ (FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_5[49])));
  assign FpAdd_8U_23U_and_37_tmp = alu_loop_op_6_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1
      & alu_loop_op_6_FpMantRNE_49U_24U_else_and_1_tmp;
  assign alu_loop_op_6_FpMantRNE_49U_24U_else_and_1_tmp = FpMantRNE_49U_24U_else_carry_6_sva
      & (FpAdd_8U_23U_int_mant_7_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign nl_FpAdd_8U_23U_o_expo_7_sva_4 = ({FpAdd_8U_23U_o_expo_7_lpi_1_dfm_2_7_4
      , FpAdd_8U_23U_o_expo_7_lpi_1_dfm_2_3_0}) + 8'b1;
  assign FpAdd_8U_23U_o_expo_7_sva_4 = nl_FpAdd_8U_23U_o_expo_7_sva_4[7:0];
  assign FpAdd_8U_23U_o_expo_7_lpi_1_dfm_1 = MUX_v_8_2_2(8'b00000000, z_out_6, FpNormalize_8U_49U_oelse_not_45);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_13_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      alu_loop_op_7_FpNormalize_8U_49U_else_lshift_itm, FpNormalize_8U_49U_oelse_not_45);
  assign FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_13_nl),
      (FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_5[49:1]), FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_5[49]);
  assign FpMantRNE_49U_24U_else_carry_7_sva = (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[25]));
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_6_nl = FpAdd_8U_23U_is_inf_7_lpi_1_dfm
      | (~ alu_loop_op_7_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1);
  assign FpAdd_8U_23U_is_inf_7_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_is_inf_7_lpi_1_dfm,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_6_nl), alu_loop_op_7_FpMantRNE_49U_24U_else_and_tmp);
  assign nl_alu_loop_op_7_FpAdd_8U_23U_if_4_if_acc_1_nl = ({1'b1 , FpAdd_8U_23U_o_expo_7_lpi_1_dfm_2_7_4
      , (FpAdd_8U_23U_o_expo_7_lpi_1_dfm_2_3_0[3:1])}) + 8'b1;
  assign alu_loop_op_7_FpAdd_8U_23U_if_4_if_acc_1_nl = nl_alu_loop_op_7_FpAdd_8U_23U_if_4_if_acc_1_nl[7:0];
  assign alu_loop_op_7_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1 = readslicef_8_1_7((alu_loop_op_7_FpAdd_8U_23U_if_4_if_acc_1_nl));
  assign FpAdd_8U_23U_o_expo_7_lpi_1_dfm_2_7_4 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_7_lpi_1_dfm_1[7:4]),
      FpAdd_8U_23U_qr_8_lpi_1_dfm_5_7_4_1, (z_out_6[7:4]), {(~ (FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_280 , FpAdd_8U_23U_asn_282});
  assign FpAdd_8U_23U_is_inf_7_lpi_1_dfm = ~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_7_sva_2
      | (~ (FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_5[49])));
  assign FpAdd_8U_23U_and_38_tmp = alu_loop_op_7_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1
      & alu_loop_op_7_FpMantRNE_49U_24U_else_and_tmp;
  assign alu_loop_op_7_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_else_carry_7_sva
      & (FpAdd_8U_23U_int_mant_8_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign nl_FpAdd_8U_23U_o_expo_8_sva_4 = ({FpAdd_8U_23U_o_expo_8_lpi_1_dfm_2_7_4
      , FpAdd_8U_23U_o_expo_8_lpi_1_dfm_2_3_0}) + 8'b1;
  assign FpAdd_8U_23U_o_expo_8_sva_4 = nl_FpAdd_8U_23U_o_expo_8_sva_4[7:0];
  assign FpAdd_8U_23U_o_expo_8_lpi_1_dfm_1 = MUX_v_8_2_2(8'b00000000, z_out_7, FpNormalize_8U_49U_oelse_not_47);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_15_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      alu_loop_op_8_FpNormalize_8U_49U_else_lshift_1_itm, FpNormalize_8U_49U_oelse_not_47);
  assign FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_15_nl),
      (FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_5[49:1]), FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_5[49]);
  assign FpMantRNE_49U_24U_else_carry_8_sva = (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[25]));
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_7_nl = FpAdd_8U_23U_is_inf_8_lpi_1_dfm
      | (~ alu_loop_op_8_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1);
  assign FpAdd_8U_23U_is_inf_8_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_is_inf_8_lpi_1_dfm,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_7_nl), alu_loop_op_8_FpMantRNE_49U_24U_else_and_1_tmp);
  assign nl_alu_loop_op_8_FpAdd_8U_23U_if_4_if_acc_2_nl = ({1'b1 , FpAdd_8U_23U_o_expo_8_lpi_1_dfm_2_7_4
      , (FpAdd_8U_23U_o_expo_8_lpi_1_dfm_2_3_0[3:1])}) + 8'b1;
  assign alu_loop_op_8_FpAdd_8U_23U_if_4_if_acc_2_nl = nl_alu_loop_op_8_FpAdd_8U_23U_if_4_if_acc_2_nl[7:0];
  assign alu_loop_op_8_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1 = readslicef_8_1_7((alu_loop_op_8_FpAdd_8U_23U_if_4_if_acc_2_nl));
  assign FpAdd_8U_23U_o_expo_8_lpi_1_dfm_2_7_4 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_8_lpi_1_dfm_1[7:4]),
      FpAdd_8U_23U_qr_9_lpi_1_dfm_5_7_4_1, (z_out_7[7:4]), {(~ (FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_284 , FpAdd_8U_23U_asn_286});
  assign FpAdd_8U_23U_is_inf_8_lpi_1_dfm = ~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_8_sva_2
      | (~ (FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_5[49])));
  assign FpAdd_8U_23U_and_39_tmp = alu_loop_op_8_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1
      & alu_loop_op_8_FpMantRNE_49U_24U_else_and_1_tmp;
  assign alu_loop_op_8_FpMantRNE_49U_24U_else_and_1_tmp = FpMantRNE_49U_24U_else_carry_8_sva
      & (FpAdd_8U_23U_int_mant_9_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign nl_FpAdd_8U_23U_o_expo_9_sva_4 = ({FpAdd_8U_23U_o_expo_9_lpi_1_dfm_2_7_4
      , FpAdd_8U_23U_o_expo_9_lpi_1_dfm_2_3_0}) + 8'b1;
  assign FpAdd_8U_23U_o_expo_9_sva_4 = nl_FpAdd_8U_23U_o_expo_9_sva_4[7:0];
  assign FpAdd_8U_23U_o_expo_9_lpi_1_dfm_1 = MUX_v_8_2_2(8'b00000000, z_out_8, FpNormalize_8U_49U_oelse_not_49);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_17_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      alu_loop_op_9_FpNormalize_8U_49U_else_lshift_itm, FpNormalize_8U_49U_oelse_not_49);
  assign FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_17_nl),
      (FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_5[49:1]), FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_5[49]);
  assign FpMantRNE_49U_24U_else_carry_9_sva = (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[25]));
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_8_nl = FpAdd_8U_23U_is_inf_9_lpi_1_dfm
      | (~ alu_loop_op_9_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1);
  assign FpAdd_8U_23U_is_inf_9_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_is_inf_9_lpi_1_dfm,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_8_nl), alu_loop_op_9_FpMantRNE_49U_24U_else_and_tmp);
  assign nl_alu_loop_op_9_FpAdd_8U_23U_if_4_if_acc_1_nl = ({1'b1 , FpAdd_8U_23U_o_expo_9_lpi_1_dfm_2_7_4
      , (FpAdd_8U_23U_o_expo_9_lpi_1_dfm_2_3_0[3:1])}) + 8'b1;
  assign alu_loop_op_9_FpAdd_8U_23U_if_4_if_acc_1_nl = nl_alu_loop_op_9_FpAdd_8U_23U_if_4_if_acc_1_nl[7:0];
  assign alu_loop_op_9_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1 = readslicef_8_1_7((alu_loop_op_9_FpAdd_8U_23U_if_4_if_acc_1_nl));
  assign FpAdd_8U_23U_o_expo_9_lpi_1_dfm_2_7_4 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_9_lpi_1_dfm_1[7:4]),
      FpAdd_8U_23U_qr_10_lpi_1_dfm_5_7_4_1, (z_out_8[7:4]), {(~ (FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_288 , FpAdd_8U_23U_asn_290});
  assign FpAdd_8U_23U_is_inf_9_lpi_1_dfm = ~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_9_sva_2
      | (~ (FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_5[49])));
  assign FpAdd_8U_23U_and_40_tmp = alu_loop_op_9_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1
      & alu_loop_op_9_FpMantRNE_49U_24U_else_and_tmp;
  assign alu_loop_op_9_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_else_carry_9_sva
      & (FpAdd_8U_23U_int_mant_10_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign nl_FpAdd_8U_23U_o_expo_10_sva_4 = ({FpAdd_8U_23U_o_expo_10_lpi_1_dfm_2_7_4
      , FpAdd_8U_23U_o_expo_10_lpi_1_dfm_2_3_0}) + 8'b1;
  assign FpAdd_8U_23U_o_expo_10_sva_4 = nl_FpAdd_8U_23U_o_expo_10_sva_4[7:0];
  assign FpAdd_8U_23U_o_expo_10_lpi_1_dfm_1 = MUX_v_8_2_2(8'b00000000, z_out_9, FpNormalize_8U_49U_oelse_not_51);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_19_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      alu_loop_op_10_FpNormalize_8U_49U_else_lshift_1_itm, FpNormalize_8U_49U_oelse_not_51);
  assign FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_19_nl),
      (FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_5[49:1]), FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_5[49]);
  assign FpMantRNE_49U_24U_else_carry_10_sva = (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[25]));
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_9_nl = FpAdd_8U_23U_is_inf_10_lpi_1_dfm
      | (~ alu_loop_op_10_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1);
  assign FpAdd_8U_23U_is_inf_10_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_is_inf_10_lpi_1_dfm,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_9_nl), alu_loop_op_10_FpMantRNE_49U_24U_else_and_1_tmp);
  assign nl_alu_loop_op_10_FpAdd_8U_23U_if_4_if_acc_2_nl = ({1'b1 , FpAdd_8U_23U_o_expo_10_lpi_1_dfm_2_7_4
      , (FpAdd_8U_23U_o_expo_10_lpi_1_dfm_2_3_0[3:1])}) + 8'b1;
  assign alu_loop_op_10_FpAdd_8U_23U_if_4_if_acc_2_nl = nl_alu_loop_op_10_FpAdd_8U_23U_if_4_if_acc_2_nl[7:0];
  assign alu_loop_op_10_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1 = readslicef_8_1_7((alu_loop_op_10_FpAdd_8U_23U_if_4_if_acc_2_nl));
  assign FpAdd_8U_23U_o_expo_10_lpi_1_dfm_2_7_4 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_10_lpi_1_dfm_1[7:4]),
      FpAdd_8U_23U_qr_11_lpi_1_dfm_5_7_4_1, (z_out_9[7:4]), {(~ (FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_292 , FpAdd_8U_23U_asn_294});
  assign FpAdd_8U_23U_is_inf_10_lpi_1_dfm = ~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_10_sva_2
      | (~ (FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_5[49])));
  assign FpAdd_8U_23U_and_41_tmp = alu_loop_op_10_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1
      & alu_loop_op_10_FpMantRNE_49U_24U_else_and_1_tmp;
  assign alu_loop_op_10_FpMantRNE_49U_24U_else_and_1_tmp = FpMantRNE_49U_24U_else_carry_10_sva
      & (FpAdd_8U_23U_int_mant_11_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign nl_FpAdd_8U_23U_o_expo_11_sva_4 = ({FpAdd_8U_23U_o_expo_11_lpi_1_dfm_2_7_4
      , FpAdd_8U_23U_o_expo_11_lpi_1_dfm_2_3_0}) + 8'b1;
  assign FpAdd_8U_23U_o_expo_11_sva_4 = nl_FpAdd_8U_23U_o_expo_11_sva_4[7:0];
  assign FpAdd_8U_23U_o_expo_11_lpi_1_dfm_1 = MUX_v_8_2_2(8'b00000000, z_out_10,
      FpNormalize_8U_49U_oelse_not_53);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_21_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      alu_loop_op_11_FpNormalize_8U_49U_else_lshift_itm, FpNormalize_8U_49U_oelse_not_53);
  assign FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_21_nl),
      (FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_5[49:1]), FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_5[49]);
  assign FpMantRNE_49U_24U_else_carry_11_sva = (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[25]));
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_10_nl = FpAdd_8U_23U_is_inf_11_lpi_1_dfm
      | (~ alu_loop_op_11_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1);
  assign FpAdd_8U_23U_is_inf_11_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_is_inf_11_lpi_1_dfm,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_10_nl), alu_loop_op_11_FpMantRNE_49U_24U_else_and_tmp);
  assign nl_alu_loop_op_11_FpAdd_8U_23U_if_4_if_acc_1_nl = ({1'b1 , FpAdd_8U_23U_o_expo_11_lpi_1_dfm_2_7_4
      , (FpAdd_8U_23U_o_expo_11_lpi_1_dfm_2_3_0[3:1])}) + 8'b1;
  assign alu_loop_op_11_FpAdd_8U_23U_if_4_if_acc_1_nl = nl_alu_loop_op_11_FpAdd_8U_23U_if_4_if_acc_1_nl[7:0];
  assign alu_loop_op_11_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1 = readslicef_8_1_7((alu_loop_op_11_FpAdd_8U_23U_if_4_if_acc_1_nl));
  assign FpAdd_8U_23U_o_expo_11_lpi_1_dfm_2_7_4 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_11_lpi_1_dfm_1[7:4]),
      FpAdd_8U_23U_qr_12_lpi_1_dfm_5_7_4_1, (z_out_10[7:4]), {(~ (FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_296 , FpAdd_8U_23U_asn_298});
  assign FpAdd_8U_23U_is_inf_11_lpi_1_dfm = ~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_11_sva_2
      | (~ (FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_5[49])));
  assign FpAdd_8U_23U_and_42_tmp = alu_loop_op_11_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1
      & alu_loop_op_11_FpMantRNE_49U_24U_else_and_tmp;
  assign alu_loop_op_11_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_else_carry_11_sva
      & (FpAdd_8U_23U_int_mant_12_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign nl_FpAdd_8U_23U_o_expo_12_sva_4 = ({FpAdd_8U_23U_o_expo_12_lpi_1_dfm_2_7_4
      , FpAdd_8U_23U_o_expo_12_lpi_1_dfm_2_3_0}) + 8'b1;
  assign FpAdd_8U_23U_o_expo_12_sva_4 = nl_FpAdd_8U_23U_o_expo_12_sva_4[7:0];
  assign FpAdd_8U_23U_o_expo_12_lpi_1_dfm_1 = MUX_v_8_2_2(8'b00000000, z_out_11,
      FpNormalize_8U_49U_oelse_not_55);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_23_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      alu_loop_op_12_FpNormalize_8U_49U_else_lshift_1_itm, FpNormalize_8U_49U_oelse_not_55);
  assign FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_23_nl),
      (FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_5[49:1]), FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_5[49]);
  assign FpMantRNE_49U_24U_else_carry_12_sva = (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[25]));
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_11_nl = FpAdd_8U_23U_is_inf_12_lpi_1_dfm
      | (~ alu_loop_op_12_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1);
  assign FpAdd_8U_23U_is_inf_12_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_is_inf_12_lpi_1_dfm,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_11_nl), alu_loop_op_12_FpMantRNE_49U_24U_else_and_1_tmp);
  assign nl_alu_loop_op_12_FpAdd_8U_23U_if_4_if_acc_2_nl = ({1'b1 , FpAdd_8U_23U_o_expo_12_lpi_1_dfm_2_7_4
      , (FpAdd_8U_23U_o_expo_12_lpi_1_dfm_2_3_0[3:1])}) + 8'b1;
  assign alu_loop_op_12_FpAdd_8U_23U_if_4_if_acc_2_nl = nl_alu_loop_op_12_FpAdd_8U_23U_if_4_if_acc_2_nl[7:0];
  assign alu_loop_op_12_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1 = readslicef_8_1_7((alu_loop_op_12_FpAdd_8U_23U_if_4_if_acc_2_nl));
  assign FpAdd_8U_23U_o_expo_12_lpi_1_dfm_2_7_4 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_12_lpi_1_dfm_1[7:4]),
      FpAdd_8U_23U_qr_13_lpi_1_dfm_5_7_4_1, (z_out_11[7:4]), {(~ (FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_300 , FpAdd_8U_23U_asn_302});
  assign FpAdd_8U_23U_is_inf_12_lpi_1_dfm = ~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_12_sva_2
      | (~ (FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_5[49])));
  assign FpAdd_8U_23U_and_43_tmp = alu_loop_op_12_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1
      & alu_loop_op_12_FpMantRNE_49U_24U_else_and_1_tmp;
  assign alu_loop_op_12_FpMantRNE_49U_24U_else_and_1_tmp = FpMantRNE_49U_24U_else_carry_12_sva
      & (FpAdd_8U_23U_int_mant_13_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign nl_FpAdd_8U_23U_o_expo_13_sva_4 = ({FpAdd_8U_23U_o_expo_13_lpi_1_dfm_2_7_4
      , FpAdd_8U_23U_o_expo_13_lpi_1_dfm_2_3_0}) + 8'b1;
  assign FpAdd_8U_23U_o_expo_13_sva_4 = nl_FpAdd_8U_23U_o_expo_13_sva_4[7:0];
  assign FpAdd_8U_23U_o_expo_13_lpi_1_dfm_1 = MUX_v_8_2_2(8'b00000000, z_out_12,
      FpNormalize_8U_49U_oelse_not_57);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_25_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      alu_loop_op_13_FpNormalize_8U_49U_else_lshift_itm, FpNormalize_8U_49U_oelse_not_57);
  assign FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_25_nl),
      (FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_5[49:1]), FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_5[49]);
  assign FpMantRNE_49U_24U_else_carry_13_sva = (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[25]));
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_12_nl = FpAdd_8U_23U_is_inf_13_lpi_1_dfm
      | (~ alu_loop_op_13_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1);
  assign FpAdd_8U_23U_is_inf_13_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_is_inf_13_lpi_1_dfm,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_12_nl), alu_loop_op_13_FpMantRNE_49U_24U_else_and_tmp);
  assign nl_alu_loop_op_13_FpAdd_8U_23U_if_4_if_acc_1_nl = ({1'b1 , FpAdd_8U_23U_o_expo_13_lpi_1_dfm_2_7_4
      , (FpAdd_8U_23U_o_expo_13_lpi_1_dfm_2_3_0[3:1])}) + 8'b1;
  assign alu_loop_op_13_FpAdd_8U_23U_if_4_if_acc_1_nl = nl_alu_loop_op_13_FpAdd_8U_23U_if_4_if_acc_1_nl[7:0];
  assign alu_loop_op_13_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1 = readslicef_8_1_7((alu_loop_op_13_FpAdd_8U_23U_if_4_if_acc_1_nl));
  assign FpAdd_8U_23U_o_expo_13_lpi_1_dfm_2_7_4 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_13_lpi_1_dfm_1[7:4]),
      FpAdd_8U_23U_qr_14_lpi_1_dfm_5_7_4_1, (z_out_12[7:4]), {(~ (FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_304 , FpAdd_8U_23U_asn_306});
  assign FpAdd_8U_23U_is_inf_13_lpi_1_dfm = ~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_13_sva_2
      | (~ (FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_5[49])));
  assign FpAdd_8U_23U_and_44_tmp = alu_loop_op_13_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1
      & alu_loop_op_13_FpMantRNE_49U_24U_else_and_tmp;
  assign alu_loop_op_13_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_else_carry_13_sva
      & (FpAdd_8U_23U_int_mant_14_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign nl_FpAdd_8U_23U_o_expo_14_sva_4 = ({FpAdd_8U_23U_o_expo_14_lpi_1_dfm_2_7_4
      , FpAdd_8U_23U_o_expo_14_lpi_1_dfm_2_3_0}) + 8'b1;
  assign FpAdd_8U_23U_o_expo_14_sva_4 = nl_FpAdd_8U_23U_o_expo_14_sva_4[7:0];
  assign FpAdd_8U_23U_o_expo_14_lpi_1_dfm_1 = MUX_v_8_2_2(8'b00000000, z_out_13,
      FpNormalize_8U_49U_oelse_not_59);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_27_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      alu_loop_op_14_FpNormalize_8U_49U_else_lshift_1_itm, FpNormalize_8U_49U_oelse_not_59);
  assign FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_27_nl),
      (FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_5[49:1]), FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_5[49]);
  assign FpMantRNE_49U_24U_else_carry_14_sva = (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[25]));
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_13_nl = FpAdd_8U_23U_is_inf_14_lpi_1_dfm
      | (~ alu_loop_op_14_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1);
  assign FpAdd_8U_23U_is_inf_14_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_is_inf_14_lpi_1_dfm,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_13_nl), alu_loop_op_14_FpMantRNE_49U_24U_else_and_1_tmp);
  assign nl_alu_loop_op_14_FpAdd_8U_23U_if_4_if_acc_2_nl = ({1'b1 , FpAdd_8U_23U_o_expo_14_lpi_1_dfm_2_7_4
      , (FpAdd_8U_23U_o_expo_14_lpi_1_dfm_2_3_0[3:1])}) + 8'b1;
  assign alu_loop_op_14_FpAdd_8U_23U_if_4_if_acc_2_nl = nl_alu_loop_op_14_FpAdd_8U_23U_if_4_if_acc_2_nl[7:0];
  assign alu_loop_op_14_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1 = readslicef_8_1_7((alu_loop_op_14_FpAdd_8U_23U_if_4_if_acc_2_nl));
  assign FpAdd_8U_23U_o_expo_14_lpi_1_dfm_2_7_4 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_14_lpi_1_dfm_1[7:4]),
      FpAdd_8U_23U_qr_15_lpi_1_dfm_5_7_4_1, (z_out_13[7:4]), {(~ (FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_308 , FpAdd_8U_23U_asn_310});
  assign FpAdd_8U_23U_is_inf_14_lpi_1_dfm = ~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_14_sva_2
      | (~ (FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_5[49])));
  assign FpAdd_8U_23U_and_45_tmp = alu_loop_op_14_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1
      & alu_loop_op_14_FpMantRNE_49U_24U_else_and_1_tmp;
  assign alu_loop_op_14_FpMantRNE_49U_24U_else_and_1_tmp = FpMantRNE_49U_24U_else_carry_14_sva
      & (FpAdd_8U_23U_int_mant_15_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign nl_FpAdd_8U_23U_o_expo_15_sva_4 = ({FpAdd_8U_23U_o_expo_15_lpi_1_dfm_2_7_4
      , FpAdd_8U_23U_o_expo_15_lpi_1_dfm_2_3_0}) + 8'b1;
  assign FpAdd_8U_23U_o_expo_15_sva_4 = nl_FpAdd_8U_23U_o_expo_15_sva_4[7:0];
  assign FpAdd_8U_23U_o_expo_15_lpi_1_dfm_1 = MUX_v_8_2_2(8'b00000000, z_out_14,
      FpNormalize_8U_49U_oelse_not_61);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_29_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      alu_loop_op_15_FpNormalize_8U_49U_else_lshift_itm, FpNormalize_8U_49U_oelse_not_61);
  assign FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_29_nl),
      (FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_5[49:1]), FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_5[49]);
  assign FpMantRNE_49U_24U_else_carry_15_sva = (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[25]));
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_14_nl = FpAdd_8U_23U_is_inf_15_lpi_1_dfm
      | (~ alu_loop_op_15_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1);
  assign FpAdd_8U_23U_is_inf_15_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_is_inf_15_lpi_1_dfm,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_14_nl), alu_loop_op_15_FpMantRNE_49U_24U_else_and_tmp);
  assign nl_alu_loop_op_15_FpAdd_8U_23U_if_4_if_acc_1_nl = ({1'b1 , FpAdd_8U_23U_o_expo_15_lpi_1_dfm_2_7_4
      , (FpAdd_8U_23U_o_expo_15_lpi_1_dfm_2_3_0[3:1])}) + 8'b1;
  assign alu_loop_op_15_FpAdd_8U_23U_if_4_if_acc_1_nl = nl_alu_loop_op_15_FpAdd_8U_23U_if_4_if_acc_1_nl[7:0];
  assign alu_loop_op_15_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1 = readslicef_8_1_7((alu_loop_op_15_FpAdd_8U_23U_if_4_if_acc_1_nl));
  assign FpAdd_8U_23U_o_expo_15_lpi_1_dfm_2_7_4 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_15_lpi_1_dfm_1[7:4]),
      FpAdd_8U_23U_qr_16_lpi_1_dfm_5_7_4_1, (z_out_14[7:4]), {(~ (FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_312 , FpAdd_8U_23U_asn_314});
  assign FpAdd_8U_23U_is_inf_15_lpi_1_dfm = ~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_15_sva_2
      | (~ (FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_5[49])));
  assign FpAdd_8U_23U_and_46_tmp = alu_loop_op_15_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1
      & alu_loop_op_15_FpMantRNE_49U_24U_else_and_tmp;
  assign alu_loop_op_15_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_else_carry_15_sva
      & (FpAdd_8U_23U_int_mant_16_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign nl_FpAdd_8U_23U_o_expo_sva_4 = ({FpAdd_8U_23U_o_expo_lpi_1_dfm_2_7_4 , FpAdd_8U_23U_o_expo_lpi_1_dfm_2_3_0})
      + 8'b1;
  assign FpAdd_8U_23U_o_expo_sva_4 = nl_FpAdd_8U_23U_o_expo_sva_4[7:0];
  assign FpAdd_8U_23U_o_expo_lpi_1_dfm_1 = MUX_v_8_2_2(8'b00000000, z_out_15, FpNormalize_8U_49U_oelse_not_63);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_31_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      alu_loop_op_16_FpNormalize_8U_49U_else_lshift_1_itm, FpNormalize_8U_49U_oelse_not_63);
  assign FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_31_nl),
      (FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49:1]), FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49]);
  assign FpMantRNE_49U_24U_else_carry_sva = (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[25]));
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_15_nl = FpAdd_8U_23U_is_inf_lpi_1_dfm
      | (~ alu_loop_op_16_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1);
  assign FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_is_inf_lpi_1_dfm,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_15_nl), alu_loop_op_16_FpMantRNE_49U_24U_else_and_1_tmp);
  assign nl_alu_loop_op_16_FpAdd_8U_23U_if_4_if_acc_2_nl = ({1'b1 , FpAdd_8U_23U_o_expo_lpi_1_dfm_2_7_4
      , (FpAdd_8U_23U_o_expo_lpi_1_dfm_2_3_0[3:1])}) + 8'b1;
  assign alu_loop_op_16_FpAdd_8U_23U_if_4_if_acc_2_nl = nl_alu_loop_op_16_FpAdd_8U_23U_if_4_if_acc_2_nl[7:0];
  assign alu_loop_op_16_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1 = readslicef_8_1_7((alu_loop_op_16_FpAdd_8U_23U_if_4_if_acc_2_nl));
  assign FpAdd_8U_23U_o_expo_lpi_1_dfm_2_7_4 = MUX1HOT_v_4_3_2((FpAdd_8U_23U_o_expo_lpi_1_dfm_1[7:4]),
      FpAdd_8U_23U_qr_lpi_1_dfm_5_7_4_1, (z_out_15[7:4]), {(~ (FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49]))
      , FpAdd_8U_23U_asn_316 , FpAdd_8U_23U_asn_318});
  assign FpAdd_8U_23U_is_inf_lpi_1_dfm = ~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_2
      | (~ (FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49])));
  assign FpAdd_8U_23U_and_47_tmp = alu_loop_op_16_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1
      & alu_loop_op_16_FpMantRNE_49U_24U_else_and_1_tmp;
  assign alu_loop_op_16_FpMantRNE_49U_24U_else_and_1_tmp = FpMantRNE_49U_24U_else_carry_sva
      & (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign nor_7_ssc = ~(else_unequal_tmp | io_read_cfg_alu_bypass_rsc_svs_7);
  assign and_1_m1c = else_unequal_tmp & (~ io_read_cfg_alu_bypass_rsc_svs_7);
  assign alu_nan_to_zero_aelse_not_111_nl = ~ alu_nan_to_zero_land_1_lpi_1_dfm;
  assign alu_nan_to_zero_op_expo_1_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_AluOp_data_0_14_10_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_111_nl));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_1_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_16)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_1_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_1_sva[5:0];
  assign alu_nan_to_zero_aelse_not_95_nl = ~ alu_nan_to_zero_land_1_lpi_1_dfm;
  assign alu_nan_to_zero_op_mant_1_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_AluOp_data_0_9_0_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_95_nl));
  assign alu_nan_to_zero_aelse_not_110_nl = ~ alu_nan_to_zero_land_2_lpi_1_dfm;
  assign alu_nan_to_zero_op_expo_2_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_AluOp_data_1_14_10_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_110_nl));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_2_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_17)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_2_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_2_sva[5:0];
  assign alu_nan_to_zero_aelse_not_94_nl = ~ alu_nan_to_zero_land_2_lpi_1_dfm;
  assign alu_nan_to_zero_op_mant_2_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_AluOp_data_1_9_0_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_94_nl));
  assign alu_nan_to_zero_aelse_not_109_nl = ~ alu_nan_to_zero_land_3_lpi_1_dfm;
  assign alu_nan_to_zero_op_expo_3_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_AluOp_data_2_14_10_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_109_nl));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_3_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_18)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_3_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_3_sva[5:0];
  assign alu_nan_to_zero_aelse_not_93_nl = ~ alu_nan_to_zero_land_3_lpi_1_dfm;
  assign alu_nan_to_zero_op_mant_3_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_AluOp_data_2_9_0_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_93_nl));
  assign alu_nan_to_zero_aelse_not_108_nl = ~ alu_nan_to_zero_land_4_lpi_1_dfm;
  assign alu_nan_to_zero_op_expo_4_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_AluOp_data_3_14_10_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_108_nl));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_4_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_19)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_4_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_4_sva[5:0];
  assign alu_nan_to_zero_aelse_not_92_nl = ~ alu_nan_to_zero_land_4_lpi_1_dfm;
  assign alu_nan_to_zero_op_mant_4_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_AluOp_data_3_9_0_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_92_nl));
  assign alu_nan_to_zero_aelse_not_107_nl = ~ alu_nan_to_zero_land_5_lpi_1_dfm;
  assign alu_nan_to_zero_op_expo_5_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_AluOp_data_4_14_10_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_107_nl));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_5_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_20)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_5_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_5_sva[5:0];
  assign alu_nan_to_zero_aelse_not_91_nl = ~ alu_nan_to_zero_land_5_lpi_1_dfm;
  assign alu_nan_to_zero_op_mant_5_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_AluOp_data_4_9_0_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_91_nl));
  assign alu_nan_to_zero_aelse_not_106_nl = ~ alu_nan_to_zero_land_6_lpi_1_dfm;
  assign alu_nan_to_zero_op_expo_6_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_AluOp_data_5_14_10_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_106_nl));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_6_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_21)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_6_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_6_sva[5:0];
  assign alu_nan_to_zero_aelse_not_90_nl = ~ alu_nan_to_zero_land_6_lpi_1_dfm;
  assign alu_nan_to_zero_op_mant_6_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_AluOp_data_5_9_0_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_90_nl));
  assign alu_nan_to_zero_aelse_not_105_nl = ~ alu_nan_to_zero_land_7_lpi_1_dfm;
  assign alu_nan_to_zero_op_expo_7_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_AluOp_data_6_14_10_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_105_nl));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_7_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_22)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_7_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_7_sva[5:0];
  assign alu_nan_to_zero_aelse_not_89_nl = ~ alu_nan_to_zero_land_7_lpi_1_dfm;
  assign alu_nan_to_zero_op_mant_7_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_AluOp_data_6_9_0_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_89_nl));
  assign alu_nan_to_zero_aelse_not_104_nl = ~ alu_nan_to_zero_land_8_lpi_1_dfm;
  assign alu_nan_to_zero_op_expo_8_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_AluOp_data_7_14_10_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_104_nl));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_8_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_23)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_8_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_8_sva[5:0];
  assign alu_nan_to_zero_aelse_not_88_nl = ~ alu_nan_to_zero_land_8_lpi_1_dfm;
  assign alu_nan_to_zero_op_mant_8_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_AluOp_data_7_9_0_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_88_nl));
  assign alu_nan_to_zero_aelse_not_103_nl = ~ alu_nan_to_zero_land_9_lpi_1_dfm;
  assign alu_nan_to_zero_op_expo_9_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_AluOp_data_8_14_10_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_103_nl));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_9_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_24)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_9_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_9_sva[5:0];
  assign alu_nan_to_zero_aelse_not_87_nl = ~ alu_nan_to_zero_land_9_lpi_1_dfm;
  assign alu_nan_to_zero_op_mant_9_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_AluOp_data_8_9_0_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_87_nl));
  assign alu_nan_to_zero_aelse_not_102_nl = ~ alu_nan_to_zero_land_10_lpi_1_dfm;
  assign alu_nan_to_zero_op_expo_10_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_AluOp_data_9_14_10_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_102_nl));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_10_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_25)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_10_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_10_sva[5:0];
  assign alu_nan_to_zero_aelse_not_86_nl = ~ alu_nan_to_zero_land_10_lpi_1_dfm;
  assign alu_nan_to_zero_op_mant_10_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_AluOp_data_9_9_0_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_86_nl));
  assign alu_nan_to_zero_aelse_not_101_nl = ~ alu_nan_to_zero_land_11_lpi_1_dfm;
  assign alu_nan_to_zero_op_expo_11_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_AluOp_data_10_14_10_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_101_nl));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_11_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_26)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_11_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_11_sva[5:0];
  assign alu_nan_to_zero_aelse_not_85_nl = ~ alu_nan_to_zero_land_11_lpi_1_dfm;
  assign alu_nan_to_zero_op_mant_11_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_AluOp_data_10_9_0_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_85_nl));
  assign alu_nan_to_zero_aelse_not_100_nl = ~ alu_nan_to_zero_land_12_lpi_1_dfm;
  assign alu_nan_to_zero_op_expo_12_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_AluOp_data_11_14_10_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_100_nl));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_12_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_27)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_12_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_12_sva[5:0];
  assign alu_nan_to_zero_aelse_not_84_nl = ~ alu_nan_to_zero_land_12_lpi_1_dfm;
  assign alu_nan_to_zero_op_mant_12_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_AluOp_data_11_9_0_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_84_nl));
  assign alu_nan_to_zero_aelse_not_99_nl = ~ alu_nan_to_zero_land_13_lpi_1_dfm;
  assign alu_nan_to_zero_op_expo_13_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_AluOp_data_12_14_10_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_99_nl));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_13_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_28)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_13_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_13_sva[5:0];
  assign alu_nan_to_zero_aelse_not_83_nl = ~ alu_nan_to_zero_land_13_lpi_1_dfm;
  assign alu_nan_to_zero_op_mant_13_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_AluOp_data_12_9_0_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_83_nl));
  assign alu_nan_to_zero_aelse_not_98_nl = ~ alu_nan_to_zero_land_14_lpi_1_dfm;
  assign alu_nan_to_zero_op_expo_14_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_AluOp_data_13_14_10_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_98_nl));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_14_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_29)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_14_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_14_sva[5:0];
  assign alu_nan_to_zero_aelse_not_82_nl = ~ alu_nan_to_zero_land_14_lpi_1_dfm;
  assign alu_nan_to_zero_op_mant_14_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_AluOp_data_13_9_0_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_82_nl));
  assign alu_nan_to_zero_aelse_not_97_nl = ~ alu_nan_to_zero_land_15_lpi_1_dfm;
  assign alu_nan_to_zero_op_expo_15_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_AluOp_data_14_14_10_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_97_nl));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_15_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_30)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_15_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_15_sva[5:0];
  assign alu_nan_to_zero_aelse_not_81_nl = ~ alu_nan_to_zero_land_15_lpi_1_dfm;
  assign alu_nan_to_zero_op_mant_15_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_AluOp_data_14_9_0_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_81_nl));
  assign alu_nan_to_zero_aelse_not_96_nl = ~ alu_nan_to_zero_land_lpi_1_dfm;
  assign alu_nan_to_zero_op_expo_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_AluOp_data_15_14_10_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_96_nl));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_31)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_sva[5:0];
  assign alu_nan_to_zero_aelse_not_80_nl = ~ alu_nan_to_zero_land_lpi_1_dfm;
  assign alu_nan_to_zero_op_mant_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_AluOp_data_15_9_0_lpi_1_dfm_mx0,
      (alu_nan_to_zero_aelse_not_80_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_30_ssc
      = ~(IsDenorm_5U_23U_land_lpi_1_dfm | IsInf_5U_23U_land_lpi_1_dfm);
  assign IsDenorm_5U_23U_land_lpi_1_dfm = ((alu_nan_to_zero_op_mant_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_sva;
  assign IsInf_5U_23U_land_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_lpi_1_dfm!=10'b0000000000) |
      IsNaN_5U_23U_IsNaN_5U_23U_nand_15_cse);
  assign IsNaN_5U_23U_nor_15_tmp = ~((alu_nan_to_zero_op_mant_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_lpi_1_dfm = ~(IsNaN_5U_23U_nor_15_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_15_cse);
  assign IsNaN_5U_23U_aelse_not_47_nl = ~ IsNaN_5U_23U_land_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_47_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_lpi_1_dfm, IsNaN_5U_23U_land_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_15_cse = ~((alu_nan_to_zero_op_expo_lpi_1_dfm==5'b11111));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_sva = ~((alu_nan_to_zero_op_expo_lpi_1_dfm!=5'b00000));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_28_ssc
      = ~(IsDenorm_5U_23U_land_15_lpi_1_dfm | IsInf_5U_23U_land_15_lpi_1_dfm);
  assign IsDenorm_5U_23U_land_15_lpi_1_dfm = ((alu_nan_to_zero_op_mant_15_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_15_sva;
  assign IsInf_5U_23U_land_15_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_15_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_15_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_14_cse);
  assign IsNaN_5U_23U_nor_14_tmp = ~((alu_nan_to_zero_op_mant_15_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_15_lpi_1_dfm = ~(IsNaN_5U_23U_nor_14_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_14_cse);
  assign IsNaN_5U_23U_aelse_not_46_nl = ~ IsNaN_5U_23U_land_15_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_15_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_15_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_46_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_15_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_15_lpi_1_dfm, IsNaN_5U_23U_land_15_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_14_cse = ~((alu_nan_to_zero_op_expo_15_lpi_1_dfm==5'b11111));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_15_sva = ~((alu_nan_to_zero_op_expo_15_lpi_1_dfm!=5'b00000));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_26_ssc
      = ~(IsDenorm_5U_23U_land_14_lpi_1_dfm | IsInf_5U_23U_land_14_lpi_1_dfm);
  assign IsDenorm_5U_23U_land_14_lpi_1_dfm = ((alu_nan_to_zero_op_mant_14_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_14_sva;
  assign IsInf_5U_23U_land_14_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_14_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_14_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_13_cse);
  assign IsNaN_5U_23U_nor_13_tmp = ~((alu_nan_to_zero_op_mant_14_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_14_lpi_1_dfm = ~(IsNaN_5U_23U_nor_13_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_13_cse);
  assign IsNaN_5U_23U_aelse_not_45_nl = ~ IsNaN_5U_23U_land_14_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_14_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_14_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_45_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_14_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_14_lpi_1_dfm, IsNaN_5U_23U_land_14_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_13_cse = ~((alu_nan_to_zero_op_expo_14_lpi_1_dfm==5'b11111));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_14_sva = ~((alu_nan_to_zero_op_expo_14_lpi_1_dfm!=5'b00000));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_24_ssc
      = ~(IsDenorm_5U_23U_land_13_lpi_1_dfm | IsInf_5U_23U_land_13_lpi_1_dfm);
  assign IsDenorm_5U_23U_land_13_lpi_1_dfm = ((alu_nan_to_zero_op_mant_13_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_13_sva;
  assign IsInf_5U_23U_land_13_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_13_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_13_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_12_cse);
  assign IsNaN_5U_23U_nor_12_tmp = ~((alu_nan_to_zero_op_mant_13_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_13_lpi_1_dfm = ~(IsNaN_5U_23U_nor_12_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_12_cse);
  assign IsNaN_5U_23U_aelse_not_44_nl = ~ IsNaN_5U_23U_land_13_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_13_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_13_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_44_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_13_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_13_lpi_1_dfm, IsNaN_5U_23U_land_13_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_12_cse = ~((alu_nan_to_zero_op_expo_13_lpi_1_dfm==5'b11111));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_13_sva = ~((alu_nan_to_zero_op_expo_13_lpi_1_dfm!=5'b00000));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_22_ssc
      = ~(IsDenorm_5U_23U_land_12_lpi_1_dfm | IsInf_5U_23U_land_12_lpi_1_dfm);
  assign IsDenorm_5U_23U_land_12_lpi_1_dfm = ((alu_nan_to_zero_op_mant_12_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_12_sva;
  assign IsInf_5U_23U_land_12_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_12_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_12_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_11_cse);
  assign IsNaN_5U_23U_nor_11_tmp = ~((alu_nan_to_zero_op_mant_12_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_12_lpi_1_dfm = ~(IsNaN_5U_23U_nor_11_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_11_cse);
  assign IsNaN_5U_23U_aelse_not_43_nl = ~ IsNaN_5U_23U_land_12_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_12_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_12_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_43_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_12_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_12_lpi_1_dfm, IsNaN_5U_23U_land_12_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_11_cse = ~((alu_nan_to_zero_op_expo_12_lpi_1_dfm==5'b11111));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_12_sva = ~((alu_nan_to_zero_op_expo_12_lpi_1_dfm!=5'b00000));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_20_ssc
      = ~(IsDenorm_5U_23U_land_11_lpi_1_dfm | IsInf_5U_23U_land_11_lpi_1_dfm);
  assign IsDenorm_5U_23U_land_11_lpi_1_dfm = ((alu_nan_to_zero_op_mant_11_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_11_sva;
  assign IsInf_5U_23U_land_11_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_11_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_11_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_10_cse);
  assign IsNaN_5U_23U_nor_10_tmp = ~((alu_nan_to_zero_op_mant_11_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_11_lpi_1_dfm = ~(IsNaN_5U_23U_nor_10_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_10_cse);
  assign IsNaN_5U_23U_aelse_not_42_nl = ~ IsNaN_5U_23U_land_11_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_11_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_11_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_42_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_11_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_11_lpi_1_dfm, IsNaN_5U_23U_land_11_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_10_cse = ~((alu_nan_to_zero_op_expo_11_lpi_1_dfm==5'b11111));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_11_sva = ~((alu_nan_to_zero_op_expo_11_lpi_1_dfm!=5'b00000));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_18_ssc
      = ~(IsDenorm_5U_23U_land_10_lpi_1_dfm | IsInf_5U_23U_land_10_lpi_1_dfm);
  assign IsDenorm_5U_23U_land_10_lpi_1_dfm = ((alu_nan_to_zero_op_mant_10_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_10_sva;
  assign IsInf_5U_23U_land_10_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_10_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_10_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_9_cse);
  assign IsNaN_5U_23U_nor_9_tmp = ~((alu_nan_to_zero_op_mant_10_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_10_lpi_1_dfm = ~(IsNaN_5U_23U_nor_9_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_9_cse);
  assign IsNaN_5U_23U_aelse_not_41_nl = ~ IsNaN_5U_23U_land_10_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_10_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_10_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_41_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_10_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_10_lpi_1_dfm, IsNaN_5U_23U_land_10_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_9_cse = ~((alu_nan_to_zero_op_expo_10_lpi_1_dfm==5'b11111));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_10_sva = ~((alu_nan_to_zero_op_expo_10_lpi_1_dfm!=5'b00000));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_16_ssc
      = ~(IsDenorm_5U_23U_land_9_lpi_1_dfm | IsInf_5U_23U_land_9_lpi_1_dfm);
  assign IsDenorm_5U_23U_land_9_lpi_1_dfm = ((alu_nan_to_zero_op_mant_9_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_9_sva;
  assign IsInf_5U_23U_land_9_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_9_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_9_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_8_cse);
  assign IsNaN_5U_23U_nor_8_tmp = ~((alu_nan_to_zero_op_mant_9_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_9_lpi_1_dfm = ~(IsNaN_5U_23U_nor_8_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_8_cse);
  assign IsNaN_5U_23U_aelse_not_40_nl = ~ IsNaN_5U_23U_land_9_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_9_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_9_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_40_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_9_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_9_lpi_1_dfm, IsNaN_5U_23U_land_9_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_8_cse = ~((alu_nan_to_zero_op_expo_9_lpi_1_dfm==5'b11111));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_9_sva = ~((alu_nan_to_zero_op_expo_9_lpi_1_dfm!=5'b00000));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_ssc
      = ~(IsDenorm_5U_23U_land_8_lpi_1_dfm | IsInf_5U_23U_land_8_lpi_1_dfm);
  assign IsDenorm_5U_23U_land_8_lpi_1_dfm = ((alu_nan_to_zero_op_mant_8_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_8_sva;
  assign IsInf_5U_23U_land_8_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_8_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_8_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_7_cse);
  assign IsNaN_5U_23U_nor_7_tmp = ~((alu_nan_to_zero_op_mant_8_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_8_lpi_1_dfm = ~(IsNaN_5U_23U_nor_7_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_7_cse);
  assign IsNaN_5U_23U_aelse_not_39_nl = ~ IsNaN_5U_23U_land_8_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_8_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_8_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_39_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_8_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_8_lpi_1_dfm, IsNaN_5U_23U_land_8_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_7_cse = ~((alu_nan_to_zero_op_expo_8_lpi_1_dfm==5'b11111));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_8_sva = ~((alu_nan_to_zero_op_expo_8_lpi_1_dfm!=5'b00000));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_ssc
      = ~(IsDenorm_5U_23U_land_7_lpi_1_dfm | IsInf_5U_23U_land_7_lpi_1_dfm);
  assign IsDenorm_5U_23U_land_7_lpi_1_dfm = ((alu_nan_to_zero_op_mant_7_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_7_sva;
  assign IsInf_5U_23U_land_7_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_7_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_7_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_6_cse);
  assign IsNaN_5U_23U_nor_6_tmp = ~((alu_nan_to_zero_op_mant_7_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_7_lpi_1_dfm = ~(IsNaN_5U_23U_nor_6_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_6_cse);
  assign IsNaN_5U_23U_aelse_not_38_nl = ~ IsNaN_5U_23U_land_7_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_7_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_7_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_38_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_7_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_7_lpi_1_dfm, IsNaN_5U_23U_land_7_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_6_cse = ~((alu_nan_to_zero_op_expo_7_lpi_1_dfm==5'b11111));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_7_sva = ~((alu_nan_to_zero_op_expo_7_lpi_1_dfm!=5'b00000));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_ssc
      = ~(IsDenorm_5U_23U_land_6_lpi_1_dfm | IsInf_5U_23U_land_6_lpi_1_dfm);
  assign IsDenorm_5U_23U_land_6_lpi_1_dfm = ((alu_nan_to_zero_op_mant_6_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_6_sva;
  assign IsInf_5U_23U_land_6_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_6_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_6_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_5_cse);
  assign IsNaN_5U_23U_nor_5_tmp = ~((alu_nan_to_zero_op_mant_6_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_6_lpi_1_dfm = ~(IsNaN_5U_23U_nor_5_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_5_cse);
  assign IsNaN_5U_23U_aelse_not_37_nl = ~ IsNaN_5U_23U_land_6_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_6_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_6_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_37_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_6_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_6_lpi_1_dfm, IsNaN_5U_23U_land_6_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_5_cse = ~((alu_nan_to_zero_op_expo_6_lpi_1_dfm==5'b11111));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_6_sva = ~((alu_nan_to_zero_op_expo_6_lpi_1_dfm!=5'b00000));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_ssc
      = ~(IsDenorm_5U_23U_land_5_lpi_1_dfm | IsInf_5U_23U_land_5_lpi_1_dfm);
  assign IsDenorm_5U_23U_land_5_lpi_1_dfm = ((alu_nan_to_zero_op_mant_5_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_5_sva;
  assign IsInf_5U_23U_land_5_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_5_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_5_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_4_cse);
  assign IsNaN_5U_23U_nor_4_tmp = ~((alu_nan_to_zero_op_mant_5_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_5_lpi_1_dfm = ~(IsNaN_5U_23U_nor_4_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_4_cse);
  assign IsNaN_5U_23U_aelse_not_36_nl = ~ IsNaN_5U_23U_land_5_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_5_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_5_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_36_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_5_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_5_lpi_1_dfm, IsNaN_5U_23U_land_5_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_4_cse = ~((alu_nan_to_zero_op_expo_5_lpi_1_dfm==5'b11111));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_5_sva = ~((alu_nan_to_zero_op_expo_5_lpi_1_dfm!=5'b00000));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_ssc
      = ~(IsDenorm_5U_23U_land_4_lpi_1_dfm | IsInf_5U_23U_land_4_lpi_1_dfm);
  assign IsDenorm_5U_23U_land_4_lpi_1_dfm = ((alu_nan_to_zero_op_mant_4_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_4_sva;
  assign IsInf_5U_23U_land_4_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_4_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_4_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_3_cse);
  assign IsNaN_5U_23U_nor_3_tmp = ~((alu_nan_to_zero_op_mant_4_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_4_lpi_1_dfm = ~(IsNaN_5U_23U_nor_3_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_3_cse);
  assign IsNaN_5U_23U_aelse_not_35_nl = ~ IsNaN_5U_23U_land_4_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_4_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_4_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_35_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_4_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_4_lpi_1_dfm, IsNaN_5U_23U_land_4_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_3_cse = ~((alu_nan_to_zero_op_expo_4_lpi_1_dfm==5'b11111));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_4_sva = ~((alu_nan_to_zero_op_expo_4_lpi_1_dfm!=5'b00000));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_ssc
      = ~(IsDenorm_5U_23U_land_3_lpi_1_dfm | IsInf_5U_23U_land_3_lpi_1_dfm);
  assign IsDenorm_5U_23U_land_3_lpi_1_dfm = ((alu_nan_to_zero_op_mant_3_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_3_sva;
  assign IsInf_5U_23U_land_3_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_3_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_3_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_2_cse);
  assign IsNaN_5U_23U_nor_2_tmp = ~((alu_nan_to_zero_op_mant_3_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_3_lpi_1_dfm = ~(IsNaN_5U_23U_nor_2_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_2_cse);
  assign IsNaN_5U_23U_aelse_not_34_nl = ~ IsNaN_5U_23U_land_3_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_3_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_3_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_34_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_3_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_3_lpi_1_dfm, IsNaN_5U_23U_land_3_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_2_cse = ~((alu_nan_to_zero_op_expo_3_lpi_1_dfm==5'b11111));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_3_sva = ~((alu_nan_to_zero_op_expo_3_lpi_1_dfm!=5'b00000));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_ssc
      = ~(IsDenorm_5U_23U_land_2_lpi_1_dfm | IsInf_5U_23U_land_2_lpi_1_dfm);
  assign IsDenorm_5U_23U_land_2_lpi_1_dfm = ((alu_nan_to_zero_op_mant_2_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_2_sva;
  assign IsInf_5U_23U_land_2_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_2_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_2_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_1_cse);
  assign IsNaN_5U_23U_nor_1_tmp = ~((alu_nan_to_zero_op_mant_2_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_2_lpi_1_dfm = ~(IsNaN_5U_23U_nor_1_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_1_cse);
  assign IsNaN_5U_23U_aelse_not_33_nl = ~ IsNaN_5U_23U_land_2_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_2_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_2_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_33_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_2_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_2_lpi_1_dfm, IsNaN_5U_23U_land_2_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_1_cse = ~((alu_nan_to_zero_op_expo_2_lpi_1_dfm==5'b11111));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_2_sva = ~((alu_nan_to_zero_op_expo_2_lpi_1_dfm!=5'b00000));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_ssc =
      ~(IsDenorm_5U_23U_land_1_lpi_1_dfm | IsInf_5U_23U_land_1_lpi_1_dfm);
  assign IsDenorm_5U_23U_land_1_lpi_1_dfm = ((alu_nan_to_zero_op_mant_1_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_1_sva;
  assign IsInf_5U_23U_land_1_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_1_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_1_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_cse);
  assign IsNaN_5U_23U_nor_tmp = ~((alu_nan_to_zero_op_mant_1_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_1_lpi_1_dfm = ~(IsNaN_5U_23U_nor_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_cse);
  assign IsNaN_5U_23U_aelse_not_32_nl = ~ IsNaN_5U_23U_land_1_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_1_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_1_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_32_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_1_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      alu_nan_to_zero_op_mant_1_lpi_1_dfm, IsNaN_5U_23U_land_1_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_cse = ~((alu_nan_to_zero_op_expo_1_lpi_1_dfm==5'b11111));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_1_sva = ~((alu_nan_to_zero_op_expo_1_lpi_1_dfm!=5'b00000));
  assign else_AluOp_data_15_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]),
      (chn_alu_op_rsci_d_mxwt[254:250]), cfg_alu_src_1_sva_st);
  assign IsNaN_5U_10U_nor_15_tmp = ~((else_AluOp_data_15_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign alu_nan_to_zero_land_lpi_1_dfm = (~(IsNaN_5U_10U_nor_15_tmp | (else_AluOp_data_15_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_AluOp_data_15_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_alu_op_1_sva_1[9:0]),
      (chn_alu_op_rsci_d_mxwt[249:240]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_14_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]),
      (chn_alu_op_rsci_d_mxwt[238:234]), cfg_alu_src_1_sva_st);
  assign IsNaN_5U_10U_nor_14_tmp = ~((else_AluOp_data_14_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign alu_nan_to_zero_land_15_lpi_1_dfm = (~(IsNaN_5U_10U_nor_14_tmp | (else_AluOp_data_14_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_AluOp_data_14_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_alu_op_1_sva_1[9:0]),
      (chn_alu_op_rsci_d_mxwt[233:224]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_13_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]),
      (chn_alu_op_rsci_d_mxwt[222:218]), cfg_alu_src_1_sva_st);
  assign IsNaN_5U_10U_nor_13_tmp = ~((else_AluOp_data_13_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign alu_nan_to_zero_land_14_lpi_1_dfm = (~(IsNaN_5U_10U_nor_13_tmp | (else_AluOp_data_13_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_AluOp_data_13_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_alu_op_1_sva_1[9:0]),
      (chn_alu_op_rsci_d_mxwt[217:208]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_12_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]),
      (chn_alu_op_rsci_d_mxwt[206:202]), cfg_alu_src_1_sva_st);
  assign IsNaN_5U_10U_nor_12_tmp = ~((else_AluOp_data_12_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign alu_nan_to_zero_land_13_lpi_1_dfm = (~(IsNaN_5U_10U_nor_12_tmp | (else_AluOp_data_12_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_AluOp_data_12_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_alu_op_1_sva_1[9:0]),
      (chn_alu_op_rsci_d_mxwt[201:192]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_11_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]),
      (chn_alu_op_rsci_d_mxwt[190:186]), cfg_alu_src_1_sva_st);
  assign IsNaN_5U_10U_nor_11_tmp = ~((else_AluOp_data_11_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign alu_nan_to_zero_land_12_lpi_1_dfm = (~(IsNaN_5U_10U_nor_11_tmp | (else_AluOp_data_11_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_AluOp_data_11_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_alu_op_1_sva_1[9:0]),
      (chn_alu_op_rsci_d_mxwt[185:176]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_10_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]),
      (chn_alu_op_rsci_d_mxwt[174:170]), cfg_alu_src_1_sva_st);
  assign IsNaN_5U_10U_nor_10_tmp = ~((else_AluOp_data_10_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign alu_nan_to_zero_land_11_lpi_1_dfm = (~(IsNaN_5U_10U_nor_10_tmp | (else_AluOp_data_10_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_AluOp_data_10_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_alu_op_1_sva_1[9:0]),
      (chn_alu_op_rsci_d_mxwt[169:160]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_9_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]),
      (chn_alu_op_rsci_d_mxwt[158:154]), cfg_alu_src_1_sva_st);
  assign IsNaN_5U_10U_nor_9_tmp = ~((else_AluOp_data_9_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign alu_nan_to_zero_land_10_lpi_1_dfm = (~(IsNaN_5U_10U_nor_9_tmp | (else_AluOp_data_9_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_AluOp_data_9_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_alu_op_1_sva_1[9:0]),
      (chn_alu_op_rsci_d_mxwt[153:144]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_8_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]),
      (chn_alu_op_rsci_d_mxwt[142:138]), cfg_alu_src_1_sva_st);
  assign IsNaN_5U_10U_nor_8_tmp = ~((else_AluOp_data_8_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign alu_nan_to_zero_land_9_lpi_1_dfm = (~(IsNaN_5U_10U_nor_8_tmp | (else_AluOp_data_8_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_AluOp_data_8_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_alu_op_1_sva_1[9:0]),
      (chn_alu_op_rsci_d_mxwt[137:128]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_7_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]),
      (chn_alu_op_rsci_d_mxwt[126:122]), cfg_alu_src_1_sva_st);
  assign IsNaN_5U_10U_nor_7_tmp = ~((else_AluOp_data_7_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign alu_nan_to_zero_land_8_lpi_1_dfm = (~(IsNaN_5U_10U_nor_7_tmp | (else_AluOp_data_7_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_AluOp_data_7_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_alu_op_1_sva_1[9:0]),
      (chn_alu_op_rsci_d_mxwt[121:112]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_6_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]),
      (chn_alu_op_rsci_d_mxwt[110:106]), cfg_alu_src_1_sva_st);
  assign IsNaN_5U_10U_nor_6_tmp = ~((else_AluOp_data_6_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign alu_nan_to_zero_land_7_lpi_1_dfm = (~(IsNaN_5U_10U_nor_6_tmp | (else_AluOp_data_6_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_AluOp_data_6_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_alu_op_1_sva_1[9:0]),
      (chn_alu_op_rsci_d_mxwt[105:96]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_5_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]),
      (chn_alu_op_rsci_d_mxwt[94:90]), cfg_alu_src_1_sva_st);
  assign IsNaN_5U_10U_nor_5_tmp = ~((else_AluOp_data_5_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign alu_nan_to_zero_land_6_lpi_1_dfm = (~(IsNaN_5U_10U_nor_5_tmp | (else_AluOp_data_5_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_AluOp_data_5_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_alu_op_1_sva_1[9:0]),
      (chn_alu_op_rsci_d_mxwt[89:80]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_4_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]),
      (chn_alu_op_rsci_d_mxwt[78:74]), cfg_alu_src_1_sva_st);
  assign IsNaN_5U_10U_nor_4_tmp = ~((else_AluOp_data_4_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign alu_nan_to_zero_land_5_lpi_1_dfm = (~(IsNaN_5U_10U_nor_4_tmp | (else_AluOp_data_4_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_AluOp_data_4_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_alu_op_1_sva_1[9:0]),
      (chn_alu_op_rsci_d_mxwt[73:64]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_3_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]),
      (chn_alu_op_rsci_d_mxwt[62:58]), cfg_alu_src_1_sva_st);
  assign IsNaN_5U_10U_nor_3_tmp = ~((else_AluOp_data_3_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign alu_nan_to_zero_land_4_lpi_1_dfm = (~(IsNaN_5U_10U_nor_3_tmp | (else_AluOp_data_3_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_AluOp_data_3_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_alu_op_1_sva_1[9:0]),
      (chn_alu_op_rsci_d_mxwt[57:48]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_2_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]),
      (chn_alu_op_rsci_d_mxwt[46:42]), cfg_alu_src_1_sva_st);
  assign IsNaN_5U_10U_nor_2_tmp = ~((else_AluOp_data_2_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign alu_nan_to_zero_land_3_lpi_1_dfm = (~(IsNaN_5U_10U_nor_2_tmp | (else_AluOp_data_2_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_AluOp_data_2_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_alu_op_1_sva_1[9:0]),
      (chn_alu_op_rsci_d_mxwt[41:32]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_1_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]),
      (chn_alu_op_rsci_d_mxwt[30:26]), cfg_alu_src_1_sva_st);
  assign IsNaN_5U_10U_nor_1_tmp = ~((else_AluOp_data_1_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign alu_nan_to_zero_land_2_lpi_1_dfm = (~(IsNaN_5U_10U_nor_1_tmp | (else_AluOp_data_1_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_AluOp_data_1_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_alu_op_1_sva_1[9:0]),
      (chn_alu_op_rsci_d_mxwt[25:16]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_0_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]),
      (chn_alu_op_rsci_d_mxwt[14:10]), cfg_alu_src_1_sva_st);
  assign IsNaN_5U_10U_nor_tmp = ~((else_AluOp_data_0_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign alu_nan_to_zero_land_1_lpi_1_dfm = (~(IsNaN_5U_10U_nor_tmp | (else_AluOp_data_0_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_AluOp_data_0_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_alu_op_1_sva_1[9:0]),
      (chn_alu_op_rsci_d_mxwt[9:0]), cfg_alu_src_1_sva_st);
  assign and_91_tmp = chn_alu_in_rsci_bawt & or_4_cse & or_5_cse & or_6_cse & or_7_cse
      & or_8_cse & or_9_cse & or_cse_2;
  assign or_4_cse = chn_alu_op_rsci_bawt | (~(cfg_alu_src_1_sva_st_1 & (~ io_read_cfg_alu_bypass_rsc_svs_st_1)
      & main_stage_v_1));
  assign or_5_cse = cfg_alu_shift_value_rsc_triosy_obj_bawt | (~ main_stage_v_1);
  assign or_6_cse = cfg_alu_src_rsc_triosy_obj_bawt | (~ main_stage_v_1);
  assign or_7_cse = cfg_alu_algo_rsc_triosy_obj_bawt | (~ main_stage_v_1);
  assign or_8_cse = cfg_alu_bypass_rsc_triosy_obj_bawt | (~ main_stage_v_1);
  assign or_9_cse = cfg_alu_op_rsc_triosy_obj_bawt | (~ main_stage_v_1);
  assign FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_16,
      FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w4);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_158_nl = ~ FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w4;
  assign FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_16,
      (FpAdd_8U_23U_is_a_greater_oelse_not_158_nl));
  assign FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_18,
      FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w4);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_159_nl = ~ FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w4;
  assign FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_18,
      (FpAdd_8U_23U_is_a_greater_oelse_not_159_nl));
  assign FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_20,
      FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w4);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_160_nl = ~ FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w4;
  assign FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_20,
      (FpAdd_8U_23U_is_a_greater_oelse_not_160_nl));
  assign FpAdd_8U_23U_b_right_shift_qr_4_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_22,
      FpAdd_8U_23U_is_a_greater_lor_4_lpi_1_dfm_1_mx0w4);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_161_nl = ~ FpAdd_8U_23U_is_a_greater_lor_4_lpi_1_dfm_1_mx0w4;
  assign FpAdd_8U_23U_a_right_shift_qr_4_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_22,
      (FpAdd_8U_23U_is_a_greater_oelse_not_161_nl));
  assign FpAdd_8U_23U_b_right_shift_qr_5_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_24,
      FpAdd_8U_23U_is_a_greater_lor_5_lpi_1_dfm_1_mx0w4);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_162_nl = ~ FpAdd_8U_23U_is_a_greater_lor_5_lpi_1_dfm_1_mx0w4;
  assign FpAdd_8U_23U_a_right_shift_qr_5_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_24,
      (FpAdd_8U_23U_is_a_greater_oelse_not_162_nl));
  assign FpAdd_8U_23U_b_right_shift_qr_6_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_26,
      FpAdd_8U_23U_is_a_greater_lor_6_lpi_1_dfm_1_mx0w4);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_163_nl = ~ FpAdd_8U_23U_is_a_greater_lor_6_lpi_1_dfm_1_mx0w4;
  assign FpAdd_8U_23U_a_right_shift_qr_6_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_26,
      (FpAdd_8U_23U_is_a_greater_oelse_not_163_nl));
  assign FpAdd_8U_23U_b_right_shift_qr_7_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_28,
      FpAdd_8U_23U_is_a_greater_lor_7_lpi_1_dfm_1_mx0w4);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_164_nl = ~ FpAdd_8U_23U_is_a_greater_lor_7_lpi_1_dfm_1_mx0w4;
  assign FpAdd_8U_23U_a_right_shift_qr_7_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_28,
      (FpAdd_8U_23U_is_a_greater_oelse_not_164_nl));
  assign FpAdd_8U_23U_b_right_shift_qr_8_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_30,
      FpAdd_8U_23U_is_a_greater_lor_8_lpi_1_dfm_1_mx0w4);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_165_nl = ~ FpAdd_8U_23U_is_a_greater_lor_8_lpi_1_dfm_1_mx0w4;
  assign FpAdd_8U_23U_a_right_shift_qr_8_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_30,
      (FpAdd_8U_23U_is_a_greater_oelse_not_165_nl));
  assign FpAdd_8U_23U_b_right_shift_qr_9_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_31,
      FpAdd_8U_23U_is_a_greater_lor_9_lpi_1_dfm_1_mx0w4);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_166_nl = ~ FpAdd_8U_23U_is_a_greater_lor_9_lpi_1_dfm_1_mx0w4;
  assign FpAdd_8U_23U_a_right_shift_qr_9_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_31,
      (FpAdd_8U_23U_is_a_greater_oelse_not_166_nl));
  assign FpAdd_8U_23U_b_right_shift_qr_10_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_29,
      FpAdd_8U_23U_is_a_greater_lor_10_lpi_1_dfm_1_mx0w4);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_167_nl = ~ FpAdd_8U_23U_is_a_greater_lor_10_lpi_1_dfm_1_mx0w4;
  assign FpAdd_8U_23U_a_right_shift_qr_10_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_29,
      (FpAdd_8U_23U_is_a_greater_oelse_not_167_nl));
  assign FpAdd_8U_23U_b_right_shift_qr_11_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_27,
      FpAdd_8U_23U_is_a_greater_lor_11_lpi_1_dfm_1_mx0w4);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_168_nl = ~ FpAdd_8U_23U_is_a_greater_lor_11_lpi_1_dfm_1_mx0w4;
  assign FpAdd_8U_23U_a_right_shift_qr_11_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_27,
      (FpAdd_8U_23U_is_a_greater_oelse_not_168_nl));
  assign FpAdd_8U_23U_b_right_shift_qr_12_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_25,
      FpAdd_8U_23U_is_a_greater_lor_12_lpi_1_dfm_1_mx0w4);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_169_nl = ~ FpAdd_8U_23U_is_a_greater_lor_12_lpi_1_dfm_1_mx0w4;
  assign FpAdd_8U_23U_a_right_shift_qr_12_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_25,
      (FpAdd_8U_23U_is_a_greater_oelse_not_169_nl));
  assign FpAdd_8U_23U_b_right_shift_qr_13_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_23,
      FpAdd_8U_23U_is_a_greater_lor_13_lpi_1_dfm_1_mx0w4);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_170_nl = ~ FpAdd_8U_23U_is_a_greater_lor_13_lpi_1_dfm_1_mx0w4;
  assign FpAdd_8U_23U_a_right_shift_qr_13_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_23,
      (FpAdd_8U_23U_is_a_greater_oelse_not_170_nl));
  assign FpAdd_8U_23U_b_right_shift_qr_14_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_21,
      FpAdd_8U_23U_is_a_greater_lor_14_lpi_1_dfm_1_mx0w4);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_171_nl = ~ FpAdd_8U_23U_is_a_greater_lor_14_lpi_1_dfm_1_mx0w4;
  assign FpAdd_8U_23U_a_right_shift_qr_14_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_21,
      (FpAdd_8U_23U_is_a_greater_oelse_not_171_nl));
  assign FpAdd_8U_23U_b_right_shift_qr_15_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_19,
      FpAdd_8U_23U_is_a_greater_lor_15_lpi_1_dfm_1_mx0w4);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_172_nl = ~ FpAdd_8U_23U_is_a_greater_lor_15_lpi_1_dfm_1_mx0w4;
  assign FpAdd_8U_23U_a_right_shift_qr_15_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_19,
      (FpAdd_8U_23U_is_a_greater_oelse_not_172_nl));
  assign FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_17,
      FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w4);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_173_nl = ~ FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w4;
  assign FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_17,
      (FpAdd_8U_23U_is_a_greater_oelse_not_173_nl));
  assign FpCmp_8U_23U_true_is_a_greater_1_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_mx0w3,
      FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_mx0w2, AluIn_data_sva_501[31]);
  assign FpCmp_8U_23U_false_is_a_greater_1_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_mx0w1,
      FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_mx0w0, AluIn_data_sva_501[31]);
  assign FpCmp_8U_23U_true_is_a_greater_2_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_1_mx0w3,
      FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_1_mx0w2, AluIn_data_sva_501[63]);
  assign FpCmp_8U_23U_false_is_a_greater_2_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_1_mx0w1,
      FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_1_mx0w0, AluIn_data_sva_501[63]);
  assign FpCmp_8U_23U_true_is_a_greater_3_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_2_mx0w3,
      FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_2_mx0w2, AluIn_data_sva_501[95]);
  assign FpCmp_8U_23U_false_is_a_greater_3_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_2_mx0w1,
      FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_2_mx0w0, AluIn_data_sva_501[95]);
  assign FpCmp_8U_23U_true_is_a_greater_4_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_3_mx0w3,
      FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_3_mx0w2, AluIn_data_sva_501[127]);
  assign FpCmp_8U_23U_false_is_a_greater_4_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_3_mx0w1,
      FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_3_mx0w0, AluIn_data_sva_501[127]);
  assign FpCmp_8U_23U_true_is_a_greater_5_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_4_mx0w3,
      FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_4_mx0w2, AluIn_data_sva_501[159]);
  assign FpCmp_8U_23U_false_is_a_greater_5_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_4_mx0w1,
      FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_4_mx0w0, AluIn_data_sva_501[159]);
  assign FpCmp_8U_23U_true_is_a_greater_6_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_5_mx0w3,
      FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_5_mx0w2, AluIn_data_sva_501[191]);
  assign FpCmp_8U_23U_false_is_a_greater_6_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_5_mx0w1,
      FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_5_mx0w0, AluIn_data_sva_501[191]);
  assign FpCmp_8U_23U_true_is_a_greater_7_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_6_mx0w3,
      FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_6_mx0w2, AluIn_data_sva_501[223]);
  assign FpCmp_8U_23U_false_is_a_greater_7_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_6_mx0w1,
      FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_6_mx0w0, AluIn_data_sva_501[223]);
  assign FpCmp_8U_23U_true_is_a_greater_8_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_7_mx0w3,
      FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_7_mx0w2, AluIn_data_sva_501[255]);
  assign FpCmp_8U_23U_false_is_a_greater_8_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_7_mx0w1,
      FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_7_mx0w0, AluIn_data_sva_501[255]);
  assign FpCmp_8U_23U_true_is_a_greater_9_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_8_mx0w3,
      FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_8_mx0w2, AluIn_data_sva_501[287]);
  assign FpCmp_8U_23U_false_is_a_greater_9_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_8_mx0w1,
      FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_8_mx0w0, AluIn_data_sva_501[287]);
  assign FpCmp_8U_23U_true_is_a_greater_10_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_9_mx0w3,
      FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_9_mx0w2, AluIn_data_sva_501[319]);
  assign FpCmp_8U_23U_false_is_a_greater_10_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_9_mx0w1,
      FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_9_mx0w0, AluIn_data_sva_501[319]);
  assign FpCmp_8U_23U_true_is_a_greater_11_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_10_mx0w3,
      FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_10_mx0w2, AluIn_data_sva_501[351]);
  assign FpCmp_8U_23U_false_is_a_greater_11_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_10_mx0w1,
      FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_10_mx0w0, AluIn_data_sva_501[351]);
  assign FpCmp_8U_23U_true_is_a_greater_12_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_11_mx0w3,
      FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_11_mx0w2, AluIn_data_sva_501[383]);
  assign FpCmp_8U_23U_false_is_a_greater_12_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_11_mx0w1,
      FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_11_mx0w0, AluIn_data_sva_501[383]);
  assign FpCmp_8U_23U_true_is_a_greater_13_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_12_mx0w3,
      FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_12_mx0w2, AluIn_data_sva_501[415]);
  assign FpCmp_8U_23U_false_is_a_greater_13_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_12_mx0w1,
      FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_12_mx0w0, AluIn_data_sva_501[415]);
  assign FpCmp_8U_23U_true_is_a_greater_14_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_13_mx0w3,
      FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_13_mx0w2, AluIn_data_sva_501[447]);
  assign FpCmp_8U_23U_false_is_a_greater_14_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_13_mx0w1,
      FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_13_mx0w0, AluIn_data_sva_501[447]);
  assign FpCmp_8U_23U_true_is_a_greater_15_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_14_mx0w3,
      FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_14_mx0w2, AluIn_data_sva_501[479]);
  assign FpCmp_8U_23U_false_is_a_greater_15_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_14_mx0w1,
      FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_14_mx0w0, AluIn_data_sva_501[479]);
  assign FpCmp_8U_23U_true_is_a_greater_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_15_mx0w3,
      FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_15_mx0w2, AluIn_data_sva_501[511]);
  assign FpCmp_8U_23U_false_is_a_greater_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_15_mx0w1,
      FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_15_mx0w0, AluIn_data_sva_501[511]);
  assign FpCmp_8U_23U_true_else_if_mux_1_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_16_itm_8_1,
      alu_loop_op_1_FpCmp_8U_23U_true_else_slc_8_svs, alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_st_2);
  assign FpCmp_8U_23U_true_is_abs_a_greater_1_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_16_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_1_nl))) | alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_3_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_16_itm_8_1,
      alu_loop_op_1_FpCmp_8U_23U_false_else_slc_8_svs, alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_st_2);
  assign FpCmp_8U_23U_false_is_abs_a_greater_1_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_16_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_3_nl))) | alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_5_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_18_itm_8_1,
      alu_loop_op_2_FpCmp_8U_23U_true_else_slc_8_1_svs, alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_st_2);
  assign FpCmp_8U_23U_true_is_abs_a_greater_2_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_18_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_5_nl))) | alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_7_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_18_itm_8_1,
      alu_loop_op_2_FpCmp_8U_23U_false_else_slc_8_1_svs, alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_st_2);
  assign FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_18_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_7_nl))) | alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_9_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_20_itm_8_1,
      alu_loop_op_3_FpCmp_8U_23U_true_else_slc_8_svs, alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_st_2);
  assign FpCmp_8U_23U_true_is_abs_a_greater_3_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_20_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_9_nl))) | alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_11_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_20_itm_8_1,
      alu_loop_op_3_FpCmp_8U_23U_false_else_slc_8_svs, alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_st_2);
  assign FpCmp_8U_23U_false_is_abs_a_greater_3_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_20_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_11_nl))) | alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_13_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_22_itm_8_1,
      alu_loop_op_4_FpCmp_8U_23U_true_else_slc_8_1_svs, alu_loop_op_4_FpCmp_8U_23U_false_slc_8_1_svs_st_2);
  assign FpCmp_8U_23U_true_is_abs_a_greater_4_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_22_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_13_nl))) | alu_loop_op_4_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_15_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_22_itm_8_1,
      alu_loop_op_4_FpCmp_8U_23U_false_else_slc_8_1_svs, alu_loop_op_4_FpCmp_8U_23U_false_slc_8_1_svs_st_2);
  assign FpCmp_8U_23U_false_is_abs_a_greater_4_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_22_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_15_nl))) | alu_loop_op_4_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_17_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_24_itm_8_1,
      alu_loop_op_5_FpCmp_8U_23U_true_else_slc_8_svs, alu_loop_op_5_FpCmp_8U_23U_false_slc_8_svs_st_2);
  assign FpCmp_8U_23U_true_is_abs_a_greater_5_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_24_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_17_nl))) | alu_loop_op_5_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_19_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_24_itm_8_1,
      alu_loop_op_5_FpCmp_8U_23U_false_else_slc_8_svs, alu_loop_op_5_FpCmp_8U_23U_false_slc_8_svs_st_2);
  assign FpCmp_8U_23U_false_is_abs_a_greater_5_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_24_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_19_nl))) | alu_loop_op_5_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_21_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_26_itm_8_1,
      alu_loop_op_6_FpCmp_8U_23U_true_else_slc_8_1_svs, alu_loop_op_6_FpCmp_8U_23U_false_slc_8_1_svs_st_2);
  assign FpCmp_8U_23U_true_is_abs_a_greater_6_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_26_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_21_nl))) | alu_loop_op_6_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_23_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_26_itm_8_1,
      alu_loop_op_6_FpCmp_8U_23U_false_else_slc_8_1_svs, alu_loop_op_6_FpCmp_8U_23U_false_slc_8_1_svs_st_2);
  assign FpCmp_8U_23U_false_is_abs_a_greater_6_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_26_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_23_nl))) | alu_loop_op_6_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_25_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_28_itm_8_1,
      alu_loop_op_7_FpCmp_8U_23U_true_else_slc_8_svs, alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_st_2);
  assign FpCmp_8U_23U_true_is_abs_a_greater_7_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_28_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_25_nl))) | alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_27_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_28_itm_8_1,
      alu_loop_op_7_FpCmp_8U_23U_false_else_slc_8_svs, alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_st_2);
  assign FpCmp_8U_23U_false_is_abs_a_greater_7_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_28_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_27_nl))) | alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_29_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_30_itm_8_1,
      alu_loop_op_8_FpCmp_8U_23U_true_else_slc_8_1_svs, alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_st_2);
  assign FpCmp_8U_23U_true_is_abs_a_greater_8_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_30_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_29_nl))) | alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_31_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_30_itm_8_1,
      alu_loop_op_8_FpCmp_8U_23U_false_else_slc_8_1_svs, alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_st_2);
  assign FpCmp_8U_23U_false_is_abs_a_greater_8_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_30_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_31_nl))) | alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_33_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_32_itm_8_1,
      alu_loop_op_9_FpCmp_8U_23U_true_else_slc_8_svs, alu_loop_op_9_FpCmp_8U_23U_false_slc_8_svs_st_2);
  assign FpCmp_8U_23U_true_is_abs_a_greater_9_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_32_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_33_nl))) | alu_loop_op_9_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_35_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_32_itm_8_1,
      alu_loop_op_9_FpCmp_8U_23U_false_else_slc_8_svs, alu_loop_op_9_FpCmp_8U_23U_false_slc_8_svs_st_2);
  assign FpCmp_8U_23U_false_is_abs_a_greater_9_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_32_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_35_nl))) | alu_loop_op_9_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_37_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_34_itm_8_1,
      alu_loop_op_10_FpCmp_8U_23U_true_else_slc_8_1_svs, alu_loop_op_10_FpCmp_8U_23U_false_slc_8_1_svs_st_2);
  assign FpCmp_8U_23U_true_is_abs_a_greater_10_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_34_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_37_nl))) | alu_loop_op_10_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_39_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_34_itm_8_1,
      alu_loop_op_10_FpCmp_8U_23U_false_else_slc_8_1_svs, alu_loop_op_10_FpCmp_8U_23U_false_slc_8_1_svs_st_2);
  assign FpCmp_8U_23U_false_is_abs_a_greater_10_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_34_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_39_nl))) | alu_loop_op_10_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_41_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_36_itm_8_1,
      alu_loop_op_11_FpCmp_8U_23U_true_else_slc_8_svs, alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_st_2);
  assign FpCmp_8U_23U_true_is_abs_a_greater_11_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_36_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_41_nl))) | alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_43_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_36_itm_8_1,
      alu_loop_op_11_FpCmp_8U_23U_false_else_slc_8_svs, alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_st_2);
  assign FpCmp_8U_23U_false_is_abs_a_greater_11_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_36_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_43_nl))) | alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_45_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_38_itm_8_1,
      alu_loop_op_12_FpCmp_8U_23U_true_else_slc_8_1_svs, alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_st_2);
  assign FpCmp_8U_23U_true_is_abs_a_greater_12_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_38_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_45_nl))) | alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_47_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_38_itm_8_1,
      alu_loop_op_12_FpCmp_8U_23U_false_else_slc_8_1_svs, alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_st_2);
  assign FpCmp_8U_23U_false_is_abs_a_greater_12_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_38_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_47_nl))) | alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_49_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_40_itm_8_1,
      alu_loop_op_13_FpCmp_8U_23U_true_else_slc_8_svs, alu_loop_op_13_FpCmp_8U_23U_false_slc_8_svs_st_2);
  assign FpCmp_8U_23U_true_is_abs_a_greater_13_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_40_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_49_nl))) | alu_loop_op_13_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_51_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_40_itm_8_1,
      alu_loop_op_13_FpCmp_8U_23U_false_else_slc_8_svs, alu_loop_op_13_FpCmp_8U_23U_false_slc_8_svs_st_2);
  assign FpCmp_8U_23U_false_is_abs_a_greater_13_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_40_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_51_nl))) | alu_loop_op_13_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_53_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_42_itm_8_1,
      alu_loop_op_14_FpCmp_8U_23U_true_else_slc_8_1_svs, alu_loop_op_14_FpCmp_8U_23U_false_slc_8_1_svs_st_2);
  assign FpCmp_8U_23U_true_is_abs_a_greater_14_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_42_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_53_nl))) | alu_loop_op_14_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_55_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_42_itm_8_1,
      alu_loop_op_14_FpCmp_8U_23U_false_else_slc_8_1_svs, alu_loop_op_14_FpCmp_8U_23U_false_slc_8_1_svs_st_2);
  assign FpCmp_8U_23U_false_is_abs_a_greater_14_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_42_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_55_nl))) | alu_loop_op_14_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_57_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_44_itm_8_1,
      alu_loop_op_15_FpCmp_8U_23U_true_else_slc_8_svs, alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_st_2);
  assign FpCmp_8U_23U_true_is_abs_a_greater_15_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_44_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_57_nl))) | alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_59_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_44_itm_8_1,
      alu_loop_op_15_FpCmp_8U_23U_false_else_slc_8_svs, alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_st_2);
  assign FpCmp_8U_23U_false_is_abs_a_greater_15_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_44_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_59_nl))) | alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_61_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_46_itm_8_1,
      alu_loop_op_16_FpCmp_8U_23U_true_else_slc_8_1_svs, alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_st_2);
  assign FpCmp_8U_23U_true_is_abs_a_greater_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_46_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_61_nl))) | alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_true_else_if_mux_63_nl = MUX_s_1_2_2(FpCmp_8U_23U_false_else_if_acc_46_itm_8_1,
      alu_loop_op_16_FpCmp_8U_23U_false_else_slc_8_1_svs, alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_st_2);
  assign FpCmp_8U_23U_false_is_abs_a_greater_lpi_1_dfm_1 = (FpCmp_8U_23U_false_else_else_if_acc_46_itm_23_1
      & (~ (FpCmp_8U_23U_true_else_if_mux_63_nl))) | alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_2;
  assign FpCmp_8U_23U_true_else_3_and_45_tmp = FpCmp_8U_23U_true_is_a_greater_lpi_1_dfm_2_mx0
      & (~ IsNaN_8U_23U_3_land_lpi_1_dfm_6);
  assign FpAlu_8U_23U_and_276_m1c = (~ IsNaN_8U_23U_4_land_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_277_cse = IsNaN_8U_23U_4_land_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_279_cse = IsNaN_8U_23U_4_land_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_false_else_3_or_45_tmp = FpCmp_8U_23U_false_is_a_greater_lpi_1_dfm_2_mx0
      | IsNaN_8U_23U_3_land_lpi_1_dfm_6;
  assign FpAlu_8U_23U_and_278_m1c = (~ IsNaN_8U_23U_4_land_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_true_else_3_and_42_tmp = FpCmp_8U_23U_true_is_a_greater_15_lpi_1_dfm_2_mx0
      & (~ IsNaN_8U_23U_3_land_15_lpi_1_dfm_6);
  assign FpAlu_8U_23U_and_262_m1c = (~ IsNaN_8U_23U_4_land_15_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_263_cse = IsNaN_8U_23U_4_land_15_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_265_cse = IsNaN_8U_23U_4_land_15_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_false_else_3_or_42_tmp = FpCmp_8U_23U_false_is_a_greater_15_lpi_1_dfm_2_mx0
      | IsNaN_8U_23U_3_land_15_lpi_1_dfm_6;
  assign FpAlu_8U_23U_and_264_m1c = (~ IsNaN_8U_23U_4_land_15_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_true_else_3_and_39_tmp = FpCmp_8U_23U_true_is_a_greater_14_lpi_1_dfm_2_mx0
      & (~ IsNaN_8U_23U_3_land_14_lpi_1_dfm_6);
  assign FpAlu_8U_23U_and_248_m1c = (~ IsNaN_8U_23U_4_land_14_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_249_cse = IsNaN_8U_23U_4_land_14_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_251_cse = IsNaN_8U_23U_4_land_14_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_false_else_3_or_39_tmp = FpCmp_8U_23U_false_is_a_greater_14_lpi_1_dfm_2_mx0
      | IsNaN_8U_23U_3_land_14_lpi_1_dfm_6;
  assign FpAlu_8U_23U_and_250_m1c = (~ IsNaN_8U_23U_4_land_14_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_true_else_3_and_36_tmp = FpCmp_8U_23U_true_is_a_greater_13_lpi_1_dfm_2_mx0
      & (~ IsNaN_8U_23U_3_land_13_lpi_1_dfm_6);
  assign FpAlu_8U_23U_and_234_m1c = (~ IsNaN_8U_23U_4_land_13_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_235_cse = IsNaN_8U_23U_4_land_13_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_237_cse = IsNaN_8U_23U_4_land_13_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_false_else_3_or_36_tmp = FpCmp_8U_23U_false_is_a_greater_13_lpi_1_dfm_2_mx0
      | IsNaN_8U_23U_3_land_13_lpi_1_dfm_6;
  assign FpAlu_8U_23U_and_236_m1c = (~ IsNaN_8U_23U_4_land_13_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_true_else_3_and_33_tmp = FpCmp_8U_23U_true_is_a_greater_12_lpi_1_dfm_2_mx0
      & (~ IsNaN_8U_23U_3_land_12_lpi_1_dfm_6);
  assign FpAlu_8U_23U_and_220_m1c = (~ IsNaN_8U_23U_4_land_12_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_221_cse = IsNaN_8U_23U_4_land_12_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_223_cse = IsNaN_8U_23U_4_land_12_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_false_else_3_or_33_tmp = FpCmp_8U_23U_false_is_a_greater_12_lpi_1_dfm_2_mx0
      | IsNaN_8U_23U_3_land_12_lpi_1_dfm_6;
  assign FpAlu_8U_23U_and_222_m1c = (~ IsNaN_8U_23U_4_land_12_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_true_else_3_and_30_tmp = FpCmp_8U_23U_true_is_a_greater_11_lpi_1_dfm_2_mx0
      & (~ IsNaN_8U_23U_3_land_11_lpi_1_dfm_6);
  assign FpAlu_8U_23U_and_206_m1c = (~ IsNaN_8U_23U_4_land_11_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_207_cse = IsNaN_8U_23U_4_land_11_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_209_cse = IsNaN_8U_23U_4_land_11_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_false_else_3_or_30_tmp = FpCmp_8U_23U_false_is_a_greater_11_lpi_1_dfm_2_mx0
      | IsNaN_8U_23U_3_land_11_lpi_1_dfm_6;
  assign FpAlu_8U_23U_and_208_m1c = (~ IsNaN_8U_23U_4_land_11_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_true_else_3_and_27_tmp = FpCmp_8U_23U_true_is_a_greater_10_lpi_1_dfm_2_mx0
      & (~ IsNaN_8U_23U_3_land_10_lpi_1_dfm_6);
  assign FpAlu_8U_23U_and_192_m1c = (~ IsNaN_8U_23U_4_land_10_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_193_cse = IsNaN_8U_23U_4_land_10_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_195_cse = IsNaN_8U_23U_4_land_10_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_false_else_3_or_27_tmp = FpCmp_8U_23U_false_is_a_greater_10_lpi_1_dfm_2_mx0
      | IsNaN_8U_23U_3_land_10_lpi_1_dfm_6;
  assign FpAlu_8U_23U_and_194_m1c = (~ IsNaN_8U_23U_4_land_10_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_true_else_3_and_24_tmp = FpCmp_8U_23U_true_is_a_greater_9_lpi_1_dfm_2_mx0
      & (~ IsNaN_8U_23U_3_land_9_lpi_1_dfm_6);
  assign FpAlu_8U_23U_and_178_m1c = (~ IsNaN_8U_23U_4_land_9_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_179_cse = IsNaN_8U_23U_4_land_9_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_181_cse = IsNaN_8U_23U_4_land_9_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_false_else_3_or_24_tmp = FpCmp_8U_23U_false_is_a_greater_9_lpi_1_dfm_2_mx0
      | IsNaN_8U_23U_3_land_9_lpi_1_dfm_6;
  assign FpAlu_8U_23U_and_180_m1c = (~ IsNaN_8U_23U_4_land_9_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_true_else_3_and_21_tmp = FpCmp_8U_23U_true_is_a_greater_8_lpi_1_dfm_2_mx0
      & (~ IsNaN_8U_23U_3_land_8_lpi_1_dfm_6);
  assign FpAlu_8U_23U_and_164_m1c = (~ IsNaN_8U_23U_4_land_8_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_165_cse = IsNaN_8U_23U_4_land_8_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_167_cse = IsNaN_8U_23U_4_land_8_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_false_else_3_or_21_tmp = FpCmp_8U_23U_false_is_a_greater_8_lpi_1_dfm_2_mx0
      | IsNaN_8U_23U_3_land_8_lpi_1_dfm_6;
  assign FpAlu_8U_23U_and_166_m1c = (~ IsNaN_8U_23U_4_land_8_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_true_else_3_and_18_tmp = FpCmp_8U_23U_true_is_a_greater_7_lpi_1_dfm_2_mx0
      & (~ IsNaN_8U_23U_3_land_7_lpi_1_dfm_6);
  assign FpAlu_8U_23U_and_150_m1c = (~ IsNaN_8U_23U_4_land_7_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_151_cse = IsNaN_8U_23U_4_land_7_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_153_cse = IsNaN_8U_23U_4_land_7_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_false_else_3_or_18_tmp = FpCmp_8U_23U_false_is_a_greater_7_lpi_1_dfm_2_mx0
      | IsNaN_8U_23U_3_land_7_lpi_1_dfm_6;
  assign FpAlu_8U_23U_and_152_m1c = (~ IsNaN_8U_23U_4_land_7_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_true_else_3_and_15_tmp = FpCmp_8U_23U_true_is_a_greater_6_lpi_1_dfm_2_mx0
      & (~ IsNaN_8U_23U_3_land_6_lpi_1_dfm_6);
  assign FpAlu_8U_23U_and_136_m1c = (~ IsNaN_8U_23U_4_land_6_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_137_cse = IsNaN_8U_23U_4_land_6_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_139_cse = IsNaN_8U_23U_4_land_6_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_false_else_3_or_15_tmp = FpCmp_8U_23U_false_is_a_greater_6_lpi_1_dfm_2_mx0
      | IsNaN_8U_23U_3_land_6_lpi_1_dfm_6;
  assign FpAlu_8U_23U_and_138_m1c = (~ IsNaN_8U_23U_4_land_6_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_true_else_3_and_12_tmp = FpCmp_8U_23U_true_is_a_greater_5_lpi_1_dfm_2_mx0
      & (~ IsNaN_8U_23U_3_land_5_lpi_1_dfm_6);
  assign FpAlu_8U_23U_and_122_m1c = (~ IsNaN_8U_23U_4_land_5_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_123_cse = IsNaN_8U_23U_4_land_5_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_125_cse = IsNaN_8U_23U_4_land_5_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_false_else_3_or_12_tmp = FpCmp_8U_23U_false_is_a_greater_5_lpi_1_dfm_2_mx0
      | IsNaN_8U_23U_3_land_5_lpi_1_dfm_6;
  assign FpAlu_8U_23U_and_124_m1c = (~ IsNaN_8U_23U_4_land_5_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_true_else_3_and_9_tmp = FpCmp_8U_23U_true_is_a_greater_4_lpi_1_dfm_2_mx0
      & (~ IsNaN_8U_23U_3_land_4_lpi_1_dfm_6);
  assign FpAlu_8U_23U_and_108_m1c = (~ IsNaN_8U_23U_4_land_4_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_109_cse = IsNaN_8U_23U_4_land_4_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_111_cse = IsNaN_8U_23U_4_land_4_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_false_else_3_or_9_tmp = FpCmp_8U_23U_false_is_a_greater_4_lpi_1_dfm_2_mx0
      | IsNaN_8U_23U_3_land_4_lpi_1_dfm_6;
  assign FpAlu_8U_23U_and_110_m1c = (~ IsNaN_8U_23U_4_land_4_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_true_else_3_and_6_tmp = FpCmp_8U_23U_true_is_a_greater_3_lpi_1_dfm_2_mx0
      & (~ IsNaN_8U_23U_3_land_3_lpi_1_dfm_6);
  assign FpAlu_8U_23U_and_94_m1c = (~ IsNaN_8U_23U_4_land_3_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_95_cse = IsNaN_8U_23U_4_land_3_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_97_cse = IsNaN_8U_23U_4_land_3_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_false_else_3_or_6_tmp = FpCmp_8U_23U_false_is_a_greater_3_lpi_1_dfm_2_mx0
      | IsNaN_8U_23U_3_land_3_lpi_1_dfm_6;
  assign FpAlu_8U_23U_and_96_m1c = (~ IsNaN_8U_23U_4_land_3_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_true_else_3_and_3_tmp = FpCmp_8U_23U_true_is_a_greater_2_lpi_1_dfm_2_mx0
      & (~ IsNaN_8U_23U_3_land_2_lpi_1_dfm_6);
  assign FpAlu_8U_23U_and_80_m1c = (~ IsNaN_8U_23U_4_land_2_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_81_cse = IsNaN_8U_23U_4_land_2_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_83_cse = IsNaN_8U_23U_4_land_2_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_false_else_3_or_3_tmp = FpCmp_8U_23U_false_is_a_greater_2_lpi_1_dfm_2_mx0
      | IsNaN_8U_23U_3_land_2_lpi_1_dfm_6;
  assign FpAlu_8U_23U_and_82_m1c = (~ IsNaN_8U_23U_4_land_2_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_true_else_3_and_tmp = FpCmp_8U_23U_true_is_a_greater_1_lpi_1_dfm_2_mx0
      & (~ IsNaN_8U_23U_3_land_1_lpi_1_dfm_6);
  assign FpAlu_8U_23U_and_66_m1c = (~ IsNaN_8U_23U_4_land_1_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_67_cse = IsNaN_8U_23U_4_land_1_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_mx0w0;
  assign FpAlu_8U_23U_and_69_cse = IsNaN_8U_23U_4_land_1_lpi_1_dfm_6 & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_false_else_3_or_tmp = FpCmp_8U_23U_false_is_a_greater_1_lpi_1_dfm_2_mx0
      | IsNaN_8U_23U_3_land_1_lpi_1_dfm_6;
  assign FpAlu_8U_23U_and_68_m1c = (~ IsNaN_8U_23U_4_land_1_lpi_1_dfm_6) & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign else_AluOp_data_15_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_alu_op_1_sva_1[15]),
      (chn_alu_op_rsci_d_mxwt[255]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_14_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_alu_op_1_sva_1[15]),
      (chn_alu_op_rsci_d_mxwt[239]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_13_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_alu_op_1_sva_1[15]),
      (chn_alu_op_rsci_d_mxwt[223]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_12_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_alu_op_1_sva_1[15]),
      (chn_alu_op_rsci_d_mxwt[207]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_11_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_alu_op_1_sva_1[15]),
      (chn_alu_op_rsci_d_mxwt[191]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_10_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_alu_op_1_sva_1[15]),
      (chn_alu_op_rsci_d_mxwt[175]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_9_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_alu_op_1_sva_1[15]),
      (chn_alu_op_rsci_d_mxwt[159]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_8_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_alu_op_1_sva_1[15]),
      (chn_alu_op_rsci_d_mxwt[143]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_7_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_alu_op_1_sva_1[15]),
      (chn_alu_op_rsci_d_mxwt[127]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_6_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_alu_op_1_sva_1[15]),
      (chn_alu_op_rsci_d_mxwt[111]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_5_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_alu_op_1_sva_1[15]),
      (chn_alu_op_rsci_d_mxwt[95]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_4_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_alu_op_1_sva_1[15]),
      (chn_alu_op_rsci_d_mxwt[79]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_3_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_alu_op_1_sva_1[15]),
      (chn_alu_op_rsci_d_mxwt[63]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_2_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_alu_op_1_sva_1[15]),
      (chn_alu_op_rsci_d_mxwt[47]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_1_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_alu_op_1_sva_1[15]),
      (chn_alu_op_rsci_d_mxwt[31]), cfg_alu_src_1_sva_st);
  assign else_AluOp_data_0_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_alu_op_1_sva_1[15]),
      (chn_alu_op_rsci_d_mxwt[15]), cfg_alu_src_1_sva_st);
  assign IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_sva = (IntShiftLeft_16U_6U_32U_mbits_fixed_sva[78])
      & (~((IntShiftLeft_16U_6U_32U_mbits_fixed_sva[77:31]==47'b11111111111111111111111111111111111111111111111)));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_sva = ~((IntShiftLeft_16U_6U_32U_mbits_fixed_sva[78])
      | (~((IntShiftLeft_16U_6U_32U_mbits_fixed_sva[77:31]!=47'b00000000000000000000000000000000000000000000000))));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_15_sva = (IntShiftLeft_16U_6U_32U_mbits_fixed_15_sva[78])
      & (~((IntShiftLeft_16U_6U_32U_mbits_fixed_15_sva[77:31]==47'b11111111111111111111111111111111111111111111111)));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_15_sva = ~((IntShiftLeft_16U_6U_32U_mbits_fixed_15_sva[78])
      | (~((IntShiftLeft_16U_6U_32U_mbits_fixed_15_sva[77:31]!=47'b00000000000000000000000000000000000000000000000))));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_14_sva = (IntShiftLeft_16U_6U_32U_mbits_fixed_14_sva[78])
      & (~((IntShiftLeft_16U_6U_32U_mbits_fixed_14_sva[77:31]==47'b11111111111111111111111111111111111111111111111)));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_14_sva = ~((IntShiftLeft_16U_6U_32U_mbits_fixed_14_sva[78])
      | (~((IntShiftLeft_16U_6U_32U_mbits_fixed_14_sva[77:31]!=47'b00000000000000000000000000000000000000000000000))));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_13_sva = (IntShiftLeft_16U_6U_32U_mbits_fixed_13_sva[78])
      & (~((IntShiftLeft_16U_6U_32U_mbits_fixed_13_sva[77:31]==47'b11111111111111111111111111111111111111111111111)));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_13_sva = ~((IntShiftLeft_16U_6U_32U_mbits_fixed_13_sva[78])
      | (~((IntShiftLeft_16U_6U_32U_mbits_fixed_13_sva[77:31]!=47'b00000000000000000000000000000000000000000000000))));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_12_sva = (IntShiftLeft_16U_6U_32U_mbits_fixed_12_sva[78])
      & (~((IntShiftLeft_16U_6U_32U_mbits_fixed_12_sva[77:31]==47'b11111111111111111111111111111111111111111111111)));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_12_sva = ~((IntShiftLeft_16U_6U_32U_mbits_fixed_12_sva[78])
      | (~((IntShiftLeft_16U_6U_32U_mbits_fixed_12_sva[77:31]!=47'b00000000000000000000000000000000000000000000000))));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_11_sva = (IntShiftLeft_16U_6U_32U_mbits_fixed_11_sva[78])
      & (~((IntShiftLeft_16U_6U_32U_mbits_fixed_11_sva[77:31]==47'b11111111111111111111111111111111111111111111111)));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_11_sva = ~((IntShiftLeft_16U_6U_32U_mbits_fixed_11_sva[78])
      | (~((IntShiftLeft_16U_6U_32U_mbits_fixed_11_sva[77:31]!=47'b00000000000000000000000000000000000000000000000))));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_10_sva = (IntShiftLeft_16U_6U_32U_mbits_fixed_10_sva[78])
      & (~((IntShiftLeft_16U_6U_32U_mbits_fixed_10_sva[77:31]==47'b11111111111111111111111111111111111111111111111)));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_10_sva = ~((IntShiftLeft_16U_6U_32U_mbits_fixed_10_sva[78])
      | (~((IntShiftLeft_16U_6U_32U_mbits_fixed_10_sva[77:31]!=47'b00000000000000000000000000000000000000000000000))));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_9_sva = (IntShiftLeft_16U_6U_32U_mbits_fixed_9_sva[78])
      & (~((IntShiftLeft_16U_6U_32U_mbits_fixed_9_sva[77:31]==47'b11111111111111111111111111111111111111111111111)));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_9_sva = ~((IntShiftLeft_16U_6U_32U_mbits_fixed_9_sva[78])
      | (~((IntShiftLeft_16U_6U_32U_mbits_fixed_9_sva[77:31]!=47'b00000000000000000000000000000000000000000000000))));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_8_sva = (IntShiftLeft_16U_6U_32U_mbits_fixed_8_sva[78])
      & (~((IntShiftLeft_16U_6U_32U_mbits_fixed_8_sva[77:31]==47'b11111111111111111111111111111111111111111111111)));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_8_sva = ~((IntShiftLeft_16U_6U_32U_mbits_fixed_8_sva[78])
      | (~((IntShiftLeft_16U_6U_32U_mbits_fixed_8_sva[77:31]!=47'b00000000000000000000000000000000000000000000000))));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_7_sva = (IntShiftLeft_16U_6U_32U_mbits_fixed_7_sva[78])
      & (~((IntShiftLeft_16U_6U_32U_mbits_fixed_7_sva[77:31]==47'b11111111111111111111111111111111111111111111111)));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_7_sva = ~((IntShiftLeft_16U_6U_32U_mbits_fixed_7_sva[78])
      | (~((IntShiftLeft_16U_6U_32U_mbits_fixed_7_sva[77:31]!=47'b00000000000000000000000000000000000000000000000))));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_6_sva = (IntShiftLeft_16U_6U_32U_mbits_fixed_6_sva[78])
      & (~((IntShiftLeft_16U_6U_32U_mbits_fixed_6_sva[77:31]==47'b11111111111111111111111111111111111111111111111)));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_6_sva = ~((IntShiftLeft_16U_6U_32U_mbits_fixed_6_sva[78])
      | (~((IntShiftLeft_16U_6U_32U_mbits_fixed_6_sva[77:31]!=47'b00000000000000000000000000000000000000000000000))));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_5_sva = (IntShiftLeft_16U_6U_32U_mbits_fixed_5_sva[78])
      & (~((IntShiftLeft_16U_6U_32U_mbits_fixed_5_sva[77:31]==47'b11111111111111111111111111111111111111111111111)));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_5_sva = ~((IntShiftLeft_16U_6U_32U_mbits_fixed_5_sva[78])
      | (~((IntShiftLeft_16U_6U_32U_mbits_fixed_5_sva[77:31]!=47'b00000000000000000000000000000000000000000000000))));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_4_sva = (IntShiftLeft_16U_6U_32U_mbits_fixed_4_sva[78])
      & (~((IntShiftLeft_16U_6U_32U_mbits_fixed_4_sva[77:31]==47'b11111111111111111111111111111111111111111111111)));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_4_sva = ~((IntShiftLeft_16U_6U_32U_mbits_fixed_4_sva[78])
      | (~((IntShiftLeft_16U_6U_32U_mbits_fixed_4_sva[77:31]!=47'b00000000000000000000000000000000000000000000000))));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_3_sva = (IntShiftLeft_16U_6U_32U_mbits_fixed_3_sva[78])
      & (~((IntShiftLeft_16U_6U_32U_mbits_fixed_3_sva[77:31]==47'b11111111111111111111111111111111111111111111111)));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_3_sva = ~((IntShiftLeft_16U_6U_32U_mbits_fixed_3_sva[78])
      | (~((IntShiftLeft_16U_6U_32U_mbits_fixed_3_sva[77:31]!=47'b00000000000000000000000000000000000000000000000))));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_2_sva = (IntShiftLeft_16U_6U_32U_mbits_fixed_2_sva[78])
      & (~((IntShiftLeft_16U_6U_32U_mbits_fixed_2_sva[77:31]==47'b11111111111111111111111111111111111111111111111)));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_2_sva = ~((IntShiftLeft_16U_6U_32U_mbits_fixed_2_sva[78])
      | (~((IntShiftLeft_16U_6U_32U_mbits_fixed_2_sva[77:31]!=47'b00000000000000000000000000000000000000000000000))));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_and_unfl_1_sva = (IntShiftLeft_16U_6U_32U_mbits_fixed_1_sva[78])
      & (~((IntShiftLeft_16U_6U_32U_mbits_fixed_1_sva[77:31]==47'b11111111111111111111111111111111111111111111111)));
  assign IntShiftLeft_16U_6U_32U_obits_fixed_nor_ovfl_1_sva = ~((IntShiftLeft_16U_6U_32U_mbits_fixed_1_sva[78])
      | (~((IntShiftLeft_16U_6U_32U_mbits_fixed_1_sva[77:31]!=47'b00000000000000000000000000000000000000000000000))));
  assign nl_FpCmp_8U_23U_false_else_else_if_acc_16_nl = ({1'b1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp_2})
      + conv_u2u_23_24(~ (AluIn_data_sva_501[22:0])) + 24'b1;
  assign FpCmp_8U_23U_false_else_else_if_acc_16_nl = nl_FpCmp_8U_23U_false_else_else_if_acc_16_nl[23:0];
  assign FpCmp_8U_23U_false_else_else_if_acc_16_itm_23_1 = readslicef_24_1_23((FpCmp_8U_23U_false_else_else_if_acc_16_nl));
  assign nl_FpCmp_8U_23U_false_else_if_acc_16_nl = ({1'b1 , (AluIn_data_sva_501[30:23])})
      + conv_u2u_8_9({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_9)}) + 9'b1;
  assign FpCmp_8U_23U_false_else_if_acc_16_nl = nl_FpCmp_8U_23U_false_else_if_acc_16_nl[8:0];
  assign FpCmp_8U_23U_false_else_if_acc_16_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_false_else_if_acc_16_nl));
  assign nl_FpCmp_8U_23U_false_else_else_if_acc_18_nl = ({1'b1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp_2})
      + conv_u2u_23_24(~ (AluIn_data_sva_501[54:32])) + 24'b1;
  assign FpCmp_8U_23U_false_else_else_if_acc_18_nl = nl_FpCmp_8U_23U_false_else_else_if_acc_18_nl[23:0];
  assign FpCmp_8U_23U_false_else_else_if_acc_18_itm_23_1 = readslicef_24_1_23((FpCmp_8U_23U_false_else_else_if_acc_18_nl));
  assign nl_FpCmp_8U_23U_false_else_if_acc_18_nl = ({1'b1 , (AluIn_data_sva_501[62:55])})
      + conv_u2u_8_9({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_9)}) + 9'b1;
  assign FpCmp_8U_23U_false_else_if_acc_18_nl = nl_FpCmp_8U_23U_false_else_if_acc_18_nl[8:0];
  assign FpCmp_8U_23U_false_else_if_acc_18_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_false_else_if_acc_18_nl));
  assign nl_FpCmp_8U_23U_false_else_else_if_acc_20_nl = ({1'b1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp_2})
      + conv_u2u_23_24(~ (AluIn_data_sva_501[86:64])) + 24'b1;
  assign FpCmp_8U_23U_false_else_else_if_acc_20_nl = nl_FpCmp_8U_23U_false_else_else_if_acc_20_nl[23:0];
  assign FpCmp_8U_23U_false_else_else_if_acc_20_itm_23_1 = readslicef_24_1_23((FpCmp_8U_23U_false_else_else_if_acc_20_nl));
  assign nl_FpCmp_8U_23U_false_else_if_acc_20_nl = ({1'b1 , (AluIn_data_sva_501[94:87])})
      + conv_u2u_8_9({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_9)}) + 9'b1;
  assign FpCmp_8U_23U_false_else_if_acc_20_nl = nl_FpCmp_8U_23U_false_else_if_acc_20_nl[8:0];
  assign FpCmp_8U_23U_false_else_if_acc_20_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_false_else_if_acc_20_nl));
  assign nl_FpCmp_8U_23U_false_else_else_if_acc_22_nl = ({1'b1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp_2})
      + conv_u2u_23_24(~ (AluIn_data_sva_501[118:96])) + 24'b1;
  assign FpCmp_8U_23U_false_else_else_if_acc_22_nl = nl_FpCmp_8U_23U_false_else_else_if_acc_22_nl[23:0];
  assign FpCmp_8U_23U_false_else_else_if_acc_22_itm_23_1 = readslicef_24_1_23((FpCmp_8U_23U_false_else_else_if_acc_22_nl));
  assign nl_FpCmp_8U_23U_false_else_if_acc_22_nl = ({1'b1 , (AluIn_data_sva_501[126:119])})
      + conv_u2u_8_9({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_9)}) + 9'b1;
  assign FpCmp_8U_23U_false_else_if_acc_22_nl = nl_FpCmp_8U_23U_false_else_if_acc_22_nl[8:0];
  assign FpCmp_8U_23U_false_else_if_acc_22_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_false_else_if_acc_22_nl));
  assign nl_FpCmp_8U_23U_false_else_else_if_acc_24_nl = ({1'b1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp_2})
      + conv_u2u_23_24(~ (AluIn_data_sva_501[150:128])) + 24'b1;
  assign FpCmp_8U_23U_false_else_else_if_acc_24_nl = nl_FpCmp_8U_23U_false_else_else_if_acc_24_nl[23:0];
  assign FpCmp_8U_23U_false_else_else_if_acc_24_itm_23_1 = readslicef_24_1_23((FpCmp_8U_23U_false_else_else_if_acc_24_nl));
  assign nl_FpCmp_8U_23U_false_else_if_acc_24_nl = ({1'b1 , (AluIn_data_sva_501[158:151])})
      + conv_u2u_8_9({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_9)}) + 9'b1;
  assign FpCmp_8U_23U_false_else_if_acc_24_nl = nl_FpCmp_8U_23U_false_else_if_acc_24_nl[8:0];
  assign FpCmp_8U_23U_false_else_if_acc_24_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_false_else_if_acc_24_nl));
  assign nl_FpCmp_8U_23U_false_else_else_if_acc_26_nl = ({1'b1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp_2})
      + conv_u2u_23_24(~ (AluIn_data_sva_501[182:160])) + 24'b1;
  assign FpCmp_8U_23U_false_else_else_if_acc_26_nl = nl_FpCmp_8U_23U_false_else_else_if_acc_26_nl[23:0];
  assign FpCmp_8U_23U_false_else_else_if_acc_26_itm_23_1 = readslicef_24_1_23((FpCmp_8U_23U_false_else_else_if_acc_26_nl));
  assign nl_FpCmp_8U_23U_false_else_if_acc_26_nl = ({1'b1 , (AluIn_data_sva_501[190:183])})
      + conv_u2u_8_9({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_9)}) + 9'b1;
  assign FpCmp_8U_23U_false_else_if_acc_26_nl = nl_FpCmp_8U_23U_false_else_if_acc_26_nl[8:0];
  assign FpCmp_8U_23U_false_else_if_acc_26_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_false_else_if_acc_26_nl));
  assign nl_FpCmp_8U_23U_false_else_else_if_acc_28_nl = ({1'b1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp_2})
      + conv_u2u_23_24(~ (AluIn_data_sva_501[214:192])) + 24'b1;
  assign FpCmp_8U_23U_false_else_else_if_acc_28_nl = nl_FpCmp_8U_23U_false_else_else_if_acc_28_nl[23:0];
  assign FpCmp_8U_23U_false_else_else_if_acc_28_itm_23_1 = readslicef_24_1_23((FpCmp_8U_23U_false_else_else_if_acc_28_nl));
  assign nl_FpCmp_8U_23U_false_else_if_acc_28_nl = ({1'b1 , (AluIn_data_sva_501[222:215])})
      + conv_u2u_8_9({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_9)}) + 9'b1;
  assign FpCmp_8U_23U_false_else_if_acc_28_nl = nl_FpCmp_8U_23U_false_else_if_acc_28_nl[8:0];
  assign FpCmp_8U_23U_false_else_if_acc_28_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_false_else_if_acc_28_nl));
  assign nl_FpCmp_8U_23U_false_else_else_if_acc_30_nl = ({1'b1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp_2})
      + conv_u2u_23_24(~ (AluIn_data_sva_501[246:224])) + 24'b1;
  assign FpCmp_8U_23U_false_else_else_if_acc_30_nl = nl_FpCmp_8U_23U_false_else_else_if_acc_30_nl[23:0];
  assign FpCmp_8U_23U_false_else_else_if_acc_30_itm_23_1 = readslicef_24_1_23((FpCmp_8U_23U_false_else_else_if_acc_30_nl));
  assign nl_FpCmp_8U_23U_false_else_if_acc_30_nl = ({1'b1 , (AluIn_data_sva_501[254:247])})
      + conv_u2u_8_9({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_9)}) + 9'b1;
  assign FpCmp_8U_23U_false_else_if_acc_30_nl = nl_FpCmp_8U_23U_false_else_if_acc_30_nl[8:0];
  assign FpCmp_8U_23U_false_else_if_acc_30_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_false_else_if_acc_30_nl));
  assign nl_FpCmp_8U_23U_false_else_else_if_acc_32_nl = ({1'b1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp_2})
      + conv_u2u_23_24(~ (AluIn_data_sva_501[278:256])) + 24'b1;
  assign FpCmp_8U_23U_false_else_else_if_acc_32_nl = nl_FpCmp_8U_23U_false_else_else_if_acc_32_nl[23:0];
  assign FpCmp_8U_23U_false_else_else_if_acc_32_itm_23_1 = readslicef_24_1_23((FpCmp_8U_23U_false_else_else_if_acc_32_nl));
  assign nl_FpCmp_8U_23U_false_else_if_acc_32_nl = ({1'b1 , (AluIn_data_sva_501[286:279])})
      + conv_u2u_8_9({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_9)}) + 9'b1;
  assign FpCmp_8U_23U_false_else_if_acc_32_nl = nl_FpCmp_8U_23U_false_else_if_acc_32_nl[8:0];
  assign FpCmp_8U_23U_false_else_if_acc_32_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_false_else_if_acc_32_nl));
  assign nl_FpCmp_8U_23U_false_else_else_if_acc_34_nl = ({1'b1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp_2})
      + conv_u2u_23_24(~ (AluIn_data_sva_501[310:288])) + 24'b1;
  assign FpCmp_8U_23U_false_else_else_if_acc_34_nl = nl_FpCmp_8U_23U_false_else_else_if_acc_34_nl[23:0];
  assign FpCmp_8U_23U_false_else_else_if_acc_34_itm_23_1 = readslicef_24_1_23((FpCmp_8U_23U_false_else_else_if_acc_34_nl));
  assign nl_FpCmp_8U_23U_false_else_if_acc_34_nl = ({1'b1 , (AluIn_data_sva_501[318:311])})
      + conv_u2u_8_9({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_9)}) + 9'b1;
  assign FpCmp_8U_23U_false_else_if_acc_34_nl = nl_FpCmp_8U_23U_false_else_if_acc_34_nl[8:0];
  assign FpCmp_8U_23U_false_else_if_acc_34_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_false_else_if_acc_34_nl));
  assign nl_FpCmp_8U_23U_false_else_else_if_acc_36_nl = ({1'b1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp_2})
      + conv_u2u_23_24(~ (AluIn_data_sva_501[342:320])) + 24'b1;
  assign FpCmp_8U_23U_false_else_else_if_acc_36_nl = nl_FpCmp_8U_23U_false_else_else_if_acc_36_nl[23:0];
  assign FpCmp_8U_23U_false_else_else_if_acc_36_itm_23_1 = readslicef_24_1_23((FpCmp_8U_23U_false_else_else_if_acc_36_nl));
  assign nl_FpCmp_8U_23U_false_else_if_acc_36_nl = ({1'b1 , (AluIn_data_sva_501[350:343])})
      + conv_u2u_8_9({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_9)}) + 9'b1;
  assign FpCmp_8U_23U_false_else_if_acc_36_nl = nl_FpCmp_8U_23U_false_else_if_acc_36_nl[8:0];
  assign FpCmp_8U_23U_false_else_if_acc_36_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_false_else_if_acc_36_nl));
  assign nl_FpCmp_8U_23U_false_else_else_if_acc_38_nl = ({1'b1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp_2})
      + conv_u2u_23_24(~ (AluIn_data_sva_501[374:352])) + 24'b1;
  assign FpCmp_8U_23U_false_else_else_if_acc_38_nl = nl_FpCmp_8U_23U_false_else_else_if_acc_38_nl[23:0];
  assign FpCmp_8U_23U_false_else_else_if_acc_38_itm_23_1 = readslicef_24_1_23((FpCmp_8U_23U_false_else_else_if_acc_38_nl));
  assign nl_FpCmp_8U_23U_false_else_if_acc_38_nl = ({1'b1 , (AluIn_data_sva_501[382:375])})
      + conv_u2u_8_9({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_9)}) + 9'b1;
  assign FpCmp_8U_23U_false_else_if_acc_38_nl = nl_FpCmp_8U_23U_false_else_if_acc_38_nl[8:0];
  assign FpCmp_8U_23U_false_else_if_acc_38_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_false_else_if_acc_38_nl));
  assign nl_FpCmp_8U_23U_false_else_else_if_acc_40_nl = ({1'b1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp_2})
      + conv_u2u_23_24(~ (AluIn_data_sva_501[406:384])) + 24'b1;
  assign FpCmp_8U_23U_false_else_else_if_acc_40_nl = nl_FpCmp_8U_23U_false_else_else_if_acc_40_nl[23:0];
  assign FpCmp_8U_23U_false_else_else_if_acc_40_itm_23_1 = readslicef_24_1_23((FpCmp_8U_23U_false_else_else_if_acc_40_nl));
  assign nl_FpCmp_8U_23U_false_else_if_acc_40_nl = ({1'b1 , (AluIn_data_sva_501[414:407])})
      + conv_u2u_8_9({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_9)}) + 9'b1;
  assign FpCmp_8U_23U_false_else_if_acc_40_nl = nl_FpCmp_8U_23U_false_else_if_acc_40_nl[8:0];
  assign FpCmp_8U_23U_false_else_if_acc_40_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_false_else_if_acc_40_nl));
  assign nl_FpCmp_8U_23U_false_else_else_if_acc_42_nl = ({1'b1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp_2})
      + conv_u2u_23_24(~ (AluIn_data_sva_501[438:416])) + 24'b1;
  assign FpCmp_8U_23U_false_else_else_if_acc_42_nl = nl_FpCmp_8U_23U_false_else_else_if_acc_42_nl[23:0];
  assign FpCmp_8U_23U_false_else_else_if_acc_42_itm_23_1 = readslicef_24_1_23((FpCmp_8U_23U_false_else_else_if_acc_42_nl));
  assign nl_FpCmp_8U_23U_false_else_if_acc_42_nl = ({1'b1 , (AluIn_data_sva_501[446:439])})
      + conv_u2u_8_9({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_9)}) + 9'b1;
  assign FpCmp_8U_23U_false_else_if_acc_42_nl = nl_FpCmp_8U_23U_false_else_if_acc_42_nl[8:0];
  assign FpCmp_8U_23U_false_else_if_acc_42_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_false_else_if_acc_42_nl));
  assign nl_FpCmp_8U_23U_false_else_else_if_acc_44_nl = ({1'b1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp_2})
      + conv_u2u_23_24(~ (AluIn_data_sva_501[470:448])) + 24'b1;
  assign FpCmp_8U_23U_false_else_else_if_acc_44_nl = nl_FpCmp_8U_23U_false_else_else_if_acc_44_nl[23:0];
  assign FpCmp_8U_23U_false_else_else_if_acc_44_itm_23_1 = readslicef_24_1_23((FpCmp_8U_23U_false_else_else_if_acc_44_nl));
  assign nl_FpCmp_8U_23U_false_else_if_acc_44_nl = ({1'b1 , (AluIn_data_sva_501[478:471])})
      + conv_u2u_8_9({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_9)}) + 9'b1;
  assign FpCmp_8U_23U_false_else_if_acc_44_nl = nl_FpCmp_8U_23U_false_else_if_acc_44_nl[8:0];
  assign FpCmp_8U_23U_false_else_if_acc_44_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_false_else_if_acc_44_nl));
  assign nl_FpCmp_8U_23U_false_else_else_if_acc_46_nl = ({1'b1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp
      , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp_2})
      + conv_u2u_23_24(~ (AluIn_data_sva_501[502:480])) + 24'b1;
  assign FpCmp_8U_23U_false_else_else_if_acc_46_nl = nl_FpCmp_8U_23U_false_else_else_if_acc_46_nl[23:0];
  assign FpCmp_8U_23U_false_else_else_if_acc_46_itm_23_1 = readslicef_24_1_23((FpCmp_8U_23U_false_else_else_if_acc_46_nl));
  assign nl_FpCmp_8U_23U_false_else_if_acc_46_nl = ({1'b1 , (AluIn_data_sva_501[510:503])})
      + conv_u2u_8_9({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_9) ,
      (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_9)}) + 9'b1;
  assign FpCmp_8U_23U_false_else_if_acc_46_nl = nl_FpCmp_8U_23U_false_else_if_acc_46_nl[8:0];
  assign FpCmp_8U_23U_false_else_if_acc_46_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_false_else_if_acc_46_nl));
  assign nl_FpCmp_8U_23U_true_if_acc_16_nl = ({1'b1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_mx0w0
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w0}) + conv_u2u_8_9(~
      (AluIn_data_sva_1[30:23])) + 9'b1;
  assign FpCmp_8U_23U_true_if_acc_16_nl = nl_FpCmp_8U_23U_true_if_acc_16_nl[8:0];
  assign FpCmp_8U_23U_true_if_acc_16_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_true_if_acc_16_nl));
  assign nl_FpCmp_8U_23U_true_if_acc_18_nl = ({1'b1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_mx0w0
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w0}) + conv_u2u_8_9(~
      (AluIn_data_sva_1[62:55])) + 9'b1;
  assign FpCmp_8U_23U_true_if_acc_18_nl = nl_FpCmp_8U_23U_true_if_acc_18_nl[8:0];
  assign FpCmp_8U_23U_true_if_acc_18_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_true_if_acc_18_nl));
  assign nl_FpCmp_8U_23U_true_if_acc_20_nl = ({1'b1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_mx0w0
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w0}) + conv_u2u_8_9(~
      (AluIn_data_sva_1[94:87])) + 9'b1;
  assign FpCmp_8U_23U_true_if_acc_20_nl = nl_FpCmp_8U_23U_true_if_acc_20_nl[8:0];
  assign FpCmp_8U_23U_true_if_acc_20_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_true_if_acc_20_nl));
  assign nl_FpCmp_8U_23U_true_if_acc_22_nl = ({1'b1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_mx0w0
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3_mx0w0}) + conv_u2u_8_9(~
      (AluIn_data_sva_1[126:119])) + 9'b1;
  assign FpCmp_8U_23U_true_if_acc_22_nl = nl_FpCmp_8U_23U_true_if_acc_22_nl[8:0];
  assign FpCmp_8U_23U_true_if_acc_22_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_true_if_acc_22_nl));
  assign nl_FpCmp_8U_23U_true_if_acc_24_nl = ({1'b1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_mx0w0
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3_mx0w0}) + conv_u2u_8_9(~
      (AluIn_data_sva_1[158:151])) + 9'b1;
  assign FpCmp_8U_23U_true_if_acc_24_nl = nl_FpCmp_8U_23U_true_if_acc_24_nl[8:0];
  assign FpCmp_8U_23U_true_if_acc_24_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_true_if_acc_24_nl));
  assign nl_FpCmp_8U_23U_true_if_acc_26_nl = ({1'b1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_mx0w0
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3_mx0w0}) + conv_u2u_8_9(~
      (AluIn_data_sva_1[190:183])) + 9'b1;
  assign FpCmp_8U_23U_true_if_acc_26_nl = nl_FpCmp_8U_23U_true_if_acc_26_nl[8:0];
  assign FpCmp_8U_23U_true_if_acc_26_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_true_if_acc_26_nl));
  assign nl_FpCmp_8U_23U_true_if_acc_28_nl = ({1'b1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_mx0w0
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3_mx0w0}) + conv_u2u_8_9(~
      (AluIn_data_sva_1[222:215])) + 9'b1;
  assign FpCmp_8U_23U_true_if_acc_28_nl = nl_FpCmp_8U_23U_true_if_acc_28_nl[8:0];
  assign FpCmp_8U_23U_true_if_acc_28_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_true_if_acc_28_nl));
  assign nl_FpCmp_8U_23U_true_if_acc_30_nl = ({1'b1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_mx0w0
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3_mx0w0}) + conv_u2u_8_9(~
      (AluIn_data_sva_1[254:247])) + 9'b1;
  assign FpCmp_8U_23U_true_if_acc_30_nl = nl_FpCmp_8U_23U_true_if_acc_30_nl[8:0];
  assign FpCmp_8U_23U_true_if_acc_30_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_true_if_acc_30_nl));
  assign nl_FpCmp_8U_23U_true_if_acc_32_nl = ({1'b1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_mx0w0
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3_mx0w0}) + conv_u2u_8_9(~
      (AluIn_data_sva_1[286:279])) + 9'b1;
  assign FpCmp_8U_23U_true_if_acc_32_nl = nl_FpCmp_8U_23U_true_if_acc_32_nl[8:0];
  assign FpCmp_8U_23U_true_if_acc_32_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_true_if_acc_32_nl));
  assign nl_FpCmp_8U_23U_true_if_acc_34_nl = ({1'b1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_mx0w0
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3_mx0w0}) + conv_u2u_8_9(~
      (AluIn_data_sva_1[318:311])) + 9'b1;
  assign FpCmp_8U_23U_true_if_acc_34_nl = nl_FpCmp_8U_23U_true_if_acc_34_nl[8:0];
  assign FpCmp_8U_23U_true_if_acc_34_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_true_if_acc_34_nl));
  assign nl_FpCmp_8U_23U_true_if_acc_36_nl = ({1'b1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_mx0w0
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3_mx0w0}) + conv_u2u_8_9(~
      (AluIn_data_sva_1[350:343])) + 9'b1;
  assign FpCmp_8U_23U_true_if_acc_36_nl = nl_FpCmp_8U_23U_true_if_acc_36_nl[8:0];
  assign FpCmp_8U_23U_true_if_acc_36_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_true_if_acc_36_nl));
  assign nl_FpCmp_8U_23U_true_if_acc_38_nl = ({1'b1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_mx0w0
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3_mx0w0}) + conv_u2u_8_9(~
      (AluIn_data_sva_1[382:375])) + 9'b1;
  assign FpCmp_8U_23U_true_if_acc_38_nl = nl_FpCmp_8U_23U_true_if_acc_38_nl[8:0];
  assign FpCmp_8U_23U_true_if_acc_38_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_true_if_acc_38_nl));
  assign nl_FpCmp_8U_23U_true_if_acc_40_nl = ({1'b1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_mx0w0
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3_mx0w0}) + conv_u2u_8_9(~
      (AluIn_data_sva_1[414:407])) + 9'b1;
  assign FpCmp_8U_23U_true_if_acc_40_nl = nl_FpCmp_8U_23U_true_if_acc_40_nl[8:0];
  assign FpCmp_8U_23U_true_if_acc_40_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_true_if_acc_40_nl));
  assign nl_FpCmp_8U_23U_true_if_acc_42_nl = ({1'b1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_mx0w0
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3_mx0w0}) + conv_u2u_8_9(~
      (AluIn_data_sva_1[446:439])) + 9'b1;
  assign FpCmp_8U_23U_true_if_acc_42_nl = nl_FpCmp_8U_23U_true_if_acc_42_nl[8:0];
  assign FpCmp_8U_23U_true_if_acc_42_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_true_if_acc_42_nl));
  assign nl_FpCmp_8U_23U_true_if_acc_44_nl = ({1'b1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_mx0w0
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3_mx0w0}) + conv_u2u_8_9(~
      (AluIn_data_sva_1[478:471])) + 9'b1;
  assign FpCmp_8U_23U_true_if_acc_44_nl = nl_FpCmp_8U_23U_true_if_acc_44_nl[8:0];
  assign FpCmp_8U_23U_true_if_acc_44_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_true_if_acc_44_nl));
  assign nl_FpCmp_8U_23U_true_if_acc_46_nl = ({1'b1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_mx0w0
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w0}) + conv_u2u_8_9(~
      (AluIn_data_sva_1[510:503])) + 9'b1;
  assign FpCmp_8U_23U_true_if_acc_46_nl = nl_FpCmp_8U_23U_true_if_acc_46_nl[8:0];
  assign FpCmp_8U_23U_true_if_acc_46_itm_8_1 = readslicef_9_1_8((FpCmp_8U_23U_true_if_acc_46_nl));
  assign nl_alu_loop_op_1_FpNormalize_8U_49U_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_qr_2_lpi_1_dfm_5_7_4_1)
      , (~ FpAdd_8U_23U_qr_2_lpi_1_dfm_5_3_0_1)}) + conv_u2s_6_9(IntLeadZero_49U_leading_sign_49_0_rtn_1_sva_2)
      + 9'b1;
  assign alu_loop_op_1_FpNormalize_8U_49U_acc_nl = nl_alu_loop_op_1_FpNormalize_8U_49U_acc_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_33 = FpNormalize_8U_49U_if_or_itm_2 & (readslicef_9_1_8((alu_loop_op_1_FpNormalize_8U_49U_acc_nl)));
  assign FpAdd_8U_23U_asn_256 = (~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_2)
      & (FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49]);
  assign FpAdd_8U_23U_asn_258 = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_2
      & (FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49]);
  assign nl_alu_loop_op_2_FpNormalize_8U_49U_acc_1_nl = ({1'b1 , (~ FpAdd_8U_23U_qr_3_lpi_1_dfm_5_7_4_1)
      , (~ FpAdd_8U_23U_qr_3_lpi_1_dfm_5_3_0_1)}) + conv_u2s_6_9(IntLeadZero_49U_leading_sign_49_0_rtn_2_sva_2)
      + 9'b1;
  assign alu_loop_op_2_FpNormalize_8U_49U_acc_1_nl = nl_alu_loop_op_2_FpNormalize_8U_49U_acc_1_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_35 = FpNormalize_8U_49U_if_or_1_itm_2 & (readslicef_9_1_8((alu_loop_op_2_FpNormalize_8U_49U_acc_1_nl)));
  assign FpAdd_8U_23U_asn_260 = (~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_2)
      & (FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49]);
  assign FpAdd_8U_23U_asn_262 = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_2
      & (FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49]);
  assign nl_alu_loop_op_3_FpNormalize_8U_49U_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_qr_4_lpi_1_dfm_5_7_4_1)
      , (~ FpAdd_8U_23U_qr_4_lpi_1_dfm_5_3_0_1)}) + conv_u2s_6_9(IntLeadZero_49U_leading_sign_49_0_rtn_3_sva_2)
      + 9'b1;
  assign alu_loop_op_3_FpNormalize_8U_49U_acc_nl = nl_alu_loop_op_3_FpNormalize_8U_49U_acc_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_37 = FpNormalize_8U_49U_if_or_2_itm_2 & (readslicef_9_1_8((alu_loop_op_3_FpNormalize_8U_49U_acc_nl)));
  assign FpAdd_8U_23U_asn_264 = (~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_2)
      & (FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49]);
  assign FpAdd_8U_23U_asn_266 = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_2
      & (FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49]);
  assign nl_alu_loop_op_4_FpNormalize_8U_49U_acc_1_nl = ({1'b1 , (~ FpAdd_8U_23U_qr_5_lpi_1_dfm_5_7_4_1)
      , (~ FpAdd_8U_23U_qr_5_lpi_1_dfm_5_3_0_1)}) + conv_u2s_6_9(IntLeadZero_49U_leading_sign_49_0_rtn_4_sva_2)
      + 9'b1;
  assign alu_loop_op_4_FpNormalize_8U_49U_acc_1_nl = nl_alu_loop_op_4_FpNormalize_8U_49U_acc_1_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_39 = FpNormalize_8U_49U_if_or_3_itm_2 & (readslicef_9_1_8((alu_loop_op_4_FpNormalize_8U_49U_acc_1_nl)));
  assign FpAdd_8U_23U_asn_268 = (~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_4_sva_2)
      & (FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_5[49]);
  assign FpAdd_8U_23U_asn_270 = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_4_sva_2
      & (FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_5[49]);
  assign nl_alu_loop_op_5_FpNormalize_8U_49U_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_qr_6_lpi_1_dfm_5_7_4_1)
      , (~ FpAdd_8U_23U_qr_6_lpi_1_dfm_5_3_0_1)}) + conv_u2s_6_9(IntLeadZero_49U_leading_sign_49_0_rtn_5_sva_2)
      + 9'b1;
  assign alu_loop_op_5_FpNormalize_8U_49U_acc_nl = nl_alu_loop_op_5_FpNormalize_8U_49U_acc_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_41 = FpNormalize_8U_49U_if_or_4_itm_2 & (readslicef_9_1_8((alu_loop_op_5_FpNormalize_8U_49U_acc_nl)));
  assign FpAdd_8U_23U_asn_272 = (~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_5_sva_2)
      & (FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_5[49]);
  assign FpAdd_8U_23U_asn_274 = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_5_sva_2
      & (FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_5[49]);
  assign nl_alu_loop_op_6_FpNormalize_8U_49U_acc_1_nl = ({1'b1 , (~ FpAdd_8U_23U_qr_7_lpi_1_dfm_5_7_4_1)
      , (~ FpAdd_8U_23U_qr_7_lpi_1_dfm_5_3_0_1)}) + conv_u2s_6_9(IntLeadZero_49U_leading_sign_49_0_rtn_6_sva_2)
      + 9'b1;
  assign alu_loop_op_6_FpNormalize_8U_49U_acc_1_nl = nl_alu_loop_op_6_FpNormalize_8U_49U_acc_1_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_43 = FpNormalize_8U_49U_if_or_5_itm_2 & (readslicef_9_1_8((alu_loop_op_6_FpNormalize_8U_49U_acc_1_nl)));
  assign FpAdd_8U_23U_asn_276 = (~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_6_sva_2)
      & (FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_5[49]);
  assign FpAdd_8U_23U_asn_278 = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_6_sva_2
      & (FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_5[49]);
  assign nl_alu_loop_op_7_FpNormalize_8U_49U_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_qr_8_lpi_1_dfm_5_7_4_1)
      , (~ FpAdd_8U_23U_qr_8_lpi_1_dfm_5_3_0_1)}) + conv_u2s_6_9(IntLeadZero_49U_leading_sign_49_0_rtn_7_sva_2)
      + 9'b1;
  assign alu_loop_op_7_FpNormalize_8U_49U_acc_nl = nl_alu_loop_op_7_FpNormalize_8U_49U_acc_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_45 = FpNormalize_8U_49U_if_or_6_itm_2 & (readslicef_9_1_8((alu_loop_op_7_FpNormalize_8U_49U_acc_nl)));
  assign FpAdd_8U_23U_asn_280 = (~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_7_sva_2)
      & (FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_5[49]);
  assign FpAdd_8U_23U_asn_282 = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_7_sva_2
      & (FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_5[49]);
  assign nl_alu_loop_op_8_FpNormalize_8U_49U_acc_1_nl = ({1'b1 , (~ FpAdd_8U_23U_qr_9_lpi_1_dfm_5_7_4_1)
      , (~ FpAdd_8U_23U_qr_9_lpi_1_dfm_5_3_0_1)}) + conv_u2s_6_9(IntLeadZero_49U_leading_sign_49_0_rtn_8_sva_2)
      + 9'b1;
  assign alu_loop_op_8_FpNormalize_8U_49U_acc_1_nl = nl_alu_loop_op_8_FpNormalize_8U_49U_acc_1_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_47 = FpNormalize_8U_49U_if_or_7_itm_2 & (readslicef_9_1_8((alu_loop_op_8_FpNormalize_8U_49U_acc_1_nl)));
  assign FpAdd_8U_23U_asn_284 = (~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_8_sva_2)
      & (FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_5[49]);
  assign FpAdd_8U_23U_asn_286 = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_8_sva_2
      & (FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_5[49]);
  assign nl_alu_loop_op_9_FpNormalize_8U_49U_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_qr_10_lpi_1_dfm_5_7_4_1)
      , (~ FpAdd_8U_23U_qr_10_lpi_1_dfm_5_3_0_1)}) + conv_u2s_6_9(IntLeadZero_49U_leading_sign_49_0_rtn_9_sva_2)
      + 9'b1;
  assign alu_loop_op_9_FpNormalize_8U_49U_acc_nl = nl_alu_loop_op_9_FpNormalize_8U_49U_acc_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_49 = FpNormalize_8U_49U_if_or_8_itm_2 & (readslicef_9_1_8((alu_loop_op_9_FpNormalize_8U_49U_acc_nl)));
  assign FpAdd_8U_23U_asn_288 = (~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_9_sva_2)
      & (FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_5[49]);
  assign FpAdd_8U_23U_asn_290 = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_9_sva_2
      & (FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_5[49]);
  assign nl_alu_loop_op_10_FpNormalize_8U_49U_acc_1_nl = ({1'b1 , (~ FpAdd_8U_23U_qr_11_lpi_1_dfm_5_7_4_1)
      , (~ FpAdd_8U_23U_qr_11_lpi_1_dfm_5_3_0_1)}) + conv_u2s_6_9(IntLeadZero_49U_leading_sign_49_0_rtn_10_sva_2)
      + 9'b1;
  assign alu_loop_op_10_FpNormalize_8U_49U_acc_1_nl = nl_alu_loop_op_10_FpNormalize_8U_49U_acc_1_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_51 = FpNormalize_8U_49U_if_or_9_itm_2 & (readslicef_9_1_8((alu_loop_op_10_FpNormalize_8U_49U_acc_1_nl)));
  assign FpAdd_8U_23U_asn_292 = (~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_10_sva_2)
      & (FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_5[49]);
  assign FpAdd_8U_23U_asn_294 = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_10_sva_2
      & (FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_5[49]);
  assign nl_alu_loop_op_11_FpNormalize_8U_49U_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_qr_12_lpi_1_dfm_5_7_4_1)
      , (~ FpAdd_8U_23U_qr_12_lpi_1_dfm_5_3_0_1)}) + conv_u2s_6_9(IntLeadZero_49U_leading_sign_49_0_rtn_11_sva_2)
      + 9'b1;
  assign alu_loop_op_11_FpNormalize_8U_49U_acc_nl = nl_alu_loop_op_11_FpNormalize_8U_49U_acc_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_53 = FpNormalize_8U_49U_if_or_10_itm_2 & (readslicef_9_1_8((alu_loop_op_11_FpNormalize_8U_49U_acc_nl)));
  assign FpAdd_8U_23U_asn_296 = (~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_11_sva_2)
      & (FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_5[49]);
  assign FpAdd_8U_23U_asn_298 = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_11_sva_2
      & (FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_5[49]);
  assign nl_alu_loop_op_12_FpNormalize_8U_49U_acc_1_nl = ({1'b1 , (~ FpAdd_8U_23U_qr_13_lpi_1_dfm_5_7_4_1)
      , (~ FpAdd_8U_23U_qr_13_lpi_1_dfm_5_3_0_1)}) + conv_u2s_6_9(IntLeadZero_49U_leading_sign_49_0_rtn_12_sva_2)
      + 9'b1;
  assign alu_loop_op_12_FpNormalize_8U_49U_acc_1_nl = nl_alu_loop_op_12_FpNormalize_8U_49U_acc_1_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_55 = FpNormalize_8U_49U_if_or_11_itm_2 & (readslicef_9_1_8((alu_loop_op_12_FpNormalize_8U_49U_acc_1_nl)));
  assign FpAdd_8U_23U_asn_300 = (~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_12_sva_2)
      & (FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_5[49]);
  assign FpAdd_8U_23U_asn_302 = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_12_sva_2
      & (FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_5[49]);
  assign nl_alu_loop_op_13_FpNormalize_8U_49U_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_qr_14_lpi_1_dfm_5_7_4_1)
      , (~ FpAdd_8U_23U_qr_14_lpi_1_dfm_5_3_0_1)}) + conv_u2s_6_9(IntLeadZero_49U_leading_sign_49_0_rtn_13_sva_2)
      + 9'b1;
  assign alu_loop_op_13_FpNormalize_8U_49U_acc_nl = nl_alu_loop_op_13_FpNormalize_8U_49U_acc_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_57 = FpNormalize_8U_49U_if_or_12_itm_2 & (readslicef_9_1_8((alu_loop_op_13_FpNormalize_8U_49U_acc_nl)));
  assign FpAdd_8U_23U_asn_304 = (~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_13_sva_2)
      & (FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_5[49]);
  assign FpAdd_8U_23U_asn_306 = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_13_sva_2
      & (FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_5[49]);
  assign nl_alu_loop_op_14_FpNormalize_8U_49U_acc_1_nl = ({1'b1 , (~ FpAdd_8U_23U_qr_15_lpi_1_dfm_5_7_4_1)
      , (~ FpAdd_8U_23U_qr_15_lpi_1_dfm_5_3_0_1)}) + conv_u2s_6_9(IntLeadZero_49U_leading_sign_49_0_rtn_14_sva_2)
      + 9'b1;
  assign alu_loop_op_14_FpNormalize_8U_49U_acc_1_nl = nl_alu_loop_op_14_FpNormalize_8U_49U_acc_1_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_59 = FpNormalize_8U_49U_if_or_13_itm_2 & (readslicef_9_1_8((alu_loop_op_14_FpNormalize_8U_49U_acc_1_nl)));
  assign FpAdd_8U_23U_asn_308 = (~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_14_sva_2)
      & (FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_5[49]);
  assign FpAdd_8U_23U_asn_310 = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_14_sva_2
      & (FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_5[49]);
  assign nl_alu_loop_op_15_FpNormalize_8U_49U_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_qr_16_lpi_1_dfm_5_7_4_1)
      , (~ FpAdd_8U_23U_qr_16_lpi_1_dfm_5_3_0_1)}) + conv_u2s_6_9(IntLeadZero_49U_leading_sign_49_0_rtn_15_sva_2)
      + 9'b1;
  assign alu_loop_op_15_FpNormalize_8U_49U_acc_nl = nl_alu_loop_op_15_FpNormalize_8U_49U_acc_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_61 = FpNormalize_8U_49U_if_or_14_itm_2 & (readslicef_9_1_8((alu_loop_op_15_FpNormalize_8U_49U_acc_nl)));
  assign FpAdd_8U_23U_asn_312 = (~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_15_sva_2)
      & (FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_5[49]);
  assign FpAdd_8U_23U_asn_314 = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_15_sva_2
      & (FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_5[49]);
  assign nl_alu_loop_op_16_FpNormalize_8U_49U_acc_1_nl = ({1'b1 , (~ FpAdd_8U_23U_qr_lpi_1_dfm_5_7_4_1)
      , (~ FpAdd_8U_23U_qr_lpi_1_dfm_5_3_0_1)}) + conv_u2s_6_9(IntLeadZero_49U_leading_sign_49_0_rtn_sva_2)
      + 9'b1;
  assign alu_loop_op_16_FpNormalize_8U_49U_acc_1_nl = nl_alu_loop_op_16_FpNormalize_8U_49U_acc_1_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_63 = FpNormalize_8U_49U_if_or_15_itm_2 & (readslicef_9_1_8((alu_loop_op_16_FpNormalize_8U_49U_acc_1_nl)));
  assign FpAdd_8U_23U_asn_316 = (~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_2)
      & (FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49]);
  assign FpAdd_8U_23U_asn_318 = FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_2
      & (FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49]);
  assign asn_1837 = alu_loop_op_else_nor_tmp_82 & and_1_m1c;
  assign else_mux_47_tmp = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]), (chn_alu_op_rsci_d_mxwt[254:250]),
      cfg_alu_src_1_sva_st);
  assign else_mux_44_tmp = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]), (chn_alu_op_rsci_d_mxwt[238:234]),
      cfg_alu_src_1_sva_st);
  assign else_mux_41_tmp = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]), (chn_alu_op_rsci_d_mxwt[222:218]),
      cfg_alu_src_1_sva_st);
  assign else_mux_38_tmp = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]), (chn_alu_op_rsci_d_mxwt[206:202]),
      cfg_alu_src_1_sva_st);
  assign else_mux_35_tmp = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]), (chn_alu_op_rsci_d_mxwt[190:186]),
      cfg_alu_src_1_sva_st);
  assign else_mux_32_tmp = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]), (chn_alu_op_rsci_d_mxwt[174:170]),
      cfg_alu_src_1_sva_st);
  assign else_mux_29_tmp = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]), (chn_alu_op_rsci_d_mxwt[158:154]),
      cfg_alu_src_1_sva_st);
  assign else_mux_26_tmp = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]), (chn_alu_op_rsci_d_mxwt[142:138]),
      cfg_alu_src_1_sva_st);
  assign else_mux_23_tmp = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]), (chn_alu_op_rsci_d_mxwt[126:122]),
      cfg_alu_src_1_sva_st);
  assign else_mux_20_tmp = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]), (chn_alu_op_rsci_d_mxwt[110:106]),
      cfg_alu_src_1_sva_st);
  assign else_mux_17_tmp = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]), (chn_alu_op_rsci_d_mxwt[94:90]),
      cfg_alu_src_1_sva_st);
  assign else_mux_14_tmp = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]), (chn_alu_op_rsci_d_mxwt[78:74]),
      cfg_alu_src_1_sva_st);
  assign else_mux_11_tmp = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]), (chn_alu_op_rsci_d_mxwt[62:58]),
      cfg_alu_src_1_sva_st);
  assign else_mux_8_tmp = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]), (chn_alu_op_rsci_d_mxwt[46:42]),
      cfg_alu_src_1_sva_st);
  assign else_mux_5_tmp = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]), (chn_alu_op_rsci_d_mxwt[30:26]),
      cfg_alu_src_1_sva_st);
  assign else_mux_2_tmp = MUX_v_5_2_2((cfg_alu_op_1_sva_1[14:10]), (chn_alu_op_rsci_d_mxwt[14:10]),
      cfg_alu_src_1_sva_st);
  assign and_89_tmp = main_stage_v_1 & or_4_cse & or_5_cse & or_6_cse & or_7_cse
      & or_8_cse & or_9_cse & or_cse_2;
  assign FpAdd_8U_23U_mux_242_tmp_49 = MUX_s_1_2_2((FpAdd_8U_23U_asn_mx1w1[49]),
      (FpAdd_8U_23U_int_mant_p1_sva[49]), reg_alu_loop_op_16_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse);
  assign FpAdd_8U_23U_mux_226_tmp_49 = MUX_s_1_2_2((FpAdd_8U_23U_asn_34_mx1w1[49]),
      (FpAdd_8U_23U_int_mant_p1_15_sva[49]), reg_alu_loop_op_15_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse);
  assign FpAdd_8U_23U_mux_210_tmp_49 = MUX_s_1_2_2((FpAdd_8U_23U_asn_37_mx1w1[49]),
      (FpAdd_8U_23U_int_mant_p1_14_sva[49]), reg_alu_loop_op_14_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse);
  assign FpAdd_8U_23U_mux_194_tmp_49 = MUX_s_1_2_2((FpAdd_8U_23U_asn_40_mx1w1[49]),
      (FpAdd_8U_23U_int_mant_p1_13_sva[49]), reg_alu_loop_op_13_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse);
  assign FpAdd_8U_23U_mux_178_tmp_49 = MUX_s_1_2_2((FpAdd_8U_23U_asn_43_mx1w1[49]),
      (FpAdd_8U_23U_int_mant_p1_12_sva[49]), reg_alu_loop_op_12_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse);
  assign FpAdd_8U_23U_mux_162_tmp_49 = MUX_s_1_2_2((FpAdd_8U_23U_asn_46_mx1w1[49]),
      (FpAdd_8U_23U_int_mant_p1_11_sva[49]), reg_alu_loop_op_11_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse);
  assign FpAdd_8U_23U_mux_146_tmp_49 = MUX_s_1_2_2((FpAdd_8U_23U_asn_49_mx1w1[49]),
      (FpAdd_8U_23U_int_mant_p1_10_sva[49]), reg_alu_loop_op_10_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse);
  assign FpAdd_8U_23U_mux_130_tmp_49 = MUX_s_1_2_2((FpAdd_8U_23U_asn_52_mx1w1[49]),
      (FpAdd_8U_23U_int_mant_p1_9_sva[49]), reg_alu_loop_op_9_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse);
  assign FpAdd_8U_23U_mux_114_tmp_49 = MUX_s_1_2_2((FpAdd_8U_23U_asn_55_mx1w1[49]),
      (FpAdd_8U_23U_int_mant_p1_8_sva[49]), reg_alu_loop_op_8_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse);
  assign FpAdd_8U_23U_mux_98_tmp_49 = MUX_s_1_2_2((FpAdd_8U_23U_asn_58_mx1w1[49]),
      (FpAdd_8U_23U_int_mant_p1_7_sva[49]), reg_alu_loop_op_7_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse);
  assign FpAdd_8U_23U_mux_82_tmp_49 = MUX_s_1_2_2((FpAdd_8U_23U_asn_61_mx1w1[49]),
      (FpAdd_8U_23U_int_mant_p1_6_sva[49]), reg_alu_loop_op_6_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse);
  assign FpAdd_8U_23U_mux_66_tmp_49 = MUX_s_1_2_2((FpAdd_8U_23U_asn_64_mx1w1[49]),
      (FpAdd_8U_23U_int_mant_p1_5_sva[49]), reg_alu_loop_op_5_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse);
  assign FpAdd_8U_23U_mux_50_tmp_49 = MUX_s_1_2_2((FpAdd_8U_23U_asn_67_mx1w1[49]),
      (FpAdd_8U_23U_int_mant_p1_4_sva[49]), reg_alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse);
  assign FpAdd_8U_23U_mux_34_tmp_49 = MUX_s_1_2_2((FpAdd_8U_23U_asn_70_mx1w1[49]),
      (FpAdd_8U_23U_int_mant_p1_3_sva[49]), reg_alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse);
  assign FpAdd_8U_23U_mux_18_tmp_49 = MUX_s_1_2_2((FpAdd_8U_23U_asn_73_mx1w1[49]),
      (FpAdd_8U_23U_int_mant_p1_2_sva[49]), reg_alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse);
  assign FpAdd_8U_23U_mux_2_tmp_49 = MUX_s_1_2_2((FpAdd_8U_23U_asn_76_mx1w1[49]),
      (FpAdd_8U_23U_int_mant_p1_1_sva[49]), reg_alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse);
  assign nl_alu_loop_op_16_else_if_acc_1_nl = conv_s2u_32_33({IntShiftLeft_16U_6U_32U_return_31_sva_2
      , IntShiftLeft_16U_6U_32U_return_30_1_sva_2 , IntShiftLeft_16U_6U_32U_return_0_sva_2})
      - conv_s2u_32_33(AluIn_data_sva_501[511:480]);
  assign alu_loop_op_16_else_if_acc_1_nl = nl_alu_loop_op_16_else_if_acc_1_nl[32:0];
  assign alu_loop_op_16_else_if_acc_1_itm_32_1 = readslicef_33_1_32((alu_loop_op_16_else_if_acc_1_nl));
  assign nl_alu_loop_op_16_else_else_if_acc_1_nl = conv_s2u_32_33(AluIn_data_sva_501[511:480])
      + conv_s2u_32_33({(~ IntShiftLeft_16U_6U_32U_return_31_sva_2) , (~ IntShiftLeft_16U_6U_32U_return_30_1_sva_2)
      , (~ IntShiftLeft_16U_6U_32U_return_0_sva_2)}) + 33'b1;
  assign alu_loop_op_16_else_else_if_acc_1_nl = nl_alu_loop_op_16_else_else_if_acc_1_nl[32:0];
  assign alu_loop_op_16_else_else_if_acc_1_itm_32_1 = readslicef_33_1_32((alu_loop_op_16_else_else_if_acc_1_nl));
  assign nl_alu_loop_op_15_else_if_acc_nl = conv_s2u_32_33({IntShiftLeft_16U_6U_32U_return_31_15_sva_2
      , IntShiftLeft_16U_6U_32U_return_30_1_15_sva_2 , IntShiftLeft_16U_6U_32U_return_0_15_sva_2})
      - conv_s2u_32_33(AluIn_data_sva_501[479:448]);
  assign alu_loop_op_15_else_if_acc_nl = nl_alu_loop_op_15_else_if_acc_nl[32:0];
  assign alu_loop_op_15_else_if_acc_itm_32_1 = readslicef_33_1_32((alu_loop_op_15_else_if_acc_nl));
  assign nl_alu_loop_op_15_else_else_if_acc_nl = conv_s2u_32_33(AluIn_data_sva_501[479:448])
      + conv_s2u_32_33({(~ IntShiftLeft_16U_6U_32U_return_31_15_sva_2) , (~ IntShiftLeft_16U_6U_32U_return_30_1_15_sva_2)
      , (~ IntShiftLeft_16U_6U_32U_return_0_15_sva_2)}) + 33'b1;
  assign alu_loop_op_15_else_else_if_acc_nl = nl_alu_loop_op_15_else_else_if_acc_nl[32:0];
  assign alu_loop_op_15_else_else_if_acc_itm_32_1 = readslicef_33_1_32((alu_loop_op_15_else_else_if_acc_nl));
  assign nl_alu_loop_op_14_else_if_acc_1_nl = conv_s2u_32_33({IntShiftLeft_16U_6U_32U_return_31_14_sva_2
      , IntShiftLeft_16U_6U_32U_return_30_1_14_sva_2 , IntShiftLeft_16U_6U_32U_return_0_14_sva_2})
      - conv_s2u_32_33(AluIn_data_sva_501[447:416]);
  assign alu_loop_op_14_else_if_acc_1_nl = nl_alu_loop_op_14_else_if_acc_1_nl[32:0];
  assign alu_loop_op_14_else_if_acc_1_itm_32_1 = readslicef_33_1_32((alu_loop_op_14_else_if_acc_1_nl));
  assign nl_alu_loop_op_14_else_else_if_acc_1_nl = conv_s2u_32_33(AluIn_data_sva_501[447:416])
      + conv_s2u_32_33({(~ IntShiftLeft_16U_6U_32U_return_31_14_sva_2) , (~ IntShiftLeft_16U_6U_32U_return_30_1_14_sva_2)
      , (~ IntShiftLeft_16U_6U_32U_return_0_14_sva_2)}) + 33'b1;
  assign alu_loop_op_14_else_else_if_acc_1_nl = nl_alu_loop_op_14_else_else_if_acc_1_nl[32:0];
  assign alu_loop_op_14_else_else_if_acc_1_itm_32_1 = readslicef_33_1_32((alu_loop_op_14_else_else_if_acc_1_nl));
  assign nl_alu_loop_op_13_else_if_acc_nl = conv_s2u_32_33({IntShiftLeft_16U_6U_32U_return_31_13_sva_2
      , IntShiftLeft_16U_6U_32U_return_30_1_13_sva_2 , IntShiftLeft_16U_6U_32U_return_0_13_sva_2})
      - conv_s2u_32_33(AluIn_data_sva_501[415:384]);
  assign alu_loop_op_13_else_if_acc_nl = nl_alu_loop_op_13_else_if_acc_nl[32:0];
  assign alu_loop_op_13_else_if_acc_itm_32_1 = readslicef_33_1_32((alu_loop_op_13_else_if_acc_nl));
  assign nl_alu_loop_op_13_else_else_if_acc_nl = conv_s2u_32_33(AluIn_data_sva_501[415:384])
      + conv_s2u_32_33({(~ IntShiftLeft_16U_6U_32U_return_31_13_sva_2) , (~ IntShiftLeft_16U_6U_32U_return_30_1_13_sva_2)
      , (~ IntShiftLeft_16U_6U_32U_return_0_13_sva_2)}) + 33'b1;
  assign alu_loop_op_13_else_else_if_acc_nl = nl_alu_loop_op_13_else_else_if_acc_nl[32:0];
  assign alu_loop_op_13_else_else_if_acc_itm_32_1 = readslicef_33_1_32((alu_loop_op_13_else_else_if_acc_nl));
  assign nl_alu_loop_op_12_else_if_acc_1_nl = conv_s2u_32_33({IntShiftLeft_16U_6U_32U_return_31_12_sva_2
      , IntShiftLeft_16U_6U_32U_return_30_1_12_sva_2 , IntShiftLeft_16U_6U_32U_return_0_12_sva_2})
      - conv_s2u_32_33(AluIn_data_sva_501[383:352]);
  assign alu_loop_op_12_else_if_acc_1_nl = nl_alu_loop_op_12_else_if_acc_1_nl[32:0];
  assign alu_loop_op_12_else_if_acc_1_itm_32_1 = readslicef_33_1_32((alu_loop_op_12_else_if_acc_1_nl));
  assign nl_alu_loop_op_12_else_else_if_acc_1_nl = conv_s2u_32_33(AluIn_data_sva_501[383:352])
      + conv_s2u_32_33({(~ IntShiftLeft_16U_6U_32U_return_31_12_sva_2) , (~ IntShiftLeft_16U_6U_32U_return_30_1_12_sva_2)
      , (~ IntShiftLeft_16U_6U_32U_return_0_12_sva_2)}) + 33'b1;
  assign alu_loop_op_12_else_else_if_acc_1_nl = nl_alu_loop_op_12_else_else_if_acc_1_nl[32:0];
  assign alu_loop_op_12_else_else_if_acc_1_itm_32_1 = readslicef_33_1_32((alu_loop_op_12_else_else_if_acc_1_nl));
  assign nl_alu_loop_op_11_else_if_acc_nl = conv_s2u_32_33({IntShiftLeft_16U_6U_32U_return_31_11_sva_2
      , IntShiftLeft_16U_6U_32U_return_30_1_11_sva_2 , IntShiftLeft_16U_6U_32U_return_0_11_sva_2})
      - conv_s2u_32_33(AluIn_data_sva_501[351:320]);
  assign alu_loop_op_11_else_if_acc_nl = nl_alu_loop_op_11_else_if_acc_nl[32:0];
  assign alu_loop_op_11_else_if_acc_itm_32_1 = readslicef_33_1_32((alu_loop_op_11_else_if_acc_nl));
  assign nl_alu_loop_op_11_else_else_if_acc_nl = conv_s2u_32_33(AluIn_data_sva_501[351:320])
      + conv_s2u_32_33({(~ IntShiftLeft_16U_6U_32U_return_31_11_sva_2) , (~ IntShiftLeft_16U_6U_32U_return_30_1_11_sva_2)
      , (~ IntShiftLeft_16U_6U_32U_return_0_11_sva_2)}) + 33'b1;
  assign alu_loop_op_11_else_else_if_acc_nl = nl_alu_loop_op_11_else_else_if_acc_nl[32:0];
  assign alu_loop_op_11_else_else_if_acc_itm_32_1 = readslicef_33_1_32((alu_loop_op_11_else_else_if_acc_nl));
  assign nl_alu_loop_op_10_else_if_acc_1_nl = conv_s2u_32_33({IntShiftLeft_16U_6U_32U_return_31_10_sva_2
      , IntShiftLeft_16U_6U_32U_return_30_1_10_sva_2 , IntShiftLeft_16U_6U_32U_return_0_10_sva_2})
      - conv_s2u_32_33(AluIn_data_sva_501[319:288]);
  assign alu_loop_op_10_else_if_acc_1_nl = nl_alu_loop_op_10_else_if_acc_1_nl[32:0];
  assign alu_loop_op_10_else_if_acc_1_itm_32_1 = readslicef_33_1_32((alu_loop_op_10_else_if_acc_1_nl));
  assign nl_alu_loop_op_10_else_else_if_acc_1_nl = conv_s2u_32_33(AluIn_data_sva_501[319:288])
      + conv_s2u_32_33({(~ IntShiftLeft_16U_6U_32U_return_31_10_sva_2) , (~ IntShiftLeft_16U_6U_32U_return_30_1_10_sva_2)
      , (~ IntShiftLeft_16U_6U_32U_return_0_10_sva_2)}) + 33'b1;
  assign alu_loop_op_10_else_else_if_acc_1_nl = nl_alu_loop_op_10_else_else_if_acc_1_nl[32:0];
  assign alu_loop_op_10_else_else_if_acc_1_itm_32_1 = readslicef_33_1_32((alu_loop_op_10_else_else_if_acc_1_nl));
  assign nl_alu_loop_op_9_else_if_acc_nl = conv_s2u_32_33({IntShiftLeft_16U_6U_32U_return_31_9_sva_2
      , IntShiftLeft_16U_6U_32U_return_30_1_9_sva_2 , IntShiftLeft_16U_6U_32U_return_0_9_sva_2})
      - conv_s2u_32_33(AluIn_data_sva_501[287:256]);
  assign alu_loop_op_9_else_if_acc_nl = nl_alu_loop_op_9_else_if_acc_nl[32:0];
  assign alu_loop_op_9_else_if_acc_itm_32_1 = readslicef_33_1_32((alu_loop_op_9_else_if_acc_nl));
  assign nl_alu_loop_op_9_else_else_if_acc_nl = conv_s2u_32_33(AluIn_data_sva_501[287:256])
      + conv_s2u_32_33({(~ IntShiftLeft_16U_6U_32U_return_31_9_sva_2) , (~ IntShiftLeft_16U_6U_32U_return_30_1_9_sva_2)
      , (~ IntShiftLeft_16U_6U_32U_return_0_9_sva_2)}) + 33'b1;
  assign alu_loop_op_9_else_else_if_acc_nl = nl_alu_loop_op_9_else_else_if_acc_nl[32:0];
  assign alu_loop_op_9_else_else_if_acc_itm_32_1 = readslicef_33_1_32((alu_loop_op_9_else_else_if_acc_nl));
  assign nl_alu_loop_op_8_else_if_acc_1_nl = conv_s2u_32_33({IntShiftLeft_16U_6U_32U_return_31_8_sva_2
      , IntShiftLeft_16U_6U_32U_return_30_1_8_sva_2 , IntShiftLeft_16U_6U_32U_return_0_8_sva_2})
      - conv_s2u_32_33(AluIn_data_sva_501[255:224]);
  assign alu_loop_op_8_else_if_acc_1_nl = nl_alu_loop_op_8_else_if_acc_1_nl[32:0];
  assign alu_loop_op_8_else_if_acc_1_itm_32_1 = readslicef_33_1_32((alu_loop_op_8_else_if_acc_1_nl));
  assign nl_alu_loop_op_8_else_else_if_acc_1_nl = conv_s2u_32_33(AluIn_data_sva_501[255:224])
      + conv_s2u_32_33({(~ IntShiftLeft_16U_6U_32U_return_31_8_sva_2) , (~ IntShiftLeft_16U_6U_32U_return_30_1_8_sva_2)
      , (~ IntShiftLeft_16U_6U_32U_return_0_8_sva_2)}) + 33'b1;
  assign alu_loop_op_8_else_else_if_acc_1_nl = nl_alu_loop_op_8_else_else_if_acc_1_nl[32:0];
  assign alu_loop_op_8_else_else_if_acc_1_itm_32_1 = readslicef_33_1_32((alu_loop_op_8_else_else_if_acc_1_nl));
  assign nl_alu_loop_op_7_else_if_acc_nl = conv_s2u_32_33({IntShiftLeft_16U_6U_32U_return_31_7_sva_2
      , IntShiftLeft_16U_6U_32U_return_30_1_7_sva_2 , IntShiftLeft_16U_6U_32U_return_0_7_sva_2})
      - conv_s2u_32_33(AluIn_data_sva_501[223:192]);
  assign alu_loop_op_7_else_if_acc_nl = nl_alu_loop_op_7_else_if_acc_nl[32:0];
  assign alu_loop_op_7_else_if_acc_itm_32_1 = readslicef_33_1_32((alu_loop_op_7_else_if_acc_nl));
  assign nl_alu_loop_op_7_else_else_if_acc_nl = conv_s2u_32_33(AluIn_data_sva_501[223:192])
      + conv_s2u_32_33({(~ IntShiftLeft_16U_6U_32U_return_31_7_sva_2) , (~ IntShiftLeft_16U_6U_32U_return_30_1_7_sva_2)
      , (~ IntShiftLeft_16U_6U_32U_return_0_7_sva_2)}) + 33'b1;
  assign alu_loop_op_7_else_else_if_acc_nl = nl_alu_loop_op_7_else_else_if_acc_nl[32:0];
  assign alu_loop_op_7_else_else_if_acc_itm_32_1 = readslicef_33_1_32((alu_loop_op_7_else_else_if_acc_nl));
  assign nl_alu_loop_op_6_else_if_acc_1_nl = conv_s2u_32_33({IntShiftLeft_16U_6U_32U_return_31_6_sva_2
      , IntShiftLeft_16U_6U_32U_return_30_1_6_sva_2 , IntShiftLeft_16U_6U_32U_return_0_6_sva_2})
      - conv_s2u_32_33(AluIn_data_sva_501[191:160]);
  assign alu_loop_op_6_else_if_acc_1_nl = nl_alu_loop_op_6_else_if_acc_1_nl[32:0];
  assign alu_loop_op_6_else_if_acc_1_itm_32_1 = readslicef_33_1_32((alu_loop_op_6_else_if_acc_1_nl));
  assign nl_alu_loop_op_6_else_else_if_acc_1_nl = conv_s2u_32_33(AluIn_data_sva_501[191:160])
      + conv_s2u_32_33({(~ IntShiftLeft_16U_6U_32U_return_31_6_sva_2) , (~ IntShiftLeft_16U_6U_32U_return_30_1_6_sva_2)
      , (~ IntShiftLeft_16U_6U_32U_return_0_6_sva_2)}) + 33'b1;
  assign alu_loop_op_6_else_else_if_acc_1_nl = nl_alu_loop_op_6_else_else_if_acc_1_nl[32:0];
  assign alu_loop_op_6_else_else_if_acc_1_itm_32_1 = readslicef_33_1_32((alu_loop_op_6_else_else_if_acc_1_nl));
  assign nl_alu_loop_op_5_else_if_acc_nl = conv_s2u_32_33({IntShiftLeft_16U_6U_32U_return_31_5_sva_2
      , IntShiftLeft_16U_6U_32U_return_30_1_5_sva_2 , IntShiftLeft_16U_6U_32U_return_0_5_sva_2})
      - conv_s2u_32_33(AluIn_data_sva_501[159:128]);
  assign alu_loop_op_5_else_if_acc_nl = nl_alu_loop_op_5_else_if_acc_nl[32:0];
  assign alu_loop_op_5_else_if_acc_itm_32_1 = readslicef_33_1_32((alu_loop_op_5_else_if_acc_nl));
  assign nl_alu_loop_op_5_else_else_if_acc_nl = conv_s2u_32_33(AluIn_data_sva_501[159:128])
      + conv_s2u_32_33({(~ IntShiftLeft_16U_6U_32U_return_31_5_sva_2) , (~ IntShiftLeft_16U_6U_32U_return_30_1_5_sva_2)
      , (~ IntShiftLeft_16U_6U_32U_return_0_5_sva_2)}) + 33'b1;
  assign alu_loop_op_5_else_else_if_acc_nl = nl_alu_loop_op_5_else_else_if_acc_nl[32:0];
  assign alu_loop_op_5_else_else_if_acc_itm_32_1 = readslicef_33_1_32((alu_loop_op_5_else_else_if_acc_nl));
  assign nl_alu_loop_op_4_else_if_acc_1_nl = conv_s2u_32_33({IntShiftLeft_16U_6U_32U_return_31_4_sva_2
      , IntShiftLeft_16U_6U_32U_return_30_1_4_sva_2 , IntShiftLeft_16U_6U_32U_return_0_4_sva_2})
      - conv_s2u_32_33(AluIn_data_sva_501[127:96]);
  assign alu_loop_op_4_else_if_acc_1_nl = nl_alu_loop_op_4_else_if_acc_1_nl[32:0];
  assign alu_loop_op_4_else_if_acc_1_itm_32_1 = readslicef_33_1_32((alu_loop_op_4_else_if_acc_1_nl));
  assign nl_alu_loop_op_4_else_else_if_acc_1_nl = conv_s2u_32_33(AluIn_data_sva_501[127:96])
      + conv_s2u_32_33({(~ IntShiftLeft_16U_6U_32U_return_31_4_sva_2) , (~ IntShiftLeft_16U_6U_32U_return_30_1_4_sva_2)
      , (~ IntShiftLeft_16U_6U_32U_return_0_4_sva_2)}) + 33'b1;
  assign alu_loop_op_4_else_else_if_acc_1_nl = nl_alu_loop_op_4_else_else_if_acc_1_nl[32:0];
  assign alu_loop_op_4_else_else_if_acc_1_itm_32_1 = readslicef_33_1_32((alu_loop_op_4_else_else_if_acc_1_nl));
  assign nl_alu_loop_op_3_else_if_acc_nl = conv_s2u_32_33({IntShiftLeft_16U_6U_32U_return_31_3_sva_2
      , IntShiftLeft_16U_6U_32U_return_30_1_3_sva_2 , IntShiftLeft_16U_6U_32U_return_0_3_sva_2})
      - conv_s2u_32_33(AluIn_data_sva_501[95:64]);
  assign alu_loop_op_3_else_if_acc_nl = nl_alu_loop_op_3_else_if_acc_nl[32:0];
  assign alu_loop_op_3_else_if_acc_itm_32_1 = readslicef_33_1_32((alu_loop_op_3_else_if_acc_nl));
  assign nl_alu_loop_op_3_else_else_if_acc_nl = conv_s2u_32_33(AluIn_data_sva_501[95:64])
      + conv_s2u_32_33({(~ IntShiftLeft_16U_6U_32U_return_31_3_sva_2) , (~ IntShiftLeft_16U_6U_32U_return_30_1_3_sva_2)
      , (~ IntShiftLeft_16U_6U_32U_return_0_3_sva_2)}) + 33'b1;
  assign alu_loop_op_3_else_else_if_acc_nl = nl_alu_loop_op_3_else_else_if_acc_nl[32:0];
  assign alu_loop_op_3_else_else_if_acc_itm_32_1 = readslicef_33_1_32((alu_loop_op_3_else_else_if_acc_nl));
  assign nl_alu_loop_op_2_else_if_acc_1_nl = conv_s2u_32_33({IntShiftLeft_16U_6U_32U_return_31_2_sva_2
      , IntShiftLeft_16U_6U_32U_return_30_1_2_sva_2 , IntShiftLeft_16U_6U_32U_return_0_2_sva_2})
      - conv_s2u_32_33(AluIn_data_sva_501[63:32]);
  assign alu_loop_op_2_else_if_acc_1_nl = nl_alu_loop_op_2_else_if_acc_1_nl[32:0];
  assign alu_loop_op_2_else_if_acc_1_itm_32_1 = readslicef_33_1_32((alu_loop_op_2_else_if_acc_1_nl));
  assign nl_alu_loop_op_2_else_else_if_acc_1_nl = conv_s2u_32_33(AluIn_data_sva_501[63:32])
      + conv_s2u_32_33({(~ IntShiftLeft_16U_6U_32U_return_31_2_sva_2) , (~ IntShiftLeft_16U_6U_32U_return_30_1_2_sva_2)
      , (~ IntShiftLeft_16U_6U_32U_return_0_2_sva_2)}) + 33'b1;
  assign alu_loop_op_2_else_else_if_acc_1_nl = nl_alu_loop_op_2_else_else_if_acc_1_nl[32:0];
  assign alu_loop_op_2_else_else_if_acc_1_itm_32_1 = readslicef_33_1_32((alu_loop_op_2_else_else_if_acc_1_nl));
  assign nl_alu_loop_op_1_else_if_acc_nl = conv_s2u_32_33({IntShiftLeft_16U_6U_32U_return_31_1_sva_2
      , IntShiftLeft_16U_6U_32U_return_30_1_1_sva_2 , IntShiftLeft_16U_6U_32U_return_0_1_sva_2})
      - conv_s2u_32_33(AluIn_data_sva_501[31:0]);
  assign alu_loop_op_1_else_if_acc_nl = nl_alu_loop_op_1_else_if_acc_nl[32:0];
  assign alu_loop_op_1_else_if_acc_itm_32_1 = readslicef_33_1_32((alu_loop_op_1_else_if_acc_nl));
  assign nl_alu_loop_op_1_else_else_if_acc_nl = conv_s2u_32_33(AluIn_data_sva_501[31:0])
      + conv_s2u_32_33({(~ IntShiftLeft_16U_6U_32U_return_31_1_sva_2) , (~ IntShiftLeft_16U_6U_32U_return_30_1_1_sva_2)
      , (~ IntShiftLeft_16U_6U_32U_return_0_1_sva_2)}) + 33'b1;
  assign alu_loop_op_1_else_else_if_acc_nl = nl_alu_loop_op_1_else_else_if_acc_nl[32:0];
  assign alu_loop_op_1_else_else_if_acc_itm_32_1 = readslicef_33_1_32((alu_loop_op_1_else_else_if_acc_nl));
  assign nor_2056_nl = ~((cfg_alu_algo_1_sva_st_92!=2'b10) | io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign nor_2057_nl = ~((reg_cfg_alu_algo_1_sva_st_93_cse!=2'b10) | (~ reg_chn_alu_out_rsci_ld_core_psct_cse)
      | chn_alu_out_rsci_bawt | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign not_tmp_4 = MUX_s_1_2_2((nor_2057_nl), (nor_2056_nl), and_89_tmp);
  assign or_22_cse = (cfg_precision!=2'b10);
  assign or_tmp_20 = ((cfg_alu_algo_1_sva_st_92==2'b11)) | io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign or_32_nl = ((reg_cfg_alu_algo_1_sva_st_93_cse==2'b11)) | (~ reg_chn_alu_out_rsci_ld_core_psct_cse)
      | chn_alu_out_rsci_bawt | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign mux_16_itm = MUX_s_1_2_2((or_32_nl), or_tmp_20, and_89_tmp);
  assign or_tmp_24 = FpCmp_8U_23U_true_if_acc_18_itm_8_1 | (cfg_precision!=2'b10)
      | io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign or_tmp_39 = alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_st_2 | io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign or_tmp_55 = alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_st_2 | io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign or_tmp_76 = alu_loop_op_4_FpCmp_8U_23U_false_slc_8_1_svs_st_2 | io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign or_tmp_97 = alu_loop_op_5_FpCmp_8U_23U_false_slc_8_svs_st_2 | io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign or_tmp_263 = (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt
      | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign mux_127_itm = MUX_s_1_2_2(or_tmp_263, io_read_cfg_alu_bypass_rsc_svs_st_1,
      and_89_tmp);
  assign nor_2061_cse = ~((~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt);
  assign or_tmp_327 = nor_2061_cse | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign or_tmp_329 = (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt
      | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign or_341_nl = io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign mux_tmp_149 = MUX_s_1_2_2(or_1935_cse, (or_341_nl), or_cse_2);
  assign or_334_cse = (cfg_alu_algo_1_sva_st_204!=2'b10);
  assign nor_1962_nl = ~(io_read_cfg_alu_bypass_rsc_svs_st_5 | (reg_cfg_alu_algo_1_sva_st_93_cse[0])
      | (~((reg_cfg_alu_algo_1_sva_st_93_cse[1]) & main_stage_v_2)));
  assign not_tmp_79 = MUX_s_1_2_2(nor_1743_cse, (nor_1962_nl), or_cse_2);
  assign mux_tmp_156 = MUX_s_1_2_2(main_stage_v_3, main_stage_v_2, or_cse_2);
  assign or_350_cse = (reg_cfg_alu_algo_1_sva_st_93_cse!=2'b10);
  assign or_tmp_670 = nor_2061_cse | io_read_cfg_alu_bypass_rsc_svs_st_6 | (~ main_stage_v_3);
  assign mux_tmp_339 = MUX_s_1_2_2(or_899_cse, or_1935_cse, or_cse_2);
  assign or_878_cse = (cfg_alu_algo_1_sva_st_205!=2'b10) | (~ reg_chn_alu_out_rsci_ld_core_psct_cse)
      | chn_alu_out_rsci_bawt | io_read_cfg_alu_bypass_rsc_svs_7 | (~ main_stage_v_4);
  assign or_879_cse = (cfg_alu_algo_1_sva_st_205!=2'b10);
  assign mux_392_nl = MUX_s_1_2_2(mux_tmp_339, or_tmp_670, or_879_cse);
  assign mux_393_itm = MUX_s_1_2_2((mux_392_nl), or_878_cse, or_334_cse);
  assign or_902_nl = (cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48)
      | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6 | (~ or_cse_2);
  assign or_904_nl = (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6 | (~
      or_cse_2);
  assign mux_tmp_392 = MUX_s_1_2_2((or_904_nl), (or_902_nl), FpAlu_8U_23U_equal_tmp_146);
  assign and_224_nl = ((cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48)
      | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6) & or_cse_2;
  assign and_225_nl = or_1935_cse & or_cse_2;
  assign mux_tmp_393 = MUX_s_1_2_2((and_225_nl), (and_224_nl), FpAlu_8U_23U_equal_tmp_146);
  assign mux_414_nl = MUX_s_1_2_2(or_tmp_670, mux_tmp_339, nor_327_cse);
  assign mux_415_itm = MUX_s_1_2_2((mux_414_nl), or_878_cse, or_334_cse);
  assign or_1128_cse = (cfg_alu_algo_1_sva_st_204!=2'b10) | or_tmp_670;
  assign mux_477_cse = MUX_s_1_2_2(mux_tmp_339, or_1827_cse, or_334_cse);
  assign mux_478_itm = MUX_s_1_2_2(mux_477_cse, or_1128_cse, or_879_cse);
  assign mux_604_itm = MUX_s_1_2_2(or_1128_cse, mux_477_cse, nor_327_cse);
  assign or_tmp_1848 = cfg_alu_bypass_rsci_d | ((cfg_alu_algo_rsci_d==2'b11)) | (cfg_precision!=2'b10);
  assign mux_782_itm = MUX_s_1_2_2(io_read_cfg_alu_bypass_rsc_svs_st_1, cfg_alu_bypass_rsci_d,
      and_91_tmp);
  assign or_tmp_1857 = nor_2061_cse | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_precision!=2'b10);
  assign or_1868_nl = FpAdd_8U_23U_mux_2_tmp_49 | (cfg_alu_algo_1_sva_st_204[0])
      | or_tmp_1857;
  assign nor_1329_nl = ~((~ FpAdd_8U_23U_mux_2_tmp_49) | (cfg_alu_algo_1_sva_st_204[0])
      | or_tmp_1857);
  assign mux_784_nl = MUX_s_1_2_2((nor_1329_nl), (or_1868_nl), alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm);
  assign mux_tmp_778 = MUX_s_1_2_2(alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm,
      (mux_784_nl), cfg_alu_algo_1_sva_st_204[1]);
  assign or_1872_nl = FpAdd_8U_23U_mux_18_tmp_49 | (cfg_alu_algo_1_sva_st_204!=2'b10)
      | or_tmp_1857;
  assign nor_1327_nl = ~((~ FpAdd_8U_23U_mux_18_tmp_49) | (cfg_alu_algo_1_sva_st_204!=2'b10)
      | or_tmp_1857);
  assign mux_tmp_779 = MUX_s_1_2_2((nor_1327_nl), (or_1872_nl), alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm);
  assign or_tmp_1865 = (cfg_alu_algo_1_sva_st_204[0]) | or_tmp_1857;
  assign or_1876_nl = alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm
      | (~ or_tmp_1865);
  assign and_284_nl = alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm
      & or_tmp_1865;
  assign mux_787_nl = MUX_s_1_2_2((and_284_nl), (or_1876_nl), FpAdd_8U_23U_mux_34_tmp_49);
  assign mux_tmp_781 = MUX_s_1_2_2(alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm,
      (mux_787_nl), cfg_alu_algo_1_sva_st_204[1]);
  assign or_tmp_1868 = (cfg_alu_algo_1_sva_st_204!=2'b10) | or_tmp_1857;
  assign or_1879_nl = alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm
      | (~ or_tmp_1868);
  assign and_285_nl = alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm
      & or_tmp_1868;
  assign mux_tmp_782 = MUX_s_1_2_2((and_285_nl), (or_1879_nl), FpAdd_8U_23U_mux_50_tmp_49);
  assign or_1882_nl = alu_loop_op_5_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm
      | (~ or_tmp_1868);
  assign and_286_nl = alu_loop_op_5_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm
      & or_tmp_1868;
  assign mux_tmp_783 = MUX_s_1_2_2((and_286_nl), (or_1882_nl), FpAdd_8U_23U_mux_66_tmp_49);
  assign or_1884_nl = FpAdd_8U_23U_mux_82_tmp_49 | or_tmp_1857;
  assign and_3691_nl = FpAdd_8U_23U_mux_82_tmp_49 & (~ or_tmp_1857);
  assign mux_791_nl = MUX_s_1_2_2((and_3691_nl), (or_1884_nl), alu_loop_op_6_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm);
  assign mux_tmp_785 = MUX_s_1_2_2((mux_791_nl), alu_loop_op_6_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm,
      or_334_cse);
  assign or_1886_nl = FpAdd_8U_23U_mux_98_tmp_49 | (cfg_alu_algo_1_sva_st_204!=2'b10)
      | or_tmp_1857;
  assign nor_1326_nl = ~((~ FpAdd_8U_23U_mux_98_tmp_49) | (cfg_alu_algo_1_sva_st_204!=2'b10)
      | or_tmp_1857);
  assign mux_tmp_786 = MUX_s_1_2_2((nor_1326_nl), (or_1886_nl), alu_loop_op_7_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm);
  assign or_1890_nl = (~ (cfg_alu_algo_1_sva_st_204[1])) | FpAdd_8U_23U_mux_114_tmp_49
      | (cfg_alu_algo_1_sva_st_204[0]) | or_tmp_1857;
  assign nor_1325_nl = ~((~ (cfg_alu_algo_1_sva_st_204[1])) | (~ FpAdd_8U_23U_mux_114_tmp_49)
      | (cfg_alu_algo_1_sva_st_204[0]) | or_tmp_1857);
  assign mux_tmp_787 = MUX_s_1_2_2((nor_1325_nl), (or_1890_nl), alu_loop_op_8_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm);
  assign or_1894_nl = FpAdd_8U_23U_mux_130_tmp_49 | (cfg_alu_algo_1_sva_st_204!=2'b10)
      | or_tmp_1857;
  assign nor_1324_nl = ~((~ FpAdd_8U_23U_mux_130_tmp_49) | (cfg_alu_algo_1_sva_st_204!=2'b10)
      | or_tmp_1857);
  assign mux_tmp_788 = MUX_s_1_2_2((nor_1324_nl), (or_1894_nl), alu_loop_op_9_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm);
  assign or_1899_nl = alu_loop_op_10_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm
      | (~ or_tmp_1868);
  assign and_287_nl = alu_loop_op_10_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm
      & or_tmp_1868;
  assign mux_tmp_789 = MUX_s_1_2_2((and_287_nl), (or_1899_nl), FpAdd_8U_23U_mux_146_tmp_49);
  assign or_1901_nl = FpAdd_8U_23U_mux_162_tmp_49 | (cfg_alu_algo_1_sva_st_204!=2'b10)
      | or_tmp_1857;
  assign nor_1323_nl = ~((~ FpAdd_8U_23U_mux_162_tmp_49) | (cfg_alu_algo_1_sva_st_204!=2'b10)
      | or_tmp_1857);
  assign mux_tmp_790 = MUX_s_1_2_2((nor_1323_nl), (or_1901_nl), alu_loop_op_11_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm);
  assign or_1905_nl = FpAdd_8U_23U_mux_178_tmp_49 | (cfg_alu_algo_1_sva_st_204!=2'b10)
      | or_tmp_1857;
  assign nor_1322_nl = ~((~ FpAdd_8U_23U_mux_178_tmp_49) | (cfg_alu_algo_1_sva_st_204!=2'b10)
      | or_tmp_1857);
  assign mux_tmp_791 = MUX_s_1_2_2((nor_1322_nl), (or_1905_nl), alu_loop_op_12_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm);
  assign or_1909_nl = FpAdd_8U_23U_mux_194_tmp_49 | (cfg_alu_algo_1_sva_st_204!=2'b10)
      | or_tmp_1857;
  assign nor_1321_nl = ~((~ FpAdd_8U_23U_mux_194_tmp_49) | (cfg_alu_algo_1_sva_st_204!=2'b10)
      | or_tmp_1857);
  assign mux_tmp_792 = MUX_s_1_2_2((nor_1321_nl), (or_1909_nl), alu_loop_op_13_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm);
  assign or_1913_nl = (cfg_alu_algo_1_sva_st_204!=2'b10) | FpAdd_8U_23U_mux_210_tmp_49
      | or_tmp_1857;
  assign nor_1320_nl = ~((cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAdd_8U_23U_mux_210_tmp_49)
      | or_tmp_1857);
  assign mux_tmp_793 = MUX_s_1_2_2((nor_1320_nl), (or_1913_nl), alu_loop_op_14_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm);
  assign or_1915_nl = FpAdd_8U_23U_mux_226_tmp_49 | or_tmp_1857;
  assign and_3690_nl = FpAdd_8U_23U_mux_226_tmp_49 & (~ or_tmp_1857);
  assign mux_801_nl = MUX_s_1_2_2((and_3690_nl), (or_1915_nl), alu_loop_op_15_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm);
  assign mux_tmp_795 = MUX_s_1_2_2((mux_801_nl), alu_loop_op_15_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm,
      or_334_cse);
  assign or_1917_nl = FpAdd_8U_23U_mux_242_tmp_49 | (cfg_alu_algo_1_sva_st_204!=2'b10)
      | or_tmp_1857;
  assign nor_1319_nl = ~((~ FpAdd_8U_23U_mux_242_tmp_49) | (cfg_alu_algo_1_sva_st_204!=2'b10)
      | or_tmp_1857);
  assign mux_tmp_796 = MUX_s_1_2_2((nor_1319_nl), (or_1917_nl), alu_loop_op_16_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm);
  assign or_tmp_1915 = (reg_cfg_alu_algo_1_sva_st_93_cse[0]) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign mux_829_nl = MUX_s_1_2_2(or_1935_cse, (~ main_stage_v_2), or_cse_2);
  assign mux_tmp_823 = MUX_s_1_2_2((mux_829_nl), or_tmp_329, io_read_cfg_alu_bypass_rsc_svs_st_5);
  assign or_2494_nl = FpAlu_8U_23U_equal_tmp_2 | (~ (reg_cfg_alu_algo_1_sva_st_93_cse[0]));
  assign and_3623_nl = FpAlu_8U_23U_equal_tmp_2 & (reg_cfg_alu_algo_1_sva_st_93_cse[0]);
  assign mux_tmp_1077 = MUX_s_1_2_2((and_3623_nl), (or_2494_nl), FpAlu_8U_23U_equal_tmp);
  assign or_tmp_2842 = nor_2061_cse | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2)
      | (cfg_precision!=2'b10);
  assign or_2855_nl = (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt
      | (~ main_stage_v_2);
  assign mux_1424_nl = MUX_s_1_2_2((or_2855_nl), or_tmp_263, io_read_cfg_alu_bypass_rsc_svs_st_5);
  assign mux_1425_itm = MUX_s_1_2_2((mux_1424_nl), io_read_cfg_alu_bypass_rsc_svs_st_1,
      and_89_tmp);
  assign and_dcpl_7 = (~ chn_alu_out_rsci_bawt) & reg_chn_alu_out_rsci_ld_core_psct_cse;
  assign and_dcpl_8 = or_cse_2 & main_stage_v_4;
  assign and_dcpl_10 = (~ main_stage_v_4) & chn_alu_out_rsci_bawt & reg_chn_alu_out_rsci_ld_core_psct_cse;
  assign and_dcpl_11 = and_91_tmp & (~ cfg_alu_bypass_rsci_d);
  assign or_dcpl_3 = (~ and_91_tmp) | cfg_alu_bypass_rsci_d;
  assign and_dcpl_14 = (~ io_read_cfg_alu_bypass_rsc_svs_st_1) & and_89_tmp & cfg_alu_src_1_sva_st_1;
  assign and_dcpl_21 = (cfg_precision==2'b10);
  assign and_dcpl_22 = and_dcpl_21 & and_89_tmp;
  assign and_dcpl_23 = or_22_cse & and_89_tmp;
  assign and_dcpl_28 = (~ io_read_cfg_alu_bypass_rsc_svs_st_1) & (cfg_precision[1]);
  assign and_dcpl_29 = and_dcpl_28 & (~ (cfg_precision[0])) & and_89_tmp;
  assign or_dcpl_13 = io_read_cfg_alu_bypass_rsc_svs_st_1 | (~ (cfg_precision[1]));
  assign or_dcpl_14 = or_dcpl_13 | (cfg_precision[0]);
  assign and_dcpl_30 = or_dcpl_14 & and_89_tmp;
  assign and_dcpl_34 = or_22_cse & and_89_tmp & (cfg_alu_algo_1_sva_st_92[0]);
  assign and_dcpl_36 = and_dcpl_23 & (cfg_alu_algo_1_sva_st_92==2'b00);
  assign and_dcpl_122 = (~ (cfg_alu_algo_1_sva_st_92[1])) & and_89_tmp;
  assign and_dcpl_126 = or_22_cse & (~ (cfg_alu_algo_1_sva_st_92[0]));
  assign and_dcpl_127 = and_dcpl_126 & and_dcpl_122;
  assign and_dcpl_241 = or_22_cse & or_cse_2;
  assign and_dcpl_256 = or_cse_2 & (~ IsNaN_8U_23U_1_land_15_lpi_1_dfm_8);
  assign and_dcpl_263 = or_cse_2 & (~ IsNaN_8U_23U_2_land_14_lpi_1_dfm_8);
  assign and_dcpl_294 = or_cse_2 & (~ IsNaN_8U_23U_2_land_10_lpi_1_dfm_8);
  assign and_dcpl_309 = or_cse_2 & (~ IsNaN_8U_23U_1_land_8_lpi_1_dfm_8);
  assign and_dcpl_316 = or_cse_2 & (~ IsNaN_8U_23U_1_land_7_lpi_1_dfm_8);
  assign and_dcpl_347 = or_cse_2 & (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_8);
  assign and_dcpl_354 = or_cse_2 & (~ IsNaN_8U_23U_2_land_2_lpi_1_dfm_8);
  assign and_dcpl_361 = or_cse_2 & (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_8);
  assign or_dcpl_112 = (cfg_alu_algo_1_sva_6!=2'b01);
  assign xor_cse = or_dcpl_112 ^ (reg_cfg_alu_algo_1_sva_st_110_cse[0]);
  assign and_dcpl_369 = xor_cse & or_22_cse & or_cse_2 & (~ io_read_cfg_alu_bypass_rsc_svs_st_6)
      & (~ (reg_cfg_alu_algo_1_sva_st_110_cse[1]));
  assign or_dcpl_113 = (reg_cfg_alu_algo_1_sva_st_110_cse!=2'b01);
  assign and_dcpl_372 = (((and_dcpl_21 | or_dcpl_113) & (cfg_alu_algo_1_sva_6==2'b01))
      | io_read_cfg_alu_bypass_rsc_svs_st_6) & or_cse_2;
  assign or_dcpl_116 = (reg_cfg_alu_algo_1_sva_st_110_cse!=2'b00);
  assign and_dcpl_375 = (and_dcpl_21 | or_dcpl_116) & or_dcpl_112 & or_cse_2 & (~
      io_read_cfg_alu_bypass_rsc_svs_st_6);
  assign and_dcpl_379 = xor_cse & or_22_cse & or_cse_2 & (~(io_read_cfg_alu_bypass_rsc_svs_st_6
      | (reg_cfg_alu_algo_1_sva_st_110_cse[1])));
  assign and_dcpl_394 = and_dcpl_21 & and_91_tmp;
  assign and_dcpl_395 = or_22_cse & and_91_tmp;
  assign and_dcpl_397 = (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10);
  assign and_dcpl_398 = and_dcpl_21 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5);
  assign and_dcpl_401 = FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w4 & or_cse_2;
  assign and_dcpl_402 = and_dcpl_401 & and_dcpl_398 & and_dcpl_397;
  assign and_dcpl_404 = (~ alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_2) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10);
  assign and_dcpl_406 = (~((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_itm_23_1) &
      alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2)) & or_cse_2;
  assign and_dcpl_407 = and_dcpl_406 & and_dcpl_398 & and_dcpl_404;
  assign or_dcpl_131 = or_22_cse | io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign and_dcpl_408 = (or_dcpl_131 | or_350_cse) & or_cse_2;
  assign or_dcpl_137 = or_22_cse | or_1935_cse | and_dcpl_7 | or_334_cse;
  assign and_3551_nl = (~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_itm_23_1) & alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_st_2;
  assign mux_tmp_1500 = MUX_s_1_2_2(alu_loop_op_2_FpAdd_8U_23U_is_a_greater_slc_8_1_svs_st_2,
      (~ alu_loop_op_2_FpAdd_8U_23U_is_a_greater_slc_8_1_svs_st_2), and_3551_nl);
  assign and_dcpl_416 = ((mux_tmp_1500 & alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2)
      | alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_2) & or_cse_2;
  assign and_dcpl_417 = and_dcpl_416 & and_dcpl_398 & and_dcpl_397;
  assign and_dcpl_419 = (~ alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_2) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10);
  assign and_dcpl_421 = (~(mux_tmp_1500 & alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2))
      & or_cse_2;
  assign and_dcpl_422 = and_dcpl_421 & and_dcpl_398 & and_dcpl_419;
  assign and_dcpl_431 = FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w4 & or_cse_2;
  assign and_dcpl_432 = and_dcpl_431 & and_dcpl_398 & and_dcpl_397;
  assign and_dcpl_434 = (~ alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_2) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10);
  assign and_dcpl_436 = (~((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_itm_23_1)
      & alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2)) & or_cse_2;
  assign and_dcpl_437 = and_dcpl_436 & and_dcpl_398 & and_dcpl_434;
  assign and_dcpl_446 = FpAdd_8U_23U_is_a_greater_lor_4_lpi_1_dfm_1_mx0w4 & or_cse_2;
  assign and_dcpl_447 = and_dcpl_446 & and_dcpl_398 & and_dcpl_397;
  assign and_dcpl_449 = (~ alu_loop_op_4_FpCmp_8U_23U_false_slc_8_1_svs_2) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10);
  assign and_dcpl_451 = (~((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_itm_23_1)
      & alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2)) & or_cse_2;
  assign and_dcpl_452 = and_dcpl_451 & and_dcpl_398 & and_dcpl_449;
  assign and_dcpl_473 = FpAdd_8U_23U_is_a_greater_lor_8_lpi_1_dfm_1_mx0w4 & or_cse_2;
  assign and_dcpl_474 = and_dcpl_473 & and_dcpl_398 & and_dcpl_397;
  assign and_dcpl_476 = (~ alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_2) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10);
  assign and_dcpl_478 = (~((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_7_itm_23_1)
      & alu_loop_op_8_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2)) & or_cse_2;
  assign and_dcpl_479 = and_dcpl_478 & and_dcpl_398 & and_dcpl_476;
  assign and_dcpl_504 = FpAdd_8U_23U_is_a_greater_lor_13_lpi_1_dfm_1_mx0w4 & or_cse_2;
  assign and_dcpl_505 = and_dcpl_504 & and_dcpl_398 & and_dcpl_397;
  assign and_dcpl_507 = (~ alu_loop_op_13_FpCmp_8U_23U_false_slc_8_svs_2) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10);
  assign and_dcpl_509 = (~((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_12_itm_23_1)
      & alu_loop_op_13_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2)) & or_cse_2;
  assign and_dcpl_510 = and_dcpl_509 & and_dcpl_398 & and_dcpl_507;
  assign and_dcpl_519 = FpAdd_8U_23U_is_a_greater_lor_14_lpi_1_dfm_1_mx0w4 & or_cse_2;
  assign and_dcpl_520 = and_dcpl_519 & and_dcpl_398 & and_dcpl_397;
  assign and_dcpl_522 = (~ alu_loop_op_14_FpCmp_8U_23U_false_slc_8_1_svs_2) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10);
  assign and_dcpl_524 = (~((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_13_itm_23_1)
      & alu_loop_op_14_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2)) & or_cse_2;
  assign and_dcpl_525 = and_dcpl_524 & and_dcpl_398 & and_dcpl_522;
  assign and_dcpl_534 = FpAdd_8U_23U_is_a_greater_lor_15_lpi_1_dfm_1_mx0w4 & or_cse_2;
  assign and_dcpl_535 = and_dcpl_534 & and_dcpl_398 & and_dcpl_397;
  assign and_dcpl_537 = (reg_cfg_alu_algo_1_sva_st_93_cse[1]) & (~ alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_2)
      & (~ (reg_cfg_alu_algo_1_sva_st_93_cse[0]));
  assign and_dcpl_539 = (~((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_14_itm_23_1)
      & alu_loop_op_15_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2)) & or_cse_2;
  assign and_dcpl_540 = and_dcpl_539 & and_dcpl_398 & and_dcpl_537;
  assign and_dcpl_549 = FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w4 & or_cse_2;
  assign and_dcpl_550 = and_dcpl_549 & and_dcpl_398 & and_dcpl_397;
  assign and_dcpl_552 = (~ alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_2) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10);
  assign and_dcpl_554 = (~((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_15_itm_23_1)
      & alu_loop_op_16_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2)) & or_cse_2;
  assign and_dcpl_555 = and_dcpl_554 & and_dcpl_398 & and_dcpl_552;
  assign or_dcpl_219 = and_dcpl_21 | or_1935_cse;
  assign and_dcpl_564 = FpAdd_8U_23U_is_a_greater_lor_5_lpi_1_dfm_1_mx0w4 & or_cse_2;
  assign and_dcpl_565 = and_dcpl_564 & and_dcpl_398 & and_dcpl_397;
  assign and_dcpl_567 = (~ alu_loop_op_5_FpCmp_8U_23U_false_slc_8_svs_2) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10);
  assign and_dcpl_569 = (~((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_itm_23_1)
      & alu_loop_op_5_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2)) & or_cse_2;
  assign and_dcpl_570 = and_dcpl_569 & and_dcpl_398 & and_dcpl_567;
  assign and_dcpl_575 = FpAdd_8U_23U_is_a_greater_lor_6_lpi_1_dfm_1_mx0w4 & or_cse_2;
  assign and_dcpl_576 = and_dcpl_575 & and_dcpl_398 & and_dcpl_397;
  assign and_dcpl_578 = (~ alu_loop_op_6_FpCmp_8U_23U_false_slc_8_1_svs_2) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10);
  assign and_dcpl_580 = (~((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_5_itm_23_1)
      & alu_loop_op_6_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2)) & or_cse_2;
  assign and_dcpl_581 = and_dcpl_580 & and_dcpl_398 & and_dcpl_578;
  assign and_dcpl_586 = FpAdd_8U_23U_is_a_greater_lor_7_lpi_1_dfm_1_mx0w4 & or_cse_2;
  assign and_dcpl_587 = and_dcpl_586 & and_dcpl_398 & and_dcpl_397;
  assign and_dcpl_589 = (~ alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_2) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10);
  assign and_dcpl_591 = (~((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_itm_23_1)
      & alu_loop_op_7_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2)) & or_cse_2;
  assign and_dcpl_592 = and_dcpl_591 & and_dcpl_398 & and_dcpl_589;
  assign and_dcpl_597 = FpAdd_8U_23U_is_a_greater_lor_9_lpi_1_dfm_1_mx0w4 & or_cse_2;
  assign and_dcpl_598 = and_dcpl_597 & and_dcpl_398 & and_dcpl_397;
  assign and_dcpl_600 = (~ alu_loop_op_9_FpCmp_8U_23U_false_slc_8_svs_2) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10);
  assign and_dcpl_602 = (~((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_itm_23_1)
      & alu_loop_op_9_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2)) & or_cse_2;
  assign and_dcpl_603 = and_dcpl_602 & and_dcpl_398 & and_dcpl_600;
  assign and_dcpl_608 = FpAdd_8U_23U_is_a_greater_lor_10_lpi_1_dfm_1_mx0w4 & or_cse_2;
  assign and_dcpl_609 = and_dcpl_608 & and_dcpl_398 & and_dcpl_397;
  assign and_dcpl_611 = (~ alu_loop_op_10_FpCmp_8U_23U_false_slc_8_1_svs_2) & (reg_cfg_alu_algo_1_sva_st_93_cse==2'b10);
  assign and_dcpl_613 = (~((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_9_itm_23_1)
      & alu_loop_op_10_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2)) & or_cse_2;
  assign and_dcpl_614 = and_dcpl_613 & and_dcpl_398 & and_dcpl_611;
  assign and_dcpl_619 = FpAdd_8U_23U_is_a_greater_lor_11_lpi_1_dfm_1_mx0w4 & or_cse_2;
  assign and_dcpl_620 = and_dcpl_619 & and_dcpl_398 & and_dcpl_397;
  assign and_dcpl_622 = (reg_cfg_alu_algo_1_sva_st_93_cse[1]) & (~ alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_2)
      & (~ (reg_cfg_alu_algo_1_sva_st_93_cse[0]));
  assign and_dcpl_624 = (~((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_itm_23_1)
      & alu_loop_op_11_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2)) & or_cse_2;
  assign and_dcpl_625 = and_dcpl_624 & and_dcpl_398 & and_dcpl_622;
  assign and_dcpl_630 = FpAdd_8U_23U_is_a_greater_lor_12_lpi_1_dfm_1_mx0w4 & or_cse_2;
  assign and_dcpl_631 = and_dcpl_630 & and_dcpl_398 & and_dcpl_397;
  assign and_dcpl_633 = (reg_cfg_alu_algo_1_sva_st_93_cse[1]) & (~ alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_2)
      & (~ (reg_cfg_alu_algo_1_sva_st_93_cse[0]));
  assign and_dcpl_635 = (~((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_11_itm_23_1)
      & alu_loop_op_12_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2)) & or_cse_2;
  assign and_dcpl_636 = and_dcpl_635 & and_dcpl_398 & and_dcpl_633;
  assign and_dcpl_638 = and_dcpl_28 & (~ (cfg_precision[0]));
  assign or_dcpl_295 = (cfg_alu_algo_1_sva_st_92!=2'b10);
  assign and_dcpl_676 = ~((reg_cfg_alu_algo_1_sva_st_93_cse!=2'b00));
  assign and_dcpl_695 = ~(io_read_cfg_alu_bypass_rsc_svs_st_5 | (reg_cfg_alu_algo_1_sva_st_157_cse[1]));
  assign or_3303_cse = (cfg_alu_algo_1_sva_5!=2'b01);
  assign nor_913_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | (~ alu_loop_op_3_else_if_acc_itm_32_1));
  assign and_3550_nl = (reg_cfg_alu_algo_1_sva_st_157_cse[0]) & alu_loop_op_3_else_else_if_acc_itm_32_1;
  assign mux_1522_nl = MUX_s_1_2_2((and_3550_nl), (nor_913_nl), or_3303_cse);
  assign and_dcpl_698 = (mux_1522_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_911_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | alu_loop_op_3_else_if_acc_itm_32_1);
  assign nor_912_nl = ~((~ (reg_cfg_alu_algo_1_sva_st_157_cse[0])) | alu_loop_op_3_else_else_if_acc_itm_32_1);
  assign mux_1523_nl = MUX_s_1_2_2((nor_912_nl), (nor_911_nl), or_3303_cse);
  assign and_dcpl_701 = (mux_1523_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign and_dcpl_704 = (((and_dcpl_21 | (reg_cfg_alu_algo_1_sva_st_157_cse!=2'b01))
      & FpAlu_8U_23U_equal_tmp_2_mx0w0) | io_read_cfg_alu_bypass_rsc_svs_st_5) &
      or_cse_2;
  assign and_dcpl_707 = (and_dcpl_21 | (reg_cfg_alu_algo_1_sva_st_157_cse!=2'b00))
      & or_cse_2 & (~((~((cfg_alu_algo_1_sva_5!=2'b01))) | io_read_cfg_alu_bypass_rsc_svs_st_5));
  assign nor_910_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | (~ alu_loop_op_5_else_if_acc_itm_32_1));
  assign and_3549_nl = (reg_cfg_alu_algo_1_sva_st_157_cse[0]) & alu_loop_op_5_else_else_if_acc_itm_32_1;
  assign mux_1524_nl = MUX_s_1_2_2((and_3549_nl), (nor_910_nl), or_3303_cse);
  assign and_dcpl_711 = (mux_1524_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_908_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | alu_loop_op_5_else_if_acc_itm_32_1);
  assign nor_909_nl = ~((~ (reg_cfg_alu_algo_1_sva_st_157_cse[0])) | alu_loop_op_5_else_else_if_acc_itm_32_1);
  assign mux_1525_nl = MUX_s_1_2_2((nor_909_nl), (nor_908_nl), or_3303_cse);
  assign and_dcpl_714 = (mux_1525_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_907_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | (~ alu_loop_op_6_else_if_acc_1_itm_32_1));
  assign and_3548_nl = (reg_cfg_alu_algo_1_sva_st_157_cse[0]) & alu_loop_op_6_else_else_if_acc_1_itm_32_1;
  assign mux_1526_nl = MUX_s_1_2_2((and_3548_nl), (nor_907_nl), or_3303_cse);
  assign and_dcpl_722 = (mux_1526_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_905_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | alu_loop_op_6_else_if_acc_1_itm_32_1);
  assign nor_906_nl = ~((~ (reg_cfg_alu_algo_1_sva_st_157_cse[0])) | alu_loop_op_6_else_else_if_acc_1_itm_32_1);
  assign mux_1527_nl = MUX_s_1_2_2((nor_906_nl), (nor_905_nl), or_3303_cse);
  assign and_dcpl_725 = (mux_1527_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_904_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | (~ alu_loop_op_7_else_if_acc_itm_32_1));
  assign and_3547_nl = (reg_cfg_alu_algo_1_sva_st_157_cse[0]) & alu_loop_op_7_else_else_if_acc_itm_32_1;
  assign mux_1528_nl = MUX_s_1_2_2((and_3547_nl), (nor_904_nl), or_3303_cse);
  assign and_dcpl_733 = (mux_1528_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_902_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | alu_loop_op_7_else_if_acc_itm_32_1);
  assign nor_903_nl = ~((~ (reg_cfg_alu_algo_1_sva_st_157_cse[0])) | alu_loop_op_7_else_else_if_acc_itm_32_1);
  assign mux_1529_nl = MUX_s_1_2_2((nor_903_nl), (nor_902_nl), or_3303_cse);
  assign and_dcpl_736 = (mux_1529_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_901_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | (~ alu_loop_op_8_else_if_acc_1_itm_32_1));
  assign and_3546_nl = (reg_cfg_alu_algo_1_sva_st_157_cse[0]) & alu_loop_op_8_else_else_if_acc_1_itm_32_1;
  assign mux_1530_nl = MUX_s_1_2_2((and_3546_nl), (nor_901_nl), or_3303_cse);
  assign and_dcpl_744 = (mux_1530_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_899_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | alu_loop_op_8_else_if_acc_1_itm_32_1);
  assign nor_900_nl = ~((~ (reg_cfg_alu_algo_1_sva_st_157_cse[0])) | alu_loop_op_8_else_else_if_acc_1_itm_32_1);
  assign mux_1531_nl = MUX_s_1_2_2((nor_900_nl), (nor_899_nl), or_3303_cse);
  assign and_dcpl_747 = (mux_1531_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_898_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | (~ alu_loop_op_9_else_if_acc_itm_32_1));
  assign and_3545_nl = (reg_cfg_alu_algo_1_sva_st_157_cse[0]) & alu_loop_op_9_else_else_if_acc_itm_32_1;
  assign mux_1532_nl = MUX_s_1_2_2((and_3545_nl), (nor_898_nl), or_3303_cse);
  assign and_dcpl_755 = (mux_1532_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_896_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | alu_loop_op_9_else_if_acc_itm_32_1);
  assign nor_897_nl = ~((~ (reg_cfg_alu_algo_1_sva_st_157_cse[0])) | alu_loop_op_9_else_else_if_acc_itm_32_1);
  assign mux_1533_nl = MUX_s_1_2_2((nor_897_nl), (nor_896_nl), or_3303_cse);
  assign and_dcpl_758 = (mux_1533_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_895_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | (~ alu_loop_op_10_else_if_acc_1_itm_32_1));
  assign and_3544_nl = (reg_cfg_alu_algo_1_sva_st_157_cse[0]) & alu_loop_op_10_else_else_if_acc_1_itm_32_1;
  assign mux_1534_nl = MUX_s_1_2_2((and_3544_nl), (nor_895_nl), or_3303_cse);
  assign and_dcpl_766 = (mux_1534_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_893_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | alu_loop_op_10_else_if_acc_1_itm_32_1);
  assign nor_894_nl = ~((~ (reg_cfg_alu_algo_1_sva_st_157_cse[0])) | alu_loop_op_10_else_else_if_acc_1_itm_32_1);
  assign mux_1535_nl = MUX_s_1_2_2((nor_894_nl), (nor_893_nl), or_3303_cse);
  assign and_dcpl_769 = (mux_1535_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_892_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | (~ alu_loop_op_11_else_if_acc_itm_32_1));
  assign and_3543_nl = (reg_cfg_alu_algo_1_sva_st_157_cse[0]) & alu_loop_op_11_else_else_if_acc_itm_32_1;
  assign mux_1536_nl = MUX_s_1_2_2((and_3543_nl), (nor_892_nl), or_3303_cse);
  assign and_dcpl_777 = (mux_1536_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_890_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | alu_loop_op_11_else_if_acc_itm_32_1);
  assign nor_891_nl = ~((~ (reg_cfg_alu_algo_1_sva_st_157_cse[0])) | alu_loop_op_11_else_else_if_acc_itm_32_1);
  assign mux_1537_nl = MUX_s_1_2_2((nor_891_nl), (nor_890_nl), or_3303_cse);
  assign and_dcpl_780 = (mux_1537_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_889_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | (~ alu_loop_op_12_else_if_acc_1_itm_32_1));
  assign and_3542_nl = (reg_cfg_alu_algo_1_sva_st_157_cse[0]) & alu_loop_op_12_else_else_if_acc_1_itm_32_1;
  assign mux_1538_nl = MUX_s_1_2_2((and_3542_nl), (nor_889_nl), or_3303_cse);
  assign and_dcpl_788 = (mux_1538_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_887_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | alu_loop_op_12_else_if_acc_1_itm_32_1);
  assign nor_888_nl = ~((~ (reg_cfg_alu_algo_1_sva_st_157_cse[0])) | alu_loop_op_12_else_else_if_acc_1_itm_32_1);
  assign mux_1539_nl = MUX_s_1_2_2((nor_888_nl), (nor_887_nl), or_3303_cse);
  assign and_dcpl_791 = (mux_1539_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_886_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | (~ alu_loop_op_13_else_if_acc_itm_32_1));
  assign and_3541_nl = (reg_cfg_alu_algo_1_sva_st_157_cse[0]) & alu_loop_op_13_else_else_if_acc_itm_32_1;
  assign mux_1540_nl = MUX_s_1_2_2((and_3541_nl), (nor_886_nl), or_3303_cse);
  assign and_dcpl_799 = (mux_1540_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_884_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | alu_loop_op_13_else_if_acc_itm_32_1);
  assign nor_885_nl = ~((~ (reg_cfg_alu_algo_1_sva_st_157_cse[0])) | alu_loop_op_13_else_else_if_acc_itm_32_1);
  assign mux_1541_nl = MUX_s_1_2_2((nor_885_nl), (nor_884_nl), or_3303_cse);
  assign and_dcpl_802 = (mux_1541_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_883_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | (~ alu_loop_op_14_else_if_acc_1_itm_32_1));
  assign and_3540_nl = (reg_cfg_alu_algo_1_sva_st_157_cse[0]) & alu_loop_op_14_else_else_if_acc_1_itm_32_1;
  assign mux_1542_nl = MUX_s_1_2_2((and_3540_nl), (nor_883_nl), or_3303_cse);
  assign and_dcpl_810 = (mux_1542_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_881_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | alu_loop_op_14_else_if_acc_1_itm_32_1);
  assign nor_882_nl = ~((~ (reg_cfg_alu_algo_1_sva_st_157_cse[0])) | alu_loop_op_14_else_else_if_acc_1_itm_32_1);
  assign mux_1543_nl = MUX_s_1_2_2((nor_882_nl), (nor_881_nl), or_3303_cse);
  assign and_dcpl_813 = (mux_1543_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_880_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | (~ alu_loop_op_15_else_if_acc_itm_32_1));
  assign and_3539_nl = (reg_cfg_alu_algo_1_sva_st_157_cse[0]) & alu_loop_op_15_else_else_if_acc_itm_32_1;
  assign mux_1544_nl = MUX_s_1_2_2((and_3539_nl), (nor_880_nl), or_3303_cse);
  assign and_dcpl_821 = (mux_1544_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign nor_878_nl = ~((reg_cfg_alu_algo_1_sva_st_157_cse[0]) | alu_loop_op_15_else_if_acc_itm_32_1);
  assign nor_879_nl = ~((~ (reg_cfg_alu_algo_1_sva_st_157_cse[0])) | alu_loop_op_15_else_else_if_acc_itm_32_1);
  assign mux_1545_nl = MUX_s_1_2_2((nor_879_nl), (nor_878_nl), or_3303_cse);
  assign and_dcpl_824 = (mux_1545_nl) & or_22_cse & or_cse_2 & and_dcpl_695;
  assign and_dcpl_830 = and_dcpl_695 & or_cse_2;
  assign nor_tmp_847 = alu_loop_op_16_else_else_if_acc_1_itm_32_1 & (reg_cfg_alu_algo_1_sva_st_157_cse[0]);
  assign nor_877_nl = ~((~ alu_loop_op_16_else_if_acc_1_itm_32_1) | (reg_cfg_alu_algo_1_sva_st_157_cse[0]));
  assign mux_1546_nl = MUX_s_1_2_2(nor_tmp_847, (nor_877_nl), or_3303_cse);
  assign and_dcpl_832 = (mux_1546_nl) & or_22_cse & and_dcpl_830;
  assign nor_875_nl = ~(alu_loop_op_16_else_if_acc_1_itm_32_1 | (reg_cfg_alu_algo_1_sva_st_157_cse[0]));
  assign nor_876_nl = ~(alu_loop_op_16_else_else_if_acc_1_itm_32_1 | (~ (reg_cfg_alu_algo_1_sva_st_157_cse[0])));
  assign mux_1547_nl = MUX_s_1_2_2((nor_876_nl), (nor_875_nl), or_3303_cse);
  assign and_dcpl_834 = (mux_1547_nl) & or_22_cse & and_dcpl_830;
  assign and_dcpl_840 = or_dcpl_131 & or_cse_2;
  assign and_dcpl_843 = (~ (reg_cfg_alu_algo_1_sva_st_93_cse[1])) & (cfg_alu_algo_1_sva_5[0]);
  assign and_dcpl_844 = or_cse_2 & (AluIn_data_sva_501[31]);
  assign and_dcpl_846 = or_cse_2 & (~ (AluIn_data_sva_501[31]));
  assign and_dcpl_848 = ~((reg_cfg_alu_algo_1_sva_st_93_cse[1]) | (cfg_alu_algo_1_sva_5[0]));
  assign and_dcpl_856 = or_cse_2 & (AluIn_data_sva_501[63]);
  assign and_dcpl_858 = or_cse_2 & (~ (AluIn_data_sva_501[63]));
  assign and_dcpl_879 = or_cse_2 & (cfg_precision[1]);
  assign and_dcpl_884 = or_cse_2 & (AluIn_data_sva_501[127]);
  assign and_dcpl_886 = or_cse_2 & (~ (AluIn_data_sva_501[127]));
  assign and_dcpl_897 = or_cse_2 & (AluIn_data_sva_501[159]);
  assign and_dcpl_899 = or_cse_2 & (~ (AluIn_data_sva_501[159]));
  assign and_dcpl_924 = or_cse_2 & (AluIn_data_sva_501[223]);
  assign and_dcpl_926 = or_cse_2 & (~ (AluIn_data_sva_501[223]));
  assign and_dcpl_946 = or_cse_2 & (AluIn_data_sva_501[287]);
  assign and_dcpl_948 = or_cse_2 & (~ (AluIn_data_sva_501[287]));
  assign and_dcpl_971 = or_cse_2 & (~ (reg_cfg_alu_algo_1_sva_st_93_cse[1]));
  assign and_dcpl_1036 = or_cse_2 & (AluIn_data_sva_501[511]);
  assign and_dcpl_1038 = or_cse_2 & (~ (AluIn_data_sva_501[511]));
  assign mux_tmp_1541 = MUX_s_1_2_2(alu_loop_op_1_else_if_acc_itm_32_1, alu_loop_op_1_else_else_if_acc_itm_32_1,
      reg_cfg_alu_algo_1_sva_st_157_cse[0]);
  assign and_dcpl_1044 = mux_tmp_1541 & or_22_cse & or_cse_2;
  assign and_dcpl_1046 = (~ mux_tmp_1541) & or_22_cse & or_cse_2;
  assign and_dcpl_1048 = and_dcpl_879 & (~ (cfg_precision[0])) & (reg_cfg_alu_algo_1_sva_st_157_cse[0]);
  assign and_dcpl_1050 = and_dcpl_879 & (~ (cfg_precision[0])) & (~ (reg_cfg_alu_algo_1_sva_st_157_cse[0]));
  assign mux_tmp_1542 = MUX_s_1_2_2(alu_loop_op_2_else_if_acc_1_itm_32_1, alu_loop_op_2_else_else_if_acc_1_itm_32_1,
      reg_cfg_alu_algo_1_sva_st_157_cse[0]);
  assign and_dcpl_1052 = mux_tmp_1542 & or_22_cse & or_cse_2;
  assign and_dcpl_1054 = (~ mux_tmp_1542) & or_22_cse & or_cse_2;
  assign mux_tmp_1543 = MUX_s_1_2_2(alu_loop_op_4_else_if_acc_1_itm_32_1, alu_loop_op_4_else_else_if_acc_1_itm_32_1,
      reg_cfg_alu_algo_1_sva_st_157_cse[0]);
  assign and_dcpl_1060 = mux_tmp_1543 & or_22_cse & or_cse_2;
  assign and_dcpl_1062 = (~ mux_tmp_1543) & or_22_cse & or_cse_2;
  assign and_dcpl_1070 = (else_mux_2_tmp[4:2]==3'b111);
  assign and_dcpl_1073 = and_dcpl_638 & (IsNaN_5U_10U_nor_tmp | (~ cfg_nan_to_zero))
      & (else_mux_2_tmp[0]);
  assign or_dcpl_391 = (~((else_mux_2_tmp[0]) & (else_mux_2_tmp[3]))) | (~((else_mux_2_tmp[4])
      & (else_mux_2_tmp[2]))) | ((~ IsNaN_5U_10U_nor_tmp) & cfg_nan_to_zero) | (~
      (else_mux_2_tmp[1])) | IsNaN_5U_23U_nor_tmp;
  assign or_dcpl_393 = or_dcpl_13 | (cfg_precision[0]) | (~ and_89_tmp);
  assign and_dcpl_1079 = and_dcpl_1073 & and_dcpl_1070 & (else_mux_2_tmp[1]) & (~
      IsNaN_5U_23U_nor_tmp);
  assign and_dcpl_1080 = or_dcpl_391 & and_dcpl_638;
  assign or_dcpl_394 = (~ and_89_tmp) | (cfg_alu_algo_1_sva_st_92[0]);
  assign and_dcpl_1084 = (else_mux_5_tmp[4:2]==3'b111);
  assign and_dcpl_1087 = and_dcpl_638 & (IsNaN_5U_10U_nor_1_tmp | (~ cfg_nan_to_zero))
      & (else_mux_5_tmp[1]);
  assign or_dcpl_411 = (else_mux_5_tmp[4:1]!=4'b1111) | ((~ IsNaN_5U_10U_nor_1_tmp)
      & cfg_nan_to_zero) | (~ (else_mux_5_tmp[0])) | IsNaN_5U_23U_nor_1_tmp;
  assign and_dcpl_1093 = and_dcpl_1087 & and_dcpl_1084 & (else_mux_5_tmp[0]) & (~
      IsNaN_5U_23U_nor_1_tmp);
  assign and_dcpl_1094 = or_dcpl_411 & and_dcpl_638;
  assign or_dcpl_413 = or_dcpl_394 | (~ (cfg_alu_algo_1_sva_st_92[1]));
  assign or_dcpl_414 = or_dcpl_14 | or_dcpl_413;
  assign and_dcpl_1098 = (else_mux_8_tmp[3:1]==3'b111);
  assign and_dcpl_1101 = and_dcpl_638 & (IsNaN_5U_10U_nor_2_tmp | (~ cfg_nan_to_zero))
      & (else_mux_8_tmp[4]);
  assign or_dcpl_429 = (else_mux_8_tmp[4:1]!=4'b1111) | ((~ IsNaN_5U_10U_nor_2_tmp)
      & cfg_nan_to_zero) | (~ (else_mux_8_tmp[0])) | IsNaN_5U_23U_nor_2_tmp;
  assign and_dcpl_1107 = and_dcpl_1101 & and_dcpl_1098 & (else_mux_8_tmp[0]) & (~
      IsNaN_5U_23U_nor_2_tmp);
  assign and_dcpl_1108 = or_dcpl_429 & and_dcpl_638;
  assign and_dcpl_1112 = (else_mux_11_tmp[3:1]==3'b111);
  assign and_dcpl_1115 = and_dcpl_638 & (IsNaN_5U_10U_nor_3_tmp | (~ cfg_nan_to_zero))
      & (else_mux_11_tmp[4]);
  assign or_dcpl_447 = (else_mux_11_tmp[4:1]!=4'b1111) | ((~ IsNaN_5U_10U_nor_3_tmp)
      & cfg_nan_to_zero) | (~ (else_mux_11_tmp[0])) | IsNaN_5U_23U_nor_3_tmp;
  assign and_dcpl_1121 = and_dcpl_1115 & and_dcpl_1112 & (else_mux_11_tmp[0]) & (~
      IsNaN_5U_23U_nor_3_tmp);
  assign and_dcpl_1122 = or_dcpl_447 & and_dcpl_638;
  assign and_dcpl_1123 = (else_mux_14_tmp[1:0]==2'b11);
  assign and_dcpl_1126 = (~ IsNaN_5U_23U_nor_4_tmp) & (else_mux_14_tmp[3:2]==2'b11);
  assign and_dcpl_1129 = and_dcpl_638 & (IsNaN_5U_10U_nor_4_tmp | (~ cfg_nan_to_zero))
      & (else_mux_14_tmp[4]);
  assign or_dcpl_465 = (~ (else_mux_14_tmp[4])) | IsNaN_5U_23U_nor_4_tmp | ((~ IsNaN_5U_10U_nor_4_tmp)
      & cfg_nan_to_zero) | (else_mux_14_tmp[3:0]!=4'b1111);
  assign and_dcpl_1134 = and_dcpl_1129 & and_dcpl_1126 & and_dcpl_1123;
  assign and_dcpl_1135 = or_dcpl_465 & and_dcpl_638;
  assign or_dcpl_477 = IsNaN_5U_10U_nor_5_tmp | (~ cfg_nan_to_zero);
  assign or_dcpl_483 = (else_mux_17_tmp!=5'b11111) | IsNaN_5U_23U_nor_5_tmp | ((~
      IsNaN_5U_10U_nor_5_tmp) & cfg_nan_to_zero);
  assign and_dcpl_1152 = and_dcpl_638 & (else_mux_17_tmp==5'b11111) & (~ IsNaN_5U_23U_nor_5_tmp)
      & or_dcpl_477;
  assign and_dcpl_1153 = or_dcpl_483 & and_dcpl_638;
  assign or_dcpl_495 = (~ cfg_nan_to_zero) | IsNaN_5U_10U_nor_6_tmp;
  assign or_dcpl_501 = (else_mux_20_tmp!=5'b11111) | IsNaN_5U_23U_nor_6_tmp | (cfg_nan_to_zero
      & (~ IsNaN_5U_10U_nor_6_tmp));
  assign and_dcpl_1170 = and_dcpl_638 & (else_mux_20_tmp==5'b11111) & (~ IsNaN_5U_23U_nor_6_tmp)
      & or_dcpl_495;
  assign and_dcpl_1171 = or_dcpl_501 & and_dcpl_638;
  assign or_dcpl_513 = (~ cfg_nan_to_zero) | IsNaN_5U_10U_nor_7_tmp;
  assign or_dcpl_519 = (else_mux_23_tmp!=5'b11111) | IsNaN_5U_23U_nor_7_tmp | (cfg_nan_to_zero
      & (~ IsNaN_5U_10U_nor_7_tmp));
  assign and_dcpl_1188 = and_dcpl_638 & (else_mux_23_tmp[4:3]==2'b11) & (~ IsNaN_5U_23U_nor_7_tmp)
      & (else_mux_23_tmp[2:0]==3'b111) & or_dcpl_513;
  assign and_dcpl_1189 = or_dcpl_519 & and_dcpl_638;
  assign or_dcpl_520 = or_dcpl_295 | (~ and_89_tmp);
  assign or_dcpl_531 = (~ cfg_nan_to_zero) | IsNaN_5U_10U_nor_8_tmp;
  assign or_dcpl_537 = (else_mux_26_tmp!=5'b11111) | IsNaN_5U_23U_nor_8_tmp | (cfg_nan_to_zero
      & (~ IsNaN_5U_10U_nor_8_tmp));
  assign and_dcpl_1206 = and_dcpl_638 & (else_mux_26_tmp[4:3]==2'b11) & (~ IsNaN_5U_23U_nor_8_tmp)
      & (else_mux_26_tmp[2:0]==3'b111) & or_dcpl_531;
  assign and_dcpl_1207 = or_dcpl_537 & and_dcpl_638;
  assign and_dcpl_1211 = (else_mux_29_tmp[2:0]==3'b111);
  assign and_dcpl_1214 = and_dcpl_638 & (IsNaN_5U_10U_nor_9_tmp | (~ cfg_nan_to_zero))
      & (else_mux_29_tmp[3]);
  assign or_dcpl_555 = (else_mux_29_tmp[3:0]!=4'b1111) | ((~ IsNaN_5U_10U_nor_9_tmp)
      & cfg_nan_to_zero) | (~ (else_mux_29_tmp[4])) | IsNaN_5U_23U_nor_9_tmp;
  assign and_dcpl_1220 = and_dcpl_1214 & and_dcpl_1211 & (else_mux_29_tmp[4]) & (~
      IsNaN_5U_23U_nor_9_tmp);
  assign and_dcpl_1221 = or_dcpl_555 & and_dcpl_638;
  assign or_dcpl_567 = (~ cfg_nan_to_zero) | IsNaN_5U_10U_nor_10_tmp;
  assign or_dcpl_573 = (else_mux_32_tmp!=5'b11111) | IsNaN_5U_23U_nor_10_tmp | (cfg_nan_to_zero
      & (~ IsNaN_5U_10U_nor_10_tmp));
  assign and_dcpl_1238 = and_dcpl_638 & (else_mux_32_tmp==5'b11111) & (~ IsNaN_5U_23U_nor_10_tmp)
      & or_dcpl_567;
  assign and_dcpl_1239 = or_dcpl_573 & and_dcpl_638;
  assign or_dcpl_585 = IsNaN_5U_10U_nor_11_tmp | (~ cfg_nan_to_zero);
  assign or_dcpl_591 = (else_mux_35_tmp!=5'b11111) | IsNaN_5U_23U_nor_11_tmp | ((~
      IsNaN_5U_10U_nor_11_tmp) & cfg_nan_to_zero);
  assign and_dcpl_1256 = and_dcpl_638 & (else_mux_35_tmp==5'b11111) & (~ IsNaN_5U_23U_nor_11_tmp)
      & or_dcpl_585;
  assign and_dcpl_1257 = or_dcpl_591 & and_dcpl_638;
  assign or_dcpl_603 = IsNaN_5U_10U_nor_12_tmp | (~ cfg_nan_to_zero);
  assign or_dcpl_609 = (else_mux_38_tmp!=5'b11111) | IsNaN_5U_23U_nor_12_tmp | ((~
      IsNaN_5U_10U_nor_12_tmp) & cfg_nan_to_zero);
  assign and_dcpl_1274 = and_dcpl_638 & (else_mux_38_tmp==5'b11111) & (~ IsNaN_5U_23U_nor_12_tmp)
      & or_dcpl_603;
  assign and_dcpl_1275 = or_dcpl_609 & and_dcpl_638;
  assign and_dcpl_1279 = (else_mux_41_tmp[3:1]==3'b111);
  assign and_dcpl_1283 = (~((~(IsNaN_5U_10U_nor_13_tmp | (~ cfg_nan_to_zero))) |
      io_read_cfg_alu_bypass_rsc_svs_st_1)) & and_dcpl_21 & (else_mux_41_tmp[4]);
  assign or_dcpl_627 = ((~ IsNaN_5U_10U_nor_13_tmp) & cfg_nan_to_zero) | (else_mux_41_tmp!=5'b11111)
      | IsNaN_5U_23U_nor_13_tmp;
  assign and_dcpl_1289 = and_dcpl_1283 & and_dcpl_1279 & (else_mux_41_tmp[0]) & (~
      IsNaN_5U_23U_nor_13_tmp);
  assign and_dcpl_1290 = or_dcpl_627 & and_dcpl_638;
  assign or_dcpl_639 = (~ cfg_nan_to_zero) | IsNaN_5U_10U_nor_14_tmp;
  assign or_dcpl_645 = (else_mux_44_tmp!=5'b11111) | IsNaN_5U_23U_nor_14_tmp | (cfg_nan_to_zero
      & (~ IsNaN_5U_10U_nor_14_tmp));
  assign and_dcpl_1307 = and_dcpl_638 & (else_mux_44_tmp==5'b11111) & (~ IsNaN_5U_23U_nor_14_tmp)
      & or_dcpl_639;
  assign and_dcpl_1308 = or_dcpl_645 & and_dcpl_638;
  assign or_dcpl_657 = IsNaN_5U_10U_nor_15_tmp | (~ cfg_nan_to_zero);
  assign or_dcpl_663 = (else_mux_47_tmp!=5'b11111) | IsNaN_5U_23U_nor_15_tmp | ((~
      IsNaN_5U_10U_nor_15_tmp) & cfg_nan_to_zero);
  assign and_dcpl_1325 = and_dcpl_638 & (else_mux_47_tmp==5'b11111) & (~ IsNaN_5U_23U_nor_15_tmp)
      & or_dcpl_657;
  assign and_dcpl_1326 = or_dcpl_663 & and_dcpl_638;
  assign or_dcpl_675 = or_22_cse | or_dcpl_3;
  assign and_dcpl_1329 = and_dcpl_21 & main_stage_v_2;
  assign and_dcpl_1333 = and_dcpl_21 & main_stage_v_2 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5);
  assign and_dcpl_1335 = and_dcpl_406 & and_dcpl_1333 & and_dcpl_404;
  assign and_dcpl_1341 = and_dcpl_421 & and_dcpl_1333 & and_dcpl_419;
  assign and_dcpl_1347 = and_dcpl_436 & and_dcpl_1333 & and_dcpl_434;
  assign and_dcpl_1353 = and_dcpl_451 & and_dcpl_1333 & and_dcpl_449;
  assign and_dcpl_1359 = and_dcpl_569 & and_dcpl_1333 & and_dcpl_567;
  assign and_dcpl_1365 = and_dcpl_580 & and_dcpl_1333 & and_dcpl_578;
  assign and_dcpl_1371 = and_dcpl_591 & and_dcpl_1333 & and_dcpl_589;
  assign and_dcpl_1377 = and_dcpl_478 & and_dcpl_1333 & and_dcpl_476;
  assign and_dcpl_1383 = and_dcpl_602 & and_dcpl_1333 & and_dcpl_600;
  assign and_dcpl_1389 = and_dcpl_613 & and_dcpl_1333 & and_dcpl_611;
  assign and_dcpl_1395 = and_dcpl_624 & and_dcpl_1333 & and_dcpl_622;
  assign and_dcpl_1401 = and_dcpl_635 & and_dcpl_1333 & and_dcpl_633;
  assign and_dcpl_1407 = and_dcpl_509 & and_dcpl_1333 & and_dcpl_507;
  assign and_dcpl_1413 = and_dcpl_524 & and_dcpl_1333 & and_dcpl_522;
  assign and_dcpl_1419 = and_dcpl_539 & and_dcpl_1333 & and_dcpl_537;
  assign and_dcpl_1425 = and_dcpl_554 & and_dcpl_1333 & and_dcpl_552;
  assign or_dcpl_677 = or_22_cse | (~ main_stage_v_2);
  assign or_dcpl_678 = or_dcpl_677 | and_dcpl_7 | io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign and_dcpl_1426 = (cfg_alu_algo_1_sva_st_92==2'b10);
  assign or_dcpl_679 = or_dcpl_295 | IsNaN_8U_23U_2_land_lpi_1_dfm_st_1;
  assign or_dcpl_681 = or_dcpl_295 | IsNaN_8U_23U_2_land_15_lpi_1_dfm_st_1;
  assign or_dcpl_683 = or_dcpl_295 | IsNaN_8U_23U_2_land_14_lpi_1_dfm_st_1;
  assign or_dcpl_686 = (cfg_alu_algo_1_sva_st_92!=2'b10) | IsNaN_8U_23U_2_land_13_lpi_1_dfm_st_1;
  assign or_dcpl_688 = or_dcpl_295 | IsNaN_8U_23U_2_land_11_lpi_1_dfm_st_1;
  assign or_dcpl_692 = or_dcpl_295 | IsNaN_8U_23U_2_land_7_lpi_1_dfm_st_1;
  assign or_dcpl_694 = or_dcpl_295 | IsNaN_8U_23U_2_land_5_lpi_1_dfm_st_1;
  assign or_dcpl_696 = or_dcpl_295 | IsNaN_8U_23U_2_land_3_lpi_1_dfm_st_1;
  assign or_dcpl_699 = (cfg_alu_algo_1_sva_st_92[0]) | IsNaN_8U_23U_2_land_1_lpi_1_dfm_st_1
      | (~ (cfg_alu_algo_1_sva_st_92[1]));
  assign and_dcpl_1468 = ~((reg_cfg_alu_algo_1_sva_st_157_cse!=2'b00));
  assign and_dcpl_1471 = or_22_cse & main_stage_v_2;
  assign and_dcpl_1472 = and_dcpl_1471 & or_cse_2;
  assign and_dcpl_1476 = and_dcpl_1472 & (~(io_read_cfg_alu_bypass_rsc_svs_st_5 |
      alu_loop_op_1_else_if_acc_itm_32_1)) & and_dcpl_1468;
  assign and_dcpl_1477 = (reg_cfg_alu_algo_1_sva_st_157_cse==2'b01);
  assign and_dcpl_1483 = and_dcpl_1472 & (~(io_read_cfg_alu_bypass_rsc_svs_st_5 |
      alu_loop_op_1_else_else_if_acc_itm_32_1)) & and_dcpl_1477;
  assign and_dcpl_1490 = and_dcpl_1472 & (~(io_read_cfg_alu_bypass_rsc_svs_st_5 |
      alu_loop_op_2_else_if_acc_1_itm_32_1)) & and_dcpl_1468;
  assign and_dcpl_1497 = and_dcpl_1472 & (~(io_read_cfg_alu_bypass_rsc_svs_st_5 |
      alu_loop_op_2_else_else_if_acc_1_itm_32_1)) & and_dcpl_1477;
  assign and_dcpl_1504 = and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & (~ alu_loop_op_3_else_if_acc_itm_32_1) & and_dcpl_1468;
  assign and_dcpl_1511 = and_dcpl_1472 & (~(io_read_cfg_alu_bypass_rsc_svs_st_5 |
      alu_loop_op_3_else_else_if_acc_itm_32_1)) & and_dcpl_1477;
  assign and_dcpl_1518 = and_dcpl_1472 & (~(io_read_cfg_alu_bypass_rsc_svs_st_5 |
      alu_loop_op_4_else_if_acc_1_itm_32_1)) & and_dcpl_1468;
  assign and_dcpl_1525 = and_dcpl_1472 & (~(io_read_cfg_alu_bypass_rsc_svs_st_5 |
      alu_loop_op_4_else_else_if_acc_1_itm_32_1)) & and_dcpl_1477;
  assign and_dcpl_1532 = and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & (~ alu_loop_op_5_else_if_acc_itm_32_1) & and_dcpl_1468;
  assign and_dcpl_1539 = and_dcpl_1472 & (~(io_read_cfg_alu_bypass_rsc_svs_st_5 |
      alu_loop_op_5_else_else_if_acc_itm_32_1)) & and_dcpl_1477;
  assign and_dcpl_1546 = and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & (~ alu_loop_op_6_else_if_acc_1_itm_32_1) & and_dcpl_1468;
  assign and_dcpl_1553 = and_dcpl_1472 & (~(io_read_cfg_alu_bypass_rsc_svs_st_5 |
      alu_loop_op_6_else_else_if_acc_1_itm_32_1)) & and_dcpl_1477;
  assign and_dcpl_1560 = and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & (~ alu_loop_op_7_else_if_acc_itm_32_1) & and_dcpl_1468;
  assign and_dcpl_1567 = and_dcpl_1472 & (~(io_read_cfg_alu_bypass_rsc_svs_st_5 |
      alu_loop_op_7_else_else_if_acc_itm_32_1)) & and_dcpl_1477;
  assign and_dcpl_1574 = and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & (~ alu_loop_op_8_else_if_acc_1_itm_32_1) & and_dcpl_1468;
  assign and_dcpl_1581 = and_dcpl_1472 & (~(io_read_cfg_alu_bypass_rsc_svs_st_5 |
      alu_loop_op_8_else_else_if_acc_1_itm_32_1)) & and_dcpl_1477;
  assign and_dcpl_1588 = and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & (~ alu_loop_op_9_else_if_acc_itm_32_1) & and_dcpl_1468;
  assign and_dcpl_1595 = and_dcpl_1472 & (~(io_read_cfg_alu_bypass_rsc_svs_st_5 |
      alu_loop_op_9_else_else_if_acc_itm_32_1)) & and_dcpl_1477;
  assign and_dcpl_1602 = and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & (~ alu_loop_op_10_else_if_acc_1_itm_32_1) & and_dcpl_1468;
  assign and_dcpl_1609 = and_dcpl_1472 & (~(io_read_cfg_alu_bypass_rsc_svs_st_5 |
      alu_loop_op_10_else_else_if_acc_1_itm_32_1)) & and_dcpl_1477;
  assign and_dcpl_1616 = and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & (~ alu_loop_op_11_else_if_acc_itm_32_1) & and_dcpl_1468;
  assign and_dcpl_1623 = and_dcpl_1472 & (~(io_read_cfg_alu_bypass_rsc_svs_st_5 |
      alu_loop_op_11_else_else_if_acc_itm_32_1)) & and_dcpl_1477;
  assign and_dcpl_1630 = and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & (~ alu_loop_op_12_else_if_acc_1_itm_32_1) & and_dcpl_1468;
  assign and_dcpl_1637 = and_dcpl_1472 & (~(io_read_cfg_alu_bypass_rsc_svs_st_5 |
      alu_loop_op_12_else_else_if_acc_1_itm_32_1)) & and_dcpl_1477;
  assign and_dcpl_1644 = and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & (~ alu_loop_op_13_else_if_acc_itm_32_1) & and_dcpl_1468;
  assign and_dcpl_1651 = and_dcpl_1472 & (~(io_read_cfg_alu_bypass_rsc_svs_st_5 |
      alu_loop_op_13_else_else_if_acc_itm_32_1)) & and_dcpl_1477;
  assign and_dcpl_1658 = and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & (~ alu_loop_op_14_else_if_acc_1_itm_32_1) & and_dcpl_1468;
  assign and_dcpl_1665 = and_dcpl_1472 & (~(io_read_cfg_alu_bypass_rsc_svs_st_5 |
      alu_loop_op_14_else_else_if_acc_1_itm_32_1)) & and_dcpl_1477;
  assign and_dcpl_1672 = and_dcpl_1472 & (~ io_read_cfg_alu_bypass_rsc_svs_st_5)
      & (~ alu_loop_op_15_else_if_acc_itm_32_1) & and_dcpl_1468;
  assign and_dcpl_1679 = and_dcpl_1472 & (~(io_read_cfg_alu_bypass_rsc_svs_st_5 |
      alu_loop_op_15_else_else_if_acc_itm_32_1)) & and_dcpl_1477;
  assign and_dcpl_1682 = and_dcpl_1471 & and_dcpl_695;
  assign and_dcpl_1686 = and_dcpl_1682 & (~ (reg_cfg_alu_algo_1_sva_st_157_cse[0]))
      & (~ alu_loop_op_16_else_if_acc_1_itm_32_1) & or_cse_2;
  assign and_dcpl_1691 = and_dcpl_1682 & (reg_cfg_alu_algo_1_sva_st_157_cse[0]) &
      (~ alu_loop_op_16_else_else_if_acc_1_itm_32_1) & or_cse_2;
  assign and_dcpl_1692 = (cfg_alu_algo_1_sva_st_92[1]) & and_89_tmp;
  assign or_dcpl_775 = (cfg_alu_algo_1_sva_st_92[0]) | IsNaN_8U_23U_2_land_10_lpi_1_dfm_st_1
      | (~ (cfg_alu_algo_1_sva_st_92[1]));
  assign or_dcpl_777 = or_dcpl_295 | IsNaN_8U_23U_2_land_9_lpi_1_dfm_st_1;
  assign or_dcpl_780 = (cfg_alu_algo_1_sva_st_92!=2'b10) | IsNaN_8U_23U_2_land_6_lpi_1_dfm_st_1;
  assign or_dcpl_783 = (cfg_alu_algo_1_sva_st_92!=2'b10) | IsNaN_8U_23U_2_land_4_lpi_1_dfm_st_1;
  assign or_dcpl_785 = or_dcpl_295 | IsNaN_8U_23U_2_land_2_lpi_1_dfm_st_1;
  assign or_dcpl_787 = alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_st_2 | (reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign or_dcpl_790 = or_dcpl_677 | and_dcpl_7;
  assign or_dcpl_823 = alu_loop_op_6_FpCmp_8U_23U_false_slc_8_1_svs_st_2 | (reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign or_dcpl_830 = (reg_cfg_alu_algo_1_sva_st_93_cse[1]) | alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_st_2;
  assign or_dcpl_837 = alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_st_2 | (reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign or_dcpl_844 = alu_loop_op_9_FpCmp_8U_23U_false_slc_8_svs_st_2 | (reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign or_dcpl_851 = alu_loop_op_10_FpCmp_8U_23U_false_slc_8_1_svs_st_2 | (reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign or_dcpl_859 = io_read_cfg_alu_bypass_rsc_svs_st_5 | (reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign or_dcpl_872 = alu_loop_op_13_FpCmp_8U_23U_false_slc_8_svs_st_2 | (reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign or_dcpl_879 = alu_loop_op_14_FpCmp_8U_23U_false_slc_8_1_svs_st_2 | (reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign or_dcpl_893 = alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_st_2 | (reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign or_dcpl_901 = or_22_cse | (cfg_alu_algo_rsci_d[0]);
  assign or_tmp_3044 = and_91_tmp & (fsm_output[1]);
  assign or_tmp_3045 = and_dcpl_11 & cfg_alu_src_rsci_d & (fsm_output[1]);
  assign or_tmp_3048 = and_89_tmp & (fsm_output[1]);
  assign or_tmp_3190 = or_dcpl_391 & and_dcpl_29 & (fsm_output[1]);
  assign or_tmp_3201 = or_dcpl_411 & and_dcpl_29 & (fsm_output[1]);
  assign or_tmp_3212 = or_dcpl_429 & and_dcpl_29 & (fsm_output[1]);
  assign or_tmp_3223 = or_dcpl_447 & and_dcpl_29 & (fsm_output[1]);
  assign or_tmp_3234 = or_dcpl_465 & and_dcpl_29 & (fsm_output[1]);
  assign or_tmp_3245 = or_dcpl_483 & and_dcpl_29 & (fsm_output[1]);
  assign or_tmp_3256 = or_dcpl_501 & and_dcpl_29 & (fsm_output[1]);
  assign or_tmp_3267 = or_dcpl_519 & and_dcpl_29 & (fsm_output[1]);
  assign or_tmp_3278 = or_dcpl_537 & and_dcpl_29 & (fsm_output[1]);
  assign or_tmp_3289 = or_dcpl_555 & and_dcpl_29 & (fsm_output[1]);
  assign or_tmp_3300 = or_dcpl_573 & and_dcpl_29 & (fsm_output[1]);
  assign or_tmp_3311 = or_dcpl_591 & and_dcpl_29 & (fsm_output[1]);
  assign or_tmp_3322 = or_dcpl_609 & and_dcpl_29 & (fsm_output[1]);
  assign or_tmp_3333 = or_dcpl_627 & and_dcpl_29 & (fsm_output[1]);
  assign or_tmp_3344 = or_dcpl_645 & and_dcpl_29 & (fsm_output[1]);
  assign or_tmp_3355 = or_dcpl_663 & and_dcpl_29 & (fsm_output[1]);
  assign or_tmp_3479 = (or_dcpl_901 | (~ (cfg_alu_algo_rsci_d[1])) | cfg_alu_bypass_rsci_d)
      & and_91_tmp & (fsm_output[1]);
  assign chn_alu_in_rsci_ld_core_psct_mx0c0 = and_91_tmp | (fsm_output[0]);
  assign chn_alu_op_rsci_ld_core_psct_mx0c1 = and_dcpl_14 & (or_dcpl_3 | (~ cfg_alu_src_rsci_d));
  assign main_stage_v_2_mx0c1 = or_cse_2 & main_stage_v_2 & (~ and_89_tmp);
  assign main_stage_v_3_mx0c1 = (~ main_stage_v_2) & main_stage_v_3 & or_cse_2;
  assign main_stage_v_4_mx0c1 = (~ main_stage_v_3) & main_stage_v_4 & or_cse_2;
  assign main_stage_v_1_mx0c1 = (~ and_91_tmp) & and_89_tmp & (fsm_output[1]);
  assign cfg_alu_src_1_sva_st_1_mx0c1 = and_91_tmp & cfg_alu_bypass_rsci_d & (fsm_output[1]);
  assign chn_alu_in_rsci_oswt_unreg = or_tmp_3044;
  assign chn_alu_op_rsci_oswt_unreg = and_dcpl_14;
  assign chn_alu_out_rsci_oswt_unreg = chn_alu_out_rsci_bawt & reg_chn_alu_out_rsci_ld_core_psct_cse;
  assign cfg_alu_op_rsc_triosy_obj_oswt_unreg_pff = or_tmp_3048;
  assign and_dcpl_1789 = nor_7_ssc & (~ FpAlu_8U_23U_equal_tmp_237);
  assign or_dcpl_1047 = (((FpAlu_8U_23U_nor_dfs_79 & IsNaN_8U_23U_land_1_lpi_1_dfm_10)
      | reg_FpAlu_8U_23U_or_752_cse) & and_dcpl_1789) | io_read_cfg_alu_bypass_rsc_svs_7;
  assign and_dcpl_1796 = FpAlu_8U_23U_or_863_cse & and_dcpl_1789;
  assign or_dcpl_1052 = (((FpAlu_8U_23U_nor_dfs_79 & IsNaN_8U_23U_land_2_lpi_1_dfm_10)
      | reg_FpAlu_8U_23U_or_755_cse) & and_dcpl_1789) | io_read_cfg_alu_bypass_rsc_svs_7;
  assign and_dcpl_1804 = FpAlu_8U_23U_or_864_cse & and_dcpl_1789;
  assign or_dcpl_1057 = (((FpAlu_8U_23U_nor_dfs_79 & IsNaN_8U_23U_land_3_lpi_1_dfm_10)
      | reg_FpAlu_8U_23U_or_758_cse) & and_dcpl_1789) | io_read_cfg_alu_bypass_rsc_svs_7;
  assign and_dcpl_1812 = FpAlu_8U_23U_or_865_cse & and_dcpl_1789;
  assign or_dcpl_1062 = (((FpAlu_8U_23U_nor_dfs_79 & IsNaN_8U_23U_land_4_lpi_1_dfm_10)
      | reg_FpAlu_8U_23U_or_761_cse) & and_dcpl_1789) | io_read_cfg_alu_bypass_rsc_svs_7;
  assign and_dcpl_1820 = FpAlu_8U_23U_or_866_cse & and_dcpl_1789;
  assign or_dcpl_1067 = (((FpAlu_8U_23U_nor_dfs_79 & IsNaN_8U_23U_land_5_lpi_1_dfm_10)
      | reg_FpAlu_8U_23U_or_764_cse) & and_dcpl_1789) | io_read_cfg_alu_bypass_rsc_svs_7;
  assign and_dcpl_1828 = FpAlu_8U_23U_or_867_cse & and_dcpl_1789;
  assign or_dcpl_1072 = (((FpAlu_8U_23U_nor_dfs_79 & IsNaN_8U_23U_land_6_lpi_1_dfm_10)
      | reg_FpAlu_8U_23U_or_767_cse) & and_dcpl_1789) | io_read_cfg_alu_bypass_rsc_svs_7;
  assign and_dcpl_1836 = FpAlu_8U_23U_or_868_cse & and_dcpl_1789;
  assign or_dcpl_1077 = (((FpAlu_8U_23U_nor_dfs_79 & IsNaN_8U_23U_land_7_lpi_1_dfm_10)
      | reg_FpAlu_8U_23U_or_770_cse) & and_dcpl_1789) | io_read_cfg_alu_bypass_rsc_svs_7;
  assign and_dcpl_1844 = FpAlu_8U_23U_or_869_cse & and_dcpl_1789;
  assign or_dcpl_1082 = (((FpAlu_8U_23U_nor_dfs_79 & IsNaN_8U_23U_land_8_lpi_1_dfm_10)
      | reg_FpAlu_8U_23U_or_773_cse) & and_dcpl_1789) | io_read_cfg_alu_bypass_rsc_svs_7;
  assign and_dcpl_1852 = FpAlu_8U_23U_or_870_cse & and_dcpl_1789;
  assign or_dcpl_1087 = (((FpAlu_8U_23U_nor_dfs_79 & IsNaN_8U_23U_land_9_lpi_1_dfm_10)
      | reg_FpAlu_8U_23U_or_776_cse) & and_dcpl_1789) | io_read_cfg_alu_bypass_rsc_svs_7;
  assign and_dcpl_1860 = FpAlu_8U_23U_or_871_cse & and_dcpl_1789;
  assign or_dcpl_1092 = (((FpAlu_8U_23U_nor_dfs_79 & IsNaN_8U_23U_land_10_lpi_1_dfm_10)
      | reg_FpAlu_8U_23U_or_779_cse) & and_dcpl_1789) | io_read_cfg_alu_bypass_rsc_svs_7;
  assign and_dcpl_1868 = FpAlu_8U_23U_or_872_cse & and_dcpl_1789;
  assign or_dcpl_1097 = (((FpAlu_8U_23U_nor_dfs_79 & IsNaN_8U_23U_land_11_lpi_1_dfm_10)
      | reg_FpAlu_8U_23U_or_782_cse) & and_dcpl_1789) | io_read_cfg_alu_bypass_rsc_svs_7;
  assign and_dcpl_1876 = FpAlu_8U_23U_or_873_cse & and_dcpl_1789;
  assign or_dcpl_1102 = (((FpAlu_8U_23U_nor_dfs_79 & IsNaN_8U_23U_land_12_lpi_1_dfm_10)
      | reg_FpAlu_8U_23U_or_785_cse) & and_dcpl_1789) | io_read_cfg_alu_bypass_rsc_svs_7;
  assign and_dcpl_1884 = FpAlu_8U_23U_or_874_cse & and_dcpl_1789;
  assign or_dcpl_1107 = (((FpAlu_8U_23U_nor_dfs_79 & IsNaN_8U_23U_land_13_lpi_1_dfm_10)
      | reg_FpAlu_8U_23U_or_788_cse) & and_dcpl_1789) | io_read_cfg_alu_bypass_rsc_svs_7;
  assign and_dcpl_1892 = FpAlu_8U_23U_or_875_cse & and_dcpl_1789;
  assign or_dcpl_1112 = (((FpAlu_8U_23U_nor_dfs_79 & IsNaN_8U_23U_land_14_lpi_1_dfm_10)
      | reg_FpAlu_8U_23U_or_791_cse) & and_dcpl_1789) | io_read_cfg_alu_bypass_rsc_svs_7;
  assign and_dcpl_1900 = FpAlu_8U_23U_or_876_cse & and_dcpl_1789;
  assign or_dcpl_1117 = (((FpAlu_8U_23U_nor_dfs_79 & IsNaN_8U_23U_land_15_lpi_1_dfm_10)
      | reg_FpAlu_8U_23U_or_794_cse) & and_dcpl_1789) | io_read_cfg_alu_bypass_rsc_svs_7;
  assign and_dcpl_1908 = FpAlu_8U_23U_or_877_cse & and_dcpl_1789;
  assign or_dcpl_1122 = (((FpAlu_8U_23U_nor_dfs_79 & IsNaN_8U_23U_land_lpi_1_dfm_10)
      | reg_FpAlu_8U_23U_or_797_cse) & and_dcpl_1789) | io_read_cfg_alu_bypass_rsc_svs_7;
  assign and_dcpl_1916 = FpAlu_8U_23U_or_878_cse & and_dcpl_1789;
  assign FpNormalize_8U_49U_else_and_tmp = (fsm_output[1]) & (~ (FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49]));
  assign FpNormalize_8U_49U_else_and_tmp_1 = (fsm_output[1]) & (~ (FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49]));
  assign FpNormalize_8U_49U_else_and_tmp_2 = (fsm_output[1]) & (~ (FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49]));
  assign FpNormalize_8U_49U_else_and_tmp_3 = (fsm_output[1]) & (~ (FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_5[49]));
  assign FpNormalize_8U_49U_else_and_tmp_4 = (fsm_output[1]) & (~ (FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_5[49]));
  assign FpNormalize_8U_49U_else_and_tmp_5 = (fsm_output[1]) & (~ (FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_5[49]));
  assign FpNormalize_8U_49U_else_and_tmp_6 = (fsm_output[1]) & (~ (FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_5[49]));
  assign FpNormalize_8U_49U_else_and_tmp_7 = (fsm_output[1]) & (~ (FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_5[49]));
  assign FpNormalize_8U_49U_else_and_tmp_8 = (fsm_output[1]) & (~ (FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_5[49]));
  assign FpNormalize_8U_49U_else_and_tmp_9 = (fsm_output[1]) & (~ (FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_5[49]));
  assign FpNormalize_8U_49U_else_and_tmp_10 = (fsm_output[1]) & (~ (FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_5[49]));
  assign FpNormalize_8U_49U_else_and_tmp_11 = (fsm_output[1]) & (~ (FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_5[49]));
  assign FpNormalize_8U_49U_else_and_tmp_12 = (fsm_output[1]) & (~ (FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_5[49]));
  assign FpNormalize_8U_49U_else_and_tmp_13 = (fsm_output[1]) & (~ (FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_5[49]));
  assign FpNormalize_8U_49U_else_and_tmp_14 = (fsm_output[1]) & (~ (FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_5[49]));
  assign FpNormalize_8U_49U_else_and_tmp_15 = (fsm_output[1]) & (~ (FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49]));
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp = (fsm_output[1]) & (~((~((~ alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2)
      | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_itm_23_1)) | alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_2));
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_1 = (fsm_output[1]) & (~((~((~
      alu_loop_op_16_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2) | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_15_itm_23_1))
      | alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_2));
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_2 = (fsm_output[1]) & (~((~((~
      alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2) | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_itm_23_1))
      | alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_2));
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_3 = (fsm_output[1]) & (~((~((~
      alu_loop_op_15_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2) | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_14_itm_23_1))
      | alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_2));
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_4 = (fsm_output[1]) & (~((~((~
      alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2) | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_itm_23_1))
      | alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_2));
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_5 = (fsm_output[1]) & (~((~((~
      alu_loop_op_14_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2) | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_13_itm_23_1))
      | alu_loop_op_14_FpCmp_8U_23U_false_slc_8_1_svs_2));
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_6 = (fsm_output[1]) & (~((~((~
      alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2) | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_itm_23_1))
      | alu_loop_op_4_FpCmp_8U_23U_false_slc_8_1_svs_2));
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_7 = (fsm_output[1]) & (~((~((~
      alu_loop_op_13_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2) | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_12_itm_23_1))
      | alu_loop_op_13_FpCmp_8U_23U_false_slc_8_svs_2));
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_8 = (fsm_output[1]) & (~((~((~
      alu_loop_op_5_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2) | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_itm_23_1))
      | alu_loop_op_5_FpCmp_8U_23U_false_slc_8_svs_2));
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_9 = (fsm_output[1]) & (~((~((~
      alu_loop_op_12_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2) | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_11_itm_23_1))
      | alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_2));
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_10 = (fsm_output[1]) & (~((~((~
      alu_loop_op_6_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2) | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_5_itm_23_1))
      | alu_loop_op_6_FpCmp_8U_23U_false_slc_8_1_svs_2));
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_11 = (fsm_output[1]) & (~((~((~
      alu_loop_op_11_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2) | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_itm_23_1))
      | alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_2));
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_12 = (fsm_output[1]) & (~((~((~
      alu_loop_op_7_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2) | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_itm_23_1))
      | alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_2));
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_13 = (fsm_output[1]) & (~((~((~
      alu_loop_op_10_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2) | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_9_itm_23_1))
      | alu_loop_op_10_FpCmp_8U_23U_false_slc_8_1_svs_2));
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_14 = (fsm_output[1]) & (~((~((~
      alu_loop_op_8_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2) | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_7_itm_23_1))
      | alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_2));
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_15 = (fsm_output[1]) & (~((~((~
      alu_loop_op_9_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2) | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_itm_23_1))
      | alu_loop_op_9_FpCmp_8U_23U_false_slc_8_svs_2));
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_in_rsci_iswt0 <= 1'b0;
      reg_cfg_alu_shift_value_rsc_triosy_obj_ld_core_psct_cse <= 1'b0;
      chn_alu_out_rsci_iswt0 <= 1'b0;
      chn_alu_op_rsci_iswt0 <= 1'b0;
    end
    else if ( core_wen ) begin
      chn_alu_in_rsci_iswt0 <= ~((~ and_91_tmp) & (fsm_output[1]));
      reg_cfg_alu_shift_value_rsc_triosy_obj_ld_core_psct_cse <= or_tmp_3044;
      chn_alu_out_rsci_iswt0 <= and_dcpl_8;
      chn_alu_op_rsci_iswt0 <= or_tmp_3045;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_in_rsci_ld_core_psct <= 1'b0;
    end
    else if ( core_wen & chn_alu_in_rsci_ld_core_psct_mx0c0 ) begin
      chn_alu_in_rsci_ld_core_psct <= chn_alu_in_rsci_ld_core_psct_mx0c0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_0 <= 1'b0;
      chn_alu_out_rsci_d_22_1 <= 22'b0;
      chn_alu_out_rsci_d_30_27 <= 4'b0;
      chn_alu_out_rsci_d_32_31 <= 2'b0;
      chn_alu_out_rsci_d_33 <= 1'b0;
      chn_alu_out_rsci_d_55_34 <= 22'b0;
      chn_alu_out_rsci_d_63_60 <= 4'b0;
      chn_alu_out_rsci_d_65_64 <= 2'b0;
      chn_alu_out_rsci_d_66 <= 1'b0;
      chn_alu_out_rsci_d_88_67 <= 22'b0;
      chn_alu_out_rsci_d_96_93 <= 4'b0;
      chn_alu_out_rsci_d_98_97 <= 2'b0;
      chn_alu_out_rsci_d_99 <= 1'b0;
      chn_alu_out_rsci_d_121_100 <= 22'b0;
      chn_alu_out_rsci_d_129_126 <= 4'b0;
      chn_alu_out_rsci_d_131_130 <= 2'b0;
      chn_alu_out_rsci_d_132 <= 1'b0;
      chn_alu_out_rsci_d_154_133 <= 22'b0;
      chn_alu_out_rsci_d_162_159 <= 4'b0;
      chn_alu_out_rsci_d_164_163 <= 2'b0;
      chn_alu_out_rsci_d_165 <= 1'b0;
      chn_alu_out_rsci_d_187_166 <= 22'b0;
      chn_alu_out_rsci_d_195_192 <= 4'b0;
      chn_alu_out_rsci_d_197_196 <= 2'b0;
      chn_alu_out_rsci_d_198 <= 1'b0;
      chn_alu_out_rsci_d_220_199 <= 22'b0;
      chn_alu_out_rsci_d_228_225 <= 4'b0;
      chn_alu_out_rsci_d_230_229 <= 2'b0;
      chn_alu_out_rsci_d_231 <= 1'b0;
      chn_alu_out_rsci_d_253_232 <= 22'b0;
      chn_alu_out_rsci_d_261_258 <= 4'b0;
      chn_alu_out_rsci_d_263_262 <= 2'b0;
      chn_alu_out_rsci_d_264 <= 1'b0;
      chn_alu_out_rsci_d_286_265 <= 22'b0;
      chn_alu_out_rsci_d_294_291 <= 4'b0;
      chn_alu_out_rsci_d_296_295 <= 2'b0;
      chn_alu_out_rsci_d_297 <= 1'b0;
      chn_alu_out_rsci_d_319_298 <= 22'b0;
      chn_alu_out_rsci_d_327_324 <= 4'b0;
      chn_alu_out_rsci_d_329_328 <= 2'b0;
      chn_alu_out_rsci_d_330 <= 1'b0;
      chn_alu_out_rsci_d_352_331 <= 22'b0;
      chn_alu_out_rsci_d_360_357 <= 4'b0;
      chn_alu_out_rsci_d_362_361 <= 2'b0;
      chn_alu_out_rsci_d_363 <= 1'b0;
      chn_alu_out_rsci_d_385_364 <= 22'b0;
      chn_alu_out_rsci_d_393_390 <= 4'b0;
      chn_alu_out_rsci_d_395_394 <= 2'b0;
      chn_alu_out_rsci_d_396 <= 1'b0;
      chn_alu_out_rsci_d_418_397 <= 22'b0;
      chn_alu_out_rsci_d_426_423 <= 4'b0;
      chn_alu_out_rsci_d_428_427 <= 2'b0;
      chn_alu_out_rsci_d_429 <= 1'b0;
      chn_alu_out_rsci_d_451_430 <= 22'b0;
      chn_alu_out_rsci_d_459_456 <= 4'b0;
      chn_alu_out_rsci_d_461_460 <= 2'b0;
      chn_alu_out_rsci_d_462 <= 1'b0;
      chn_alu_out_rsci_d_484_463 <= 22'b0;
      chn_alu_out_rsci_d_492_489 <= 4'b0;
      chn_alu_out_rsci_d_494_493 <= 2'b0;
      chn_alu_out_rsci_d_495 <= 1'b0;
      chn_alu_out_rsci_d_517_496 <= 22'b0;
      chn_alu_out_rsci_d_525_522 <= 4'b0;
      chn_alu_out_rsci_d_527_526 <= 2'b0;
    end
    else if ( chn_alu_out_and_cse ) begin
      chn_alu_out_rsci_d_0 <= MUX1HOT_s_1_7_2((FpAdd_8U_23U_o_mant_1_lpi_1_dfm_2_mx0[0]),
          (FpCmp_8U_23U_true_o_22_0_1_lpi_1_dfm_6[0]), FpAlu_8U_23U_o_0_1_sva_7,
          (FpCmp_8U_23U_false_o_22_0_1_lpi_1_dfm_6[0]), alu_loop_op_1_else_else_if_conc_itm_1_0_1,
          (AluOut_data_0_sva_8[0]), (AluIn_data_sva_503[0]), {and_149_cse , and_150_cse
          , and_151_cse , and_152_cse , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_22_1 <= MUX1HOT_v_22_4_2((FpAlu_8U_23U_and_3_nl), (alu_loop_op_1_else_else_if_conc_itm_1_30_1_1[21:0]),
          (AluOut_data_0_sva_8[22:1]), (AluIn_data_sva_503[22:1]), {nor_7_ssc , or_4809_cse
          , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_30_27 <= MUX1HOT_v_4_5_2((FpAlu_8U_23U_FpAlu_8U_23U_nor_16_nl),
          (alu_loop_op_1_else_else_if_conc_itm_1_30_1_1[29:26]), (AluOut_data_0_sva_8[30:27]),
          (AluIn_data_sva_503[30:27]), FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_11,
          {(and_4125_nl) , or_4809_cse , asn_1837 , or_dcpl_1047 , and_dcpl_1796});
      chn_alu_out_rsci_d_32_31 <= MUX1HOT_v_2_4_2(({{1{FpAlu_8U_23U_and_itm_4}},
          FpAlu_8U_23U_and_itm_4}), ({{1{alu_loop_op_1_else_else_if_conc_itm_1_31_1}},
          alu_loop_op_1_else_else_if_conc_itm_1_31_1}), (AluOut_data_0_sva_8[32:31]),
          (signext_2_1(AluIn_data_sva_503[31])), {nor_7_ssc , or_4809_cse , asn_1837
          , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_33 <= MUX1HOT_s_1_7_2((FpAdd_8U_23U_o_mant_2_lpi_1_dfm_2_mx0[0]),
          (FpCmp_8U_23U_true_o_22_0_2_lpi_1_dfm_6[0]), FpAlu_8U_23U_o_0_2_sva_7,
          (FpCmp_8U_23U_false_o_22_0_2_lpi_1_dfm_6[0]), alu_loop_op_2_else_else_if_conc_1_itm_1_0_1,
          (AluOut_data_1_sva_8[0]), (AluIn_data_sva_503[32]), {and_149_cse , and_150_cse
          , and_151_cse , and_152_cse , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_55_34 <= MUX1HOT_v_22_4_2((FpAlu_8U_23U_and_7_nl), (alu_loop_op_2_else_else_if_conc_1_itm_1_30_1_1[21:0]),
          (AluOut_data_1_sva_8[22:1]), (AluIn_data_sva_503[54:33]), {nor_7_ssc ,
          or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_63_60 <= MUX1HOT_v_4_5_2((FpAlu_8U_23U_FpAlu_8U_23U_nor_15_nl),
          (alu_loop_op_2_else_else_if_conc_1_itm_1_30_1_1[29:26]), (AluOut_data_1_sva_8[30:27]),
          (AluIn_data_sva_503[62:59]), FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_11,
          {(and_4119_nl) , or_4809_cse , asn_1837 , or_dcpl_1052 , and_dcpl_1804});
      chn_alu_out_rsci_d_65_64 <= MUX1HOT_v_2_4_2(({{1{FpAlu_8U_23U_and_4_itm_4}},
          FpAlu_8U_23U_and_4_itm_4}), ({{1{alu_loop_op_2_else_else_if_conc_1_itm_1_31_1}},
          alu_loop_op_2_else_else_if_conc_1_itm_1_31_1}), (AluOut_data_1_sva_8[32:31]),
          (signext_2_1(AluIn_data_sva_503[63])), {nor_7_ssc , or_4809_cse , asn_1837
          , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_66 <= MUX1HOT_s_1_7_2((FpAdd_8U_23U_o_mant_3_lpi_1_dfm_2_mx0[0]),
          (FpCmp_8U_23U_true_o_22_0_3_lpi_1_dfm_6[0]), FpAlu_8U_23U_o_0_3_sva_7,
          (FpCmp_8U_23U_false_o_22_0_3_lpi_1_dfm_6[0]), alu_loop_op_else_else_if_mux_8_itm_4,
          (AluOut_data_2_sva_8[0]), (AluIn_data_sva_503[64]), {and_149_cse , and_150_cse
          , and_151_cse , and_152_cse , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_88_67 <= MUX1HOT_v_22_4_2((FpAlu_8U_23U_and_11_nl), (alu_loop_op_else_else_if_mux_7_itm_4[21:0]),
          (AluOut_data_2_sva_8[22:1]), (AluIn_data_sva_503[86:65]), {nor_7_ssc ,
          or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_96_93 <= MUX1HOT_v_4_5_2((FpAlu_8U_23U_FpAlu_8U_23U_nor_14_nl),
          (alu_loop_op_else_else_if_mux_7_itm_4[29:26]), (AluOut_data_2_sva_8[30:27]),
          (AluIn_data_sva_503[94:91]), FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_11,
          {(and_4113_nl) , or_4809_cse , asn_1837 , or_dcpl_1057 , and_dcpl_1812});
      chn_alu_out_rsci_d_98_97 <= MUX1HOT_v_2_4_2(({{1{FpAlu_8U_23U_and_8_itm_4}},
          FpAlu_8U_23U_and_8_itm_4}), ({{1{alu_loop_op_else_else_if_mux_6_itm_4}},
          alu_loop_op_else_else_if_mux_6_itm_4}), (AluOut_data_2_sva_8[32:31]), (signext_2_1(AluIn_data_sva_503[95])),
          {nor_7_ssc , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_99 <= MUX1HOT_s_1_7_2((FpAdd_8U_23U_o_mant_4_lpi_1_dfm_2_mx0[0]),
          (FpCmp_8U_23U_true_o_22_0_4_lpi_1_dfm_6[0]), FpAlu_8U_23U_o_0_4_sva_7,
          (FpCmp_8U_23U_false_o_22_0_4_lpi_1_dfm_6[0]), alu_loop_op_4_else_else_if_conc_1_itm_1_0_1,
          (AluOut_data_3_sva_8[0]), (AluIn_data_sva_503[96]), {and_149_cse , and_150_cse
          , and_151_cse , and_152_cse , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_121_100 <= MUX1HOT_v_22_4_2((FpAlu_8U_23U_and_15_nl), (alu_loop_op_4_else_else_if_conc_1_itm_1_30_1_1[21:0]),
          (AluOut_data_3_sva_8[22:1]), (AluIn_data_sva_503[118:97]), {nor_7_ssc ,
          or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_129_126 <= MUX1HOT_v_4_5_2((FpAlu_8U_23U_FpAlu_8U_23U_nor_13_nl),
          (alu_loop_op_4_else_else_if_conc_1_itm_1_30_1_1[29:26]), (AluOut_data_3_sva_8[30:27]),
          (AluIn_data_sva_503[126:123]), FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_11,
          {(and_4107_nl) , or_4809_cse , asn_1837 , or_dcpl_1062 , and_dcpl_1820});
      chn_alu_out_rsci_d_131_130 <= MUX1HOT_v_2_4_2(({{1{FpAlu_8U_23U_and_12_itm_4}},
          FpAlu_8U_23U_and_12_itm_4}), ({{1{alu_loop_op_4_else_else_if_conc_1_itm_1_31_1}},
          alu_loop_op_4_else_else_if_conc_1_itm_1_31_1}), (AluOut_data_3_sva_8[32:31]),
          (signext_2_1(AluIn_data_sva_503[127])), {nor_7_ssc , or_4809_cse , asn_1837
          , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_132 <= MUX1HOT_s_1_7_2((FpAdd_8U_23U_o_mant_5_lpi_1_dfm_2_mx0[0]),
          (FpCmp_8U_23U_true_o_22_0_5_lpi_1_dfm_6[0]), FpAlu_8U_23U_o_0_5_sva_7,
          (FpCmp_8U_23U_false_o_22_0_5_lpi_1_dfm_6[0]), alu_loop_op_else_else_if_mux_14_itm_4,
          (AluOut_data_4_sva_8[0]), (AluIn_data_sva_503[128]), {and_149_cse , and_150_cse
          , and_151_cse , and_152_cse , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_154_133 <= MUX1HOT_v_22_4_2((FpAlu_8U_23U_and_19_nl), (alu_loop_op_else_else_if_mux_13_itm_4[21:0]),
          (AluOut_data_4_sva_8[22:1]), (AluIn_data_sva_503[150:129]), {nor_7_ssc
          , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_162_159 <= MUX1HOT_v_4_5_2((FpAlu_8U_23U_FpAlu_8U_23U_nor_12_nl),
          (alu_loop_op_else_else_if_mux_13_itm_4[29:26]), (AluOut_data_4_sva_8[30:27]),
          (AluIn_data_sva_503[158:155]), FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_11,
          {(and_4101_nl) , or_4809_cse , asn_1837 , or_dcpl_1067 , and_dcpl_1828});
      chn_alu_out_rsci_d_164_163 <= MUX1HOT_v_2_4_2(({{1{FpAlu_8U_23U_and_16_itm_4}},
          FpAlu_8U_23U_and_16_itm_4}), ({{1{alu_loop_op_else_else_if_mux_12_itm_4}},
          alu_loop_op_else_else_if_mux_12_itm_4}), (AluOut_data_4_sva_8[32:31]),
          (signext_2_1(AluIn_data_sva_503[159])), {nor_7_ssc , or_4809_cse , asn_1837
          , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_165 <= MUX1HOT_s_1_7_2((FpAdd_8U_23U_o_mant_6_lpi_1_dfm_2_mx0[0]),
          (FpCmp_8U_23U_true_o_22_0_6_lpi_1_dfm_6[0]), FpAlu_8U_23U_o_0_6_sva_7,
          (FpCmp_8U_23U_false_o_22_0_6_lpi_1_dfm_6[0]), alu_loop_op_else_else_if_mux_17_itm_4,
          (AluOut_data_5_sva_8[0]), (AluIn_data_sva_503[160]), {and_149_cse , and_150_cse
          , and_151_cse , and_152_cse , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_187_166 <= MUX1HOT_v_22_4_2((FpAlu_8U_23U_and_23_nl), (alu_loop_op_else_else_if_mux_16_itm_4[21:0]),
          (AluOut_data_5_sva_8[22:1]), (AluIn_data_sva_503[182:161]), {nor_7_ssc
          , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_195_192 <= MUX1HOT_v_4_5_2((FpAlu_8U_23U_FpAlu_8U_23U_nor_11_nl),
          (alu_loop_op_else_else_if_mux_16_itm_4[29:26]), (AluOut_data_5_sva_8[30:27]),
          (AluIn_data_sva_503[190:187]), FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_11,
          {(and_4095_nl) , or_4809_cse , asn_1837 , or_dcpl_1072 , and_dcpl_1836});
      chn_alu_out_rsci_d_197_196 <= MUX1HOT_v_2_4_2(({{1{FpAlu_8U_23U_and_20_itm_4}},
          FpAlu_8U_23U_and_20_itm_4}), ({{1{alu_loop_op_else_else_if_mux_15_itm_4}},
          alu_loop_op_else_else_if_mux_15_itm_4}), (AluOut_data_5_sva_8[32:31]),
          (signext_2_1(AluIn_data_sva_503[191])), {nor_7_ssc , or_4809_cse , asn_1837
          , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_198 <= MUX1HOT_s_1_7_2((FpAdd_8U_23U_o_mant_7_lpi_1_dfm_2_mx0[0]),
          (FpCmp_8U_23U_true_o_22_0_7_lpi_1_dfm_6[0]), FpAlu_8U_23U_o_0_7_sva_7,
          (FpCmp_8U_23U_false_o_22_0_7_lpi_1_dfm_6[0]), alu_loop_op_else_else_if_mux_20_itm_4,
          (AluOut_data_6_sva_8[0]), (AluIn_data_sva_503[192]), {and_149_cse , and_150_cse
          , and_151_cse , and_152_cse , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_220_199 <= MUX1HOT_v_22_4_2((FpAlu_8U_23U_and_27_nl), (alu_loop_op_else_else_if_mux_19_itm_4[21:0]),
          (AluOut_data_6_sva_8[22:1]), (AluIn_data_sva_503[214:193]), {nor_7_ssc
          , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_228_225 <= MUX1HOT_v_4_5_2((FpAlu_8U_23U_FpAlu_8U_23U_nor_10_nl),
          (alu_loop_op_else_else_if_mux_19_itm_4[29:26]), (AluOut_data_6_sva_8[30:27]),
          (AluIn_data_sva_503[222:219]), FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_11,
          {(and_4089_nl) , or_4809_cse , asn_1837 , or_dcpl_1077 , and_dcpl_1844});
      chn_alu_out_rsci_d_230_229 <= MUX1HOT_v_2_4_2(({{1{FpAlu_8U_23U_and_24_itm_4}},
          FpAlu_8U_23U_and_24_itm_4}), ({{1{alu_loop_op_else_else_if_mux_18_itm_4}},
          alu_loop_op_else_else_if_mux_18_itm_4}), (AluOut_data_6_sva_8[32:31]),
          (signext_2_1(AluIn_data_sva_503[223])), {nor_7_ssc , or_4809_cse , asn_1837
          , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_231 <= MUX1HOT_s_1_7_2((FpAdd_8U_23U_o_mant_8_lpi_1_dfm_2_mx0[0]),
          (FpCmp_8U_23U_true_o_22_0_8_lpi_1_dfm_6[0]), FpAlu_8U_23U_o_0_8_sva_7,
          (FpCmp_8U_23U_false_o_22_0_8_lpi_1_dfm_6[0]), alu_loop_op_else_else_if_mux_23_itm_4,
          (AluOut_data_7_sva_8[0]), (AluIn_data_sva_503[224]), {and_149_cse , and_150_cse
          , and_151_cse , and_152_cse , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_253_232 <= MUX1HOT_v_22_4_2((FpAlu_8U_23U_and_31_nl), (alu_loop_op_else_else_if_mux_22_itm_4[21:0]),
          (AluOut_data_7_sva_8[22:1]), (AluIn_data_sva_503[246:225]), {nor_7_ssc
          , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_261_258 <= MUX1HOT_v_4_5_2((FpAlu_8U_23U_FpAlu_8U_23U_nor_9_nl),
          (alu_loop_op_else_else_if_mux_22_itm_4[29:26]), (AluOut_data_7_sva_8[30:27]),
          (AluIn_data_sva_503[254:251]), FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_11,
          {(and_4083_nl) , or_4809_cse , asn_1837 , or_dcpl_1082 , and_dcpl_1852});
      chn_alu_out_rsci_d_263_262 <= MUX1HOT_v_2_4_2(({{1{FpAlu_8U_23U_and_28_itm_4}},
          FpAlu_8U_23U_and_28_itm_4}), ({{1{alu_loop_op_else_else_if_mux_21_itm_4}},
          alu_loop_op_else_else_if_mux_21_itm_4}), (AluOut_data_7_sva_8[32:31]),
          (signext_2_1(AluIn_data_sva_503[255])), {nor_7_ssc , or_4809_cse , asn_1837
          , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_264 <= MUX1HOT_s_1_7_2((FpAdd_8U_23U_o_mant_9_lpi_1_dfm_2_mx0[0]),
          (FpCmp_8U_23U_true_o_22_0_9_lpi_1_dfm_6[0]), FpAlu_8U_23U_o_0_9_sva_7,
          (FpCmp_8U_23U_false_o_22_0_9_lpi_1_dfm_6[0]), alu_loop_op_else_else_if_mux_26_itm_4,
          (AluOut_data_8_sva_8[0]), (AluIn_data_sva_503[256]), {and_149_cse , and_150_cse
          , and_151_cse , and_152_cse , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_286_265 <= MUX1HOT_v_22_4_2((FpAlu_8U_23U_and_35_nl), (alu_loop_op_else_else_if_mux_25_itm_4[21:0]),
          (AluOut_data_8_sva_8[22:1]), (AluIn_data_sva_503[278:257]), {nor_7_ssc
          , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_294_291 <= MUX1HOT_v_4_5_2((FpAlu_8U_23U_FpAlu_8U_23U_nor_8_nl),
          (alu_loop_op_else_else_if_mux_25_itm_4[29:26]), (AluOut_data_8_sva_8[30:27]),
          (AluIn_data_sva_503[286:283]), FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_11,
          {(and_4077_nl) , or_4809_cse , asn_1837 , or_dcpl_1087 , and_dcpl_1860});
      chn_alu_out_rsci_d_296_295 <= MUX1HOT_v_2_4_2(({{1{FpAlu_8U_23U_and_32_itm_4}},
          FpAlu_8U_23U_and_32_itm_4}), ({{1{alu_loop_op_else_else_if_mux_24_itm_4}},
          alu_loop_op_else_else_if_mux_24_itm_4}), (AluOut_data_8_sva_8[32:31]),
          (signext_2_1(AluIn_data_sva_503[287])), {nor_7_ssc , or_4809_cse , asn_1837
          , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_297 <= MUX1HOT_s_1_7_2((FpAdd_8U_23U_o_mant_10_lpi_1_dfm_2_mx0[0]),
          (FpCmp_8U_23U_true_o_22_0_10_lpi_1_dfm_6[0]), FpAlu_8U_23U_o_0_10_sva_7,
          (FpCmp_8U_23U_false_o_22_0_10_lpi_1_dfm_6[0]), alu_loop_op_else_else_if_mux_29_itm_4,
          (AluOut_data_9_sva_8[0]), (AluIn_data_sva_503[288]), {and_149_cse , and_150_cse
          , and_151_cse , and_152_cse , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_319_298 <= MUX1HOT_v_22_4_2((FpAlu_8U_23U_and_39_nl), (alu_loop_op_else_else_if_mux_28_itm_4[21:0]),
          (AluOut_data_9_sva_8[22:1]), (AluIn_data_sva_503[310:289]), {nor_7_ssc
          , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_327_324 <= MUX1HOT_v_4_5_2((FpAlu_8U_23U_FpAlu_8U_23U_nor_7_nl),
          (alu_loop_op_else_else_if_mux_28_itm_4[29:26]), (AluOut_data_9_sva_8[30:27]),
          (AluIn_data_sva_503[318:315]), FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_11,
          {(and_4071_nl) , or_4809_cse , asn_1837 , or_dcpl_1092 , and_dcpl_1868});
      chn_alu_out_rsci_d_329_328 <= MUX1HOT_v_2_4_2(({{1{FpAlu_8U_23U_and_36_itm_4}},
          FpAlu_8U_23U_and_36_itm_4}), ({{1{alu_loop_op_else_else_if_mux_27_itm_4}},
          alu_loop_op_else_else_if_mux_27_itm_4}), (AluOut_data_9_sva_8[32:31]),
          (signext_2_1(AluIn_data_sva_503[319])), {nor_7_ssc , or_4809_cse , asn_1837
          , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_330 <= MUX1HOT_s_1_7_2((FpAdd_8U_23U_o_mant_11_lpi_1_dfm_2_mx0[0]),
          (FpCmp_8U_23U_true_o_22_0_11_lpi_1_dfm_6[0]), FpAlu_8U_23U_o_0_11_sva_7,
          (FpCmp_8U_23U_false_o_22_0_11_lpi_1_dfm_6[0]), alu_loop_op_else_else_if_mux_32_itm_4,
          (AluOut_data_10_sva_8[0]), (AluIn_data_sva_503[320]), {and_149_cse , and_150_cse
          , and_151_cse , and_152_cse , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_352_331 <= MUX1HOT_v_22_4_2((FpAlu_8U_23U_and_43_nl), (alu_loop_op_else_else_if_mux_31_itm_4[21:0]),
          (AluOut_data_10_sva_8[22:1]), (AluIn_data_sva_503[342:321]), {nor_7_ssc
          , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_360_357 <= MUX1HOT_v_4_5_2((FpAlu_8U_23U_FpAlu_8U_23U_nor_6_nl),
          (alu_loop_op_else_else_if_mux_31_itm_4[29:26]), (AluOut_data_10_sva_8[30:27]),
          (AluIn_data_sva_503[350:347]), FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_11,
          {(and_4065_nl) , or_4809_cse , asn_1837 , or_dcpl_1097 , and_dcpl_1876});
      chn_alu_out_rsci_d_362_361 <= MUX1HOT_v_2_4_2(({{1{FpAlu_8U_23U_and_40_itm_4}},
          FpAlu_8U_23U_and_40_itm_4}), ({{1{alu_loop_op_else_else_if_mux_30_itm_4}},
          alu_loop_op_else_else_if_mux_30_itm_4}), (AluOut_data_10_sva_8[32:31]),
          (signext_2_1(AluIn_data_sva_503[351])), {nor_7_ssc , or_4809_cse , asn_1837
          , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_363 <= MUX1HOT_s_1_7_2((FpAdd_8U_23U_o_mant_12_lpi_1_dfm_2_mx0[0]),
          (FpCmp_8U_23U_true_o_22_0_12_lpi_1_dfm_6[0]), FpAlu_8U_23U_o_0_12_sva_7,
          (FpCmp_8U_23U_false_o_22_0_12_lpi_1_dfm_6[0]), alu_loop_op_else_else_if_mux_35_itm_4,
          (AluOut_data_11_sva_8[0]), (AluIn_data_sva_503[352]), {and_149_cse , and_150_cse
          , and_151_cse , and_152_cse , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_385_364 <= MUX1HOT_v_22_4_2((FpAlu_8U_23U_and_47_nl), (alu_loop_op_else_else_if_mux_34_itm_4[21:0]),
          (AluOut_data_11_sva_8[22:1]), (AluIn_data_sva_503[374:353]), {nor_7_ssc
          , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_393_390 <= MUX1HOT_v_4_5_2((FpAlu_8U_23U_FpAlu_8U_23U_nor_5_nl),
          (alu_loop_op_else_else_if_mux_34_itm_4[29:26]), (AluOut_data_11_sva_8[30:27]),
          (AluIn_data_sva_503[382:379]), FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_11,
          {(and_4059_nl) , or_4809_cse , asn_1837 , or_dcpl_1102 , and_dcpl_1884});
      chn_alu_out_rsci_d_395_394 <= MUX1HOT_v_2_4_2(({{1{FpAlu_8U_23U_and_44_itm_4}},
          FpAlu_8U_23U_and_44_itm_4}), ({{1{alu_loop_op_else_else_if_mux_33_itm_4}},
          alu_loop_op_else_else_if_mux_33_itm_4}), (AluOut_data_11_sva_8[32:31]),
          (signext_2_1(AluIn_data_sva_503[383])), {nor_7_ssc , or_4809_cse , asn_1837
          , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_396 <= MUX1HOT_s_1_7_2((FpAdd_8U_23U_o_mant_13_lpi_1_dfm_2_mx0[0]),
          (FpCmp_8U_23U_true_o_22_0_13_lpi_1_dfm_6[0]), FpAlu_8U_23U_o_0_13_sva_7,
          (FpCmp_8U_23U_false_o_22_0_13_lpi_1_dfm_6[0]), alu_loop_op_else_else_if_mux_38_itm_4,
          (AluOut_data_12_sva_8[0]), (AluIn_data_sva_503[384]), {and_149_cse , and_150_cse
          , and_151_cse , and_152_cse , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_418_397 <= MUX1HOT_v_22_4_2((FpAlu_8U_23U_and_51_nl), (alu_loop_op_else_else_if_mux_37_itm_4[21:0]),
          (AluOut_data_12_sva_8[22:1]), (AluIn_data_sva_503[406:385]), {nor_7_ssc
          , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_426_423 <= MUX1HOT_v_4_5_2((FpAlu_8U_23U_FpAlu_8U_23U_nor_4_nl),
          (alu_loop_op_else_else_if_mux_37_itm_4[29:26]), (AluOut_data_12_sva_8[30:27]),
          (AluIn_data_sva_503[414:411]), FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_11,
          {(and_4053_nl) , or_4809_cse , asn_1837 , or_dcpl_1107 , and_dcpl_1892});
      chn_alu_out_rsci_d_428_427 <= MUX1HOT_v_2_4_2(({{1{FpAlu_8U_23U_and_48_itm_4}},
          FpAlu_8U_23U_and_48_itm_4}), ({{1{alu_loop_op_else_else_if_mux_36_itm_4}},
          alu_loop_op_else_else_if_mux_36_itm_4}), (AluOut_data_12_sva_8[32:31]),
          (signext_2_1(AluIn_data_sva_503[415])), {nor_7_ssc , or_4809_cse , asn_1837
          , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_429 <= MUX1HOT_s_1_7_2((FpAdd_8U_23U_o_mant_14_lpi_1_dfm_2_mx0[0]),
          (FpCmp_8U_23U_true_o_22_0_14_lpi_1_dfm_6[0]), FpAlu_8U_23U_o_0_14_sva_7,
          (FpCmp_8U_23U_false_o_22_0_14_lpi_1_dfm_6[0]), alu_loop_op_else_else_if_mux_41_itm_4,
          (AluOut_data_13_sva_8[0]), (AluIn_data_sva_503[416]), {and_149_cse , and_150_cse
          , and_151_cse , and_152_cse , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_451_430 <= MUX1HOT_v_22_4_2((FpAlu_8U_23U_and_55_nl), (alu_loop_op_else_else_if_mux_40_itm_4[21:0]),
          (AluOut_data_13_sva_8[22:1]), (AluIn_data_sva_503[438:417]), {nor_7_ssc
          , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_459_456 <= MUX1HOT_v_4_5_2((FpAlu_8U_23U_FpAlu_8U_23U_nor_3_nl),
          (alu_loop_op_else_else_if_mux_40_itm_4[29:26]), (AluOut_data_13_sva_8[30:27]),
          (AluIn_data_sva_503[446:443]), FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_11,
          {(and_4047_nl) , or_4809_cse , asn_1837 , or_dcpl_1112 , and_dcpl_1900});
      chn_alu_out_rsci_d_461_460 <= MUX1HOT_v_2_4_2(({{1{FpAlu_8U_23U_and_52_itm_4}},
          FpAlu_8U_23U_and_52_itm_4}), ({{1{alu_loop_op_else_else_if_mux_39_itm_4}},
          alu_loop_op_else_else_if_mux_39_itm_4}), (AluOut_data_13_sva_8[32:31]),
          (signext_2_1(AluIn_data_sva_503[447])), {nor_7_ssc , or_4809_cse , asn_1837
          , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_462 <= MUX1HOT_s_1_7_2((FpAdd_8U_23U_o_mant_15_lpi_1_dfm_2_mx0[0]),
          (FpCmp_8U_23U_true_o_22_0_15_lpi_1_dfm_6[0]), FpAlu_8U_23U_o_0_15_sva_7,
          (FpCmp_8U_23U_false_o_22_0_15_lpi_1_dfm_6[0]), alu_loop_op_else_else_if_mux_44_itm_4,
          (AluOut_data_14_sva_8[0]), (AluIn_data_sva_503[448]), {and_149_cse , and_150_cse
          , and_151_cse , and_152_cse , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_484_463 <= MUX1HOT_v_22_4_2((FpAlu_8U_23U_and_59_nl), (alu_loop_op_else_else_if_mux_43_itm_4[21:0]),
          (AluOut_data_14_sva_8[22:1]), (AluIn_data_sva_503[470:449]), {nor_7_ssc
          , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_492_489 <= MUX1HOT_v_4_5_2((FpAlu_8U_23U_FpAlu_8U_23U_nor_2_nl),
          (alu_loop_op_else_else_if_mux_43_itm_4[29:26]), (AluOut_data_14_sva_8[30:27]),
          (AluIn_data_sva_503[478:475]), FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_11,
          {(and_4041_nl) , or_4809_cse , asn_1837 , or_dcpl_1117 , and_dcpl_1908});
      chn_alu_out_rsci_d_494_493 <= MUX1HOT_v_2_4_2(({{1{FpAlu_8U_23U_and_56_itm_4}},
          FpAlu_8U_23U_and_56_itm_4}), ({{1{alu_loop_op_else_else_if_mux_42_itm_4}},
          alu_loop_op_else_else_if_mux_42_itm_4}), (AluOut_data_14_sva_8[32:31]),
          (signext_2_1(AluIn_data_sva_503[479])), {nor_7_ssc , or_4809_cse , asn_1837
          , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_495 <= MUX1HOT_s_1_7_2((FpAdd_8U_23U_o_mant_lpi_1_dfm_2_mx0[0]),
          (FpCmp_8U_23U_true_o_22_0_lpi_1_dfm_6[0]), FpAlu_8U_23U_o_0_sva_7, (FpCmp_8U_23U_false_o_22_0_lpi_1_dfm_6[0]),
          alu_loop_op_else_else_if_mux_47_itm_4, (AluOut_data_15_sva_8[0]), (AluIn_data_sva_503[480]),
          {and_149_cse , and_150_cse , and_151_cse , and_152_cse , or_4809_cse ,
          asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_517_496 <= MUX1HOT_v_22_4_2((FpAlu_8U_23U_and_63_nl), (alu_loop_op_else_else_if_mux_46_itm_4[21:0]),
          (AluOut_data_15_sva_8[22:1]), (AluIn_data_sva_503[502:481]), {nor_7_ssc
          , or_4809_cse , asn_1837 , io_read_cfg_alu_bypass_rsc_svs_7});
      chn_alu_out_rsci_d_525_522 <= MUX1HOT_v_4_5_2((FpAlu_8U_23U_FpAlu_8U_23U_nor_1_nl),
          (alu_loop_op_else_else_if_mux_46_itm_4[29:26]), (AluOut_data_15_sva_8[30:27]),
          (AluIn_data_sva_503[510:507]), FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_11,
          {(and_4035_nl) , or_4809_cse , asn_1837 , or_dcpl_1122 , and_dcpl_1916});
      chn_alu_out_rsci_d_527_526 <= MUX1HOT_v_2_4_2(({{1{FpAlu_8U_23U_and_60_itm_4}},
          FpAlu_8U_23U_and_60_itm_4}), ({{1{alu_loop_op_else_else_if_mux_45_itm_4}},
          alu_loop_op_else_else_if_mux_45_itm_4}), (AluOut_data_15_sva_8[32:31]),
          (signext_2_1(AluIn_data_sva_503[511])), {nor_7_ssc , or_4809_cse , asn_1837
          , io_read_cfg_alu_bypass_rsc_svs_7});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_26_23 <= 4'b0;
    end
    else if ( (mux_1569_nl) & core_wen & main_stage_v_4 & or_cse_2 ) begin
      chn_alu_out_rsci_d_26_23 <= MUX1HOT_v_4_4_2((FpAlu_8U_23U_and_2_nl), (alu_loop_op_1_else_else_if_conc_itm_1_30_1_1[25:22]),
          (AluOut_data_0_sva_8[26:23]), (AluIn_data_sva_503[26:23]), {(and_4128_nl)
          , or_4809_cse , asn_1837 , or_dcpl_1047});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_59_56 <= 4'b0;
    end
    else if ( (mux_1572_nl) & core_wen & main_stage_v_4 & or_cse_2 ) begin
      chn_alu_out_rsci_d_59_56 <= MUX1HOT_v_4_4_2((FpAlu_8U_23U_and_6_nl), (alu_loop_op_2_else_else_if_conc_1_itm_1_30_1_1[25:22]),
          (AluOut_data_1_sva_8[26:23]), (AluIn_data_sva_503[58:55]), {(and_4122_nl)
          , or_4809_cse , asn_1837 , or_dcpl_1052});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_92_89 <= 4'b0;
    end
    else if ( (mux_1575_nl) & core_wen & main_stage_v_4 & or_cse_2 ) begin
      chn_alu_out_rsci_d_92_89 <= MUX1HOT_v_4_4_2((FpAlu_8U_23U_and_10_nl), (alu_loop_op_else_else_if_mux_7_itm_4[25:22]),
          (AluOut_data_2_sva_8[26:23]), (AluIn_data_sva_503[90:87]), {(and_4116_nl)
          , or_4809_cse , asn_1837 , or_dcpl_1057});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_125_122 <= 4'b0;
    end
    else if ( (mux_1578_nl) & core_wen & main_stage_v_4 & or_cse_2 ) begin
      chn_alu_out_rsci_d_125_122 <= MUX1HOT_v_4_4_2((FpAlu_8U_23U_and_14_nl), (alu_loop_op_4_else_else_if_conc_1_itm_1_30_1_1[25:22]),
          (AluOut_data_3_sva_8[26:23]), (AluIn_data_sva_503[122:119]), {(and_4110_nl)
          , or_4809_cse , asn_1837 , or_dcpl_1062});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_158_155 <= 4'b0;
    end
    else if ( (mux_1581_nl) & core_wen & main_stage_v_4 & or_cse_2 ) begin
      chn_alu_out_rsci_d_158_155 <= MUX1HOT_v_4_4_2((FpAlu_8U_23U_and_18_nl), (alu_loop_op_else_else_if_mux_13_itm_4[25:22]),
          (AluOut_data_4_sva_8[26:23]), (AluIn_data_sva_503[154:151]), {(and_4104_nl)
          , or_4809_cse , asn_1837 , or_dcpl_1067});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_191_188 <= 4'b0;
    end
    else if ( (mux_1584_nl) & core_wen & main_stage_v_4 & or_cse_2 ) begin
      chn_alu_out_rsci_d_191_188 <= MUX1HOT_v_4_4_2((FpAlu_8U_23U_and_22_nl), (alu_loop_op_else_else_if_mux_16_itm_4[25:22]),
          (AluOut_data_5_sva_8[26:23]), (AluIn_data_sva_503[186:183]), {(and_4098_nl)
          , or_4809_cse , asn_1837 , or_dcpl_1072});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_224_221 <= 4'b0;
    end
    else if ( (mux_1587_nl) & core_wen & main_stage_v_4 & or_cse_2 ) begin
      chn_alu_out_rsci_d_224_221 <= MUX1HOT_v_4_4_2((FpAlu_8U_23U_and_26_nl), (alu_loop_op_else_else_if_mux_19_itm_4[25:22]),
          (AluOut_data_6_sva_8[26:23]), (AluIn_data_sva_503[218:215]), {(and_4092_nl)
          , or_4809_cse , asn_1837 , or_dcpl_1077});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_257_254 <= 4'b0;
    end
    else if ( (mux_1590_nl) & core_wen & main_stage_v_4 & or_cse_2 ) begin
      chn_alu_out_rsci_d_257_254 <= MUX1HOT_v_4_4_2((FpAlu_8U_23U_and_30_nl), (alu_loop_op_else_else_if_mux_22_itm_4[25:22]),
          (AluOut_data_7_sva_8[26:23]), (AluIn_data_sva_503[250:247]), {(and_4086_nl)
          , or_4809_cse , asn_1837 , or_dcpl_1082});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_290_287 <= 4'b0;
    end
    else if ( (mux_1593_nl) & core_wen & main_stage_v_4 & or_cse_2 ) begin
      chn_alu_out_rsci_d_290_287 <= MUX1HOT_v_4_4_2((FpAlu_8U_23U_and_34_nl), (alu_loop_op_else_else_if_mux_25_itm_4[25:22]),
          (AluOut_data_8_sva_8[26:23]), (AluIn_data_sva_503[282:279]), {(and_4080_nl)
          , or_4809_cse , asn_1837 , or_dcpl_1087});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_323_320 <= 4'b0;
    end
    else if ( (mux_1596_nl) & core_wen & main_stage_v_4 & or_cse_2 ) begin
      chn_alu_out_rsci_d_323_320 <= MUX1HOT_v_4_4_2((FpAlu_8U_23U_and_38_nl), (alu_loop_op_else_else_if_mux_28_itm_4[25:22]),
          (AluOut_data_9_sva_8[26:23]), (AluIn_data_sva_503[314:311]), {(and_4074_nl)
          , or_4809_cse , asn_1837 , or_dcpl_1092});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_356_353 <= 4'b0;
    end
    else if ( (mux_1599_nl) & core_wen & main_stage_v_4 & or_cse_2 ) begin
      chn_alu_out_rsci_d_356_353 <= MUX1HOT_v_4_4_2((FpAlu_8U_23U_and_42_nl), (alu_loop_op_else_else_if_mux_31_itm_4[25:22]),
          (AluOut_data_10_sva_8[26:23]), (AluIn_data_sva_503[346:343]), {(and_4068_nl)
          , or_4809_cse , asn_1837 , or_dcpl_1097});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_389_386 <= 4'b0;
    end
    else if ( (mux_1602_nl) & core_wen & main_stage_v_4 & or_cse_2 ) begin
      chn_alu_out_rsci_d_389_386 <= MUX1HOT_v_4_4_2((FpAlu_8U_23U_and_46_nl), (alu_loop_op_else_else_if_mux_34_itm_4[25:22]),
          (AluOut_data_11_sva_8[26:23]), (AluIn_data_sva_503[378:375]), {(and_4062_nl)
          , or_4809_cse , asn_1837 , or_dcpl_1102});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_422_419 <= 4'b0;
    end
    else if ( (mux_1605_nl) & core_wen & main_stage_v_4 & or_cse_2 ) begin
      chn_alu_out_rsci_d_422_419 <= MUX1HOT_v_4_4_2((FpAlu_8U_23U_and_50_nl), (alu_loop_op_else_else_if_mux_37_itm_4[25:22]),
          (AluOut_data_12_sva_8[26:23]), (AluIn_data_sva_503[410:407]), {(and_4056_nl)
          , or_4809_cse , asn_1837 , or_dcpl_1107});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_455_452 <= 4'b0;
    end
    else if ( (mux_1608_nl) & core_wen & main_stage_v_4 & or_cse_2 ) begin
      chn_alu_out_rsci_d_455_452 <= MUX1HOT_v_4_4_2((FpAlu_8U_23U_and_54_nl), (alu_loop_op_else_else_if_mux_40_itm_4[25:22]),
          (AluOut_data_13_sva_8[26:23]), (AluIn_data_sva_503[442:439]), {(and_4050_nl)
          , or_4809_cse , asn_1837 , or_dcpl_1112});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_488_485 <= 4'b0;
    end
    else if ( (mux_1611_nl) & core_wen & main_stage_v_4 & or_cse_2 ) begin
      chn_alu_out_rsci_d_488_485 <= MUX1HOT_v_4_4_2((FpAlu_8U_23U_and_58_nl), (alu_loop_op_else_else_if_mux_43_itm_4[25:22]),
          (AluOut_data_14_sva_8[26:23]), (AluIn_data_sva_503[474:471]), {(and_4044_nl)
          , or_4809_cse , asn_1837 , or_dcpl_1117});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_521_518 <= 4'b0;
    end
    else if ( (mux_1614_nl) & core_wen & main_stage_v_4 & or_cse_2 ) begin
      chn_alu_out_rsci_d_521_518 <= MUX1HOT_v_4_4_2((FpAlu_8U_23U_and_62_nl), (alu_loop_op_else_else_if_mux_46_itm_4[25:22]),
          (AluOut_data_15_sva_8[26:23]), (AluIn_data_sva_503[506:503]), {(and_4038_nl)
          , or_4809_cse , asn_1837 , or_dcpl_1122});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_alu_out_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_8 | and_dcpl_10) ) begin
      reg_chn_alu_out_rsci_ld_core_psct_cse <= ~ and_dcpl_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_op_rsci_ld_core_psct <= 1'b0;
    end
    else if ( core_wen & (or_tmp_3045 | chn_alu_op_rsci_ld_core_psct_mx0c1) ) begin
      chn_alu_op_rsci_ld_core_psct <= ~ chn_alu_op_rsci_ld_core_psct_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & (or_tmp_3048 | main_stage_v_2_mx0c1) ) begin
      main_stage_v_2 <= ~ main_stage_v_2_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      AluIn_data_sva_501 <= 512'b0;
      io_read_cfg_alu_bypass_rsc_svs_st_5 <= 1'b0;
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
      alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
      alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
      alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
      alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
      alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
      alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
      alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
      alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
      alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
      alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
      alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
      alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_15_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_14_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_13_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_12_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_11_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_10_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_9_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_8_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_7_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_6_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_5_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_4_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_8 <= 1'b0;
      alu_loop_op_else_nor_tmp_80 <= 1'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp_2 <= 10'b0;
    end
    else if ( AluIn_data_and_1_cse ) begin
      AluIn_data_sva_501 <= AluIn_data_sva_1;
      io_read_cfg_alu_bypass_rsc_svs_st_5 <= io_read_cfg_alu_bypass_rsc_svs_st_1;
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
      alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
      alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
      alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
      alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
      alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
      alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
      alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
      alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
      alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
      alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
      alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
      alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1;
      IsNaN_8U_23U_land_lpi_1_dfm_8 <= IsNaN_8U_23U_land_lpi_1_dfm_4;
      IsNaN_8U_23U_land_15_lpi_1_dfm_8 <= IsNaN_8U_23U_land_15_lpi_1_dfm_4;
      IsNaN_8U_23U_land_14_lpi_1_dfm_8 <= IsNaN_8U_23U_land_14_lpi_1_dfm_4;
      IsNaN_8U_23U_land_13_lpi_1_dfm_8 <= IsNaN_8U_23U_land_13_lpi_1_dfm_4;
      IsNaN_8U_23U_land_12_lpi_1_dfm_8 <= IsNaN_8U_23U_land_12_lpi_1_dfm_4;
      IsNaN_8U_23U_land_11_lpi_1_dfm_8 <= IsNaN_8U_23U_land_11_lpi_1_dfm_4;
      IsNaN_8U_23U_land_10_lpi_1_dfm_8 <= IsNaN_8U_23U_land_10_lpi_1_dfm_4;
      IsNaN_8U_23U_land_9_lpi_1_dfm_8 <= IsNaN_8U_23U_land_9_lpi_1_dfm_4;
      IsNaN_8U_23U_land_8_lpi_1_dfm_8 <= IsNaN_8U_23U_land_8_lpi_1_dfm_4;
      IsNaN_8U_23U_land_7_lpi_1_dfm_8 <= IsNaN_8U_23U_land_7_lpi_1_dfm_4;
      IsNaN_8U_23U_land_6_lpi_1_dfm_8 <= IsNaN_8U_23U_land_6_lpi_1_dfm_4;
      IsNaN_8U_23U_land_5_lpi_1_dfm_8 <= IsNaN_8U_23U_land_5_lpi_1_dfm_4;
      IsNaN_8U_23U_land_4_lpi_1_dfm_8 <= IsNaN_8U_23U_land_4_lpi_1_dfm_4;
      IsNaN_8U_23U_land_3_lpi_1_dfm_8 <= IsNaN_8U_23U_land_3_lpi_1_dfm_4;
      IsNaN_8U_23U_land_2_lpi_1_dfm_8 <= IsNaN_8U_23U_land_2_lpi_1_dfm_4;
      IsNaN_8U_23U_land_1_lpi_1_dfm_8 <= IsNaN_8U_23U_land_1_lpi_1_dfm_4;
      alu_loop_op_else_nor_tmp_80 <= alu_loop_op_else_nor_tmp_16;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_95_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_22_13, {and_dcpl_1325
          , and_dcpl_1326 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_12_10, or_dcpl_14);
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp_2 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_94_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_9_0, {and_dcpl_1325 ,
          and_dcpl_1326 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_13_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_89_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_22_13, {and_dcpl_1274
          , and_dcpl_1275 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_12_10, or_dcpl_14);
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp_2 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_13_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_88_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_9_0, {and_dcpl_1274
          , and_dcpl_1275 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_12_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_87_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_22_13, {and_dcpl_1256
          , and_dcpl_1257 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_12_10, or_dcpl_14);
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp_2 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_12_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_86_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_9_0, {and_dcpl_1256
          , and_dcpl_1257 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_11_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_85_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_22_13, {and_dcpl_1238
          , and_dcpl_1239 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_12_10, or_dcpl_14);
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp_2 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_11_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_84_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_9_0, {and_dcpl_1238
          , and_dcpl_1239 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_10_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_83_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_22_13, {and_dcpl_1220
          , and_dcpl_1221 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_12_10, or_dcpl_14);
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp_2 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_10_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_82_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_9_0, {and_dcpl_1220
          , and_dcpl_1221 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_9_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_81_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_22_13, {and_dcpl_1206
          , and_dcpl_1207 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_12_10, or_dcpl_14);
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp_2 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_9_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_80_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_9_0, {and_dcpl_1206
          , and_dcpl_1207 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_8_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_79_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_22_13, {and_dcpl_1188
          , and_dcpl_1189 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_12_10, or_dcpl_14);
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp_2 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_8_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_78_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_9_0, {and_dcpl_1188
          , and_dcpl_1189 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_7_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_77_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_22_13, {and_dcpl_1170
          , and_dcpl_1171 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_12_10, or_dcpl_14);
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp_2 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_7_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_76_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_9_0, {and_dcpl_1170
          , and_dcpl_1171 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_6_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_75_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_22_13, {and_dcpl_1152
          , and_dcpl_1153 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_12_10, or_dcpl_14);
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp_2 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_6_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_74_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_9_0, {and_dcpl_1152
          , and_dcpl_1153 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_5_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_73_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_22_13, {and_dcpl_1134
          , and_dcpl_1135 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_12_10, or_dcpl_14);
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp_2 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_5_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_72_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_9_0, {and_dcpl_1134
          , and_dcpl_1135 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_4_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_71_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_22_13, {and_dcpl_1121
          , and_dcpl_1122 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_12_10, or_dcpl_14);
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp_2 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_4_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_70_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_9_0, {and_dcpl_1121
          , and_dcpl_1122 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_3_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_69_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_22_13, {and_dcpl_1107
          , and_dcpl_1108 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_12_10, or_dcpl_14);
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp_2 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_3_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_68_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_9_0, {and_dcpl_1107
          , and_dcpl_1108 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_2_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_67_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_22_13, {and_dcpl_1093
          , and_dcpl_1094 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_12_10, or_dcpl_14);
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp_2 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_2_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_66_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_9_0, {and_dcpl_1093
          , and_dcpl_1094 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_1_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_65_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_22_13, {and_dcpl_1079
          , and_dcpl_1080 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_12_10, or_dcpl_14);
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp_2 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_1_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_64_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_9_0, {and_dcpl_1079
          , and_dcpl_1080 , or_dcpl_14});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2 <= 1'b0;
      alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2 <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2 <= 1'b0;
      alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2 <= 1'b0;
      alu_loop_op_5_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2 <= 1'b0;
      alu_loop_op_6_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2 <= 1'b0;
      alu_loop_op_7_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2 <= 1'b0;
      alu_loop_op_8_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2 <= 1'b0;
      alu_loop_op_9_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2 <= 1'b0;
      alu_loop_op_10_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2 <= 1'b0;
      alu_loop_op_11_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2 <= 1'b0;
      alu_loop_op_12_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2 <= 1'b0;
      alu_loop_op_13_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2 <= 1'b0;
      alu_loop_op_14_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2 <= 1'b0;
      alu_loop_op_15_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2 <= 1'b0;
      alu_loop_op_16_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_is_a_greater_oelse_and_17_cse ) begin
      alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2 <= MUX_s_1_2_2(alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0,
          alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_svs, and_492_nl);
      alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2 <= MUX_s_1_2_2(alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0,
          alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs, and_509_nl);
      alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2 <= MUX_s_1_2_2(alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0,
          alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_svs, and_522_nl);
      alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2 <= MUX_s_1_2_2(alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0,
          alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs, and_535_nl);
      alu_loop_op_5_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2 <= MUX_s_1_2_2(alu_loop_op_5_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0,
          alu_loop_op_5_FpAdd_8U_23U_is_a_greater_oif_equal_svs, and_548_nl);
      alu_loop_op_6_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2 <= MUX_s_1_2_2(alu_loop_op_6_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0,
          alu_loop_op_6_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs, and_561_nl);
      alu_loop_op_7_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2 <= MUX_s_1_2_2(alu_loop_op_7_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0,
          alu_loop_op_7_FpAdd_8U_23U_is_a_greater_oif_equal_svs, and_574_nl);
      alu_loop_op_8_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2 <= MUX_s_1_2_2(alu_loop_op_8_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0,
          alu_loop_op_8_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs, and_587_nl);
      alu_loop_op_9_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2 <= MUX_s_1_2_2(alu_loop_op_9_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0,
          alu_loop_op_9_FpAdd_8U_23U_is_a_greater_oif_equal_svs, and_600_nl);
      alu_loop_op_10_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2 <= MUX_s_1_2_2(alu_loop_op_10_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0,
          alu_loop_op_10_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs, and_613_nl);
      alu_loop_op_11_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2 <= MUX_s_1_2_2(alu_loop_op_11_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0,
          alu_loop_op_11_FpAdd_8U_23U_is_a_greater_oif_equal_svs, and_626_nl);
      alu_loop_op_12_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2 <= MUX_s_1_2_2(alu_loop_op_12_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0,
          alu_loop_op_12_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs, and_639_nl);
      alu_loop_op_13_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2 <= MUX_s_1_2_2(alu_loop_op_13_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0,
          alu_loop_op_13_FpAdd_8U_23U_is_a_greater_oif_equal_svs, and_652_nl);
      alu_loop_op_14_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2 <= MUX_s_1_2_2(alu_loop_op_14_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0,
          alu_loop_op_14_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs, and_665_nl);
      alu_loop_op_15_FpAdd_8U_23U_is_a_greater_oif_equal_svs_2 <= MUX_s_1_2_2(alu_loop_op_15_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0,
          alu_loop_op_15_FpAdd_8U_23U_is_a_greater_oif_equal_svs, and_678_nl);
      alu_loop_op_16_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_2 <= MUX_s_1_2_2(alu_loop_op_16_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0,
          alu_loop_op_16_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs, and_691_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_9 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3, and_dcpl_30);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3, and_dcpl_30);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_st_2 <= 1'b0;
      alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_st_2 <= 1'b0;
      alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_st_2 <= 1'b0;
      alu_loop_op_4_FpCmp_8U_23U_false_slc_8_1_svs_st_2 <= 1'b0;
      alu_loop_op_5_FpCmp_8U_23U_false_slc_8_svs_st_2 <= 1'b0;
      alu_loop_op_6_FpCmp_8U_23U_false_slc_8_1_svs_st_2 <= 1'b0;
      alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_st_2 <= 1'b0;
      alu_loop_op_9_FpCmp_8U_23U_false_slc_8_svs_st_2 <= 1'b0;
      alu_loop_op_10_FpCmp_8U_23U_false_slc_8_1_svs_st_2 <= 1'b0;
      alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_st_2 <= 1'b0;
      alu_loop_op_13_FpCmp_8U_23U_false_slc_8_svs_st_2 <= 1'b0;
      alu_loop_op_14_FpCmp_8U_23U_false_slc_8_1_svs_st_2 <= 1'b0;
      alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_st_2 <= 1'b0;
      alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_st_2 <= 1'b0;
    end
    else if ( FpCmp_8U_23U_false_if_and_32_cse ) begin
      alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_st_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_16_itm_8_1,
          alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_st, alu_loop_op_1_FpCmp_8U_23U_true_slc_8_svs_st,
          IsNaN_8U_23U_2_land_1_lpi_1_dfm_st_1, {and_498_rgt , and_dcpl_34 , and_dcpl_36
          , and_543_rgt});
      alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_st_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_18_itm_8_1,
          alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_st, alu_loop_op_2_FpCmp_8U_23U_true_slc_8_1_svs_st,
          IsNaN_8U_23U_2_land_2_lpi_1_dfm_st_1, {and_498_rgt , and_dcpl_34 , and_dcpl_36
          , and_543_rgt});
      alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_st_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_20_itm_8_1,
          alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_st, alu_loop_op_3_FpCmp_8U_23U_true_slc_8_svs_st,
          IsNaN_8U_23U_2_land_3_lpi_1_dfm_st_1, {and_498_rgt , and_dcpl_34 , and_dcpl_36
          , and_543_rgt});
      alu_loop_op_4_FpCmp_8U_23U_false_slc_8_1_svs_st_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_22_itm_8_1,
          alu_loop_op_4_FpCmp_8U_23U_false_slc_8_1_svs_st, alu_loop_op_4_FpCmp_8U_23U_true_slc_8_1_svs_st,
          IsNaN_8U_23U_2_land_4_lpi_1_dfm_st_1, {and_498_rgt , and_dcpl_34 , and_dcpl_36
          , and_543_rgt});
      alu_loop_op_5_FpCmp_8U_23U_false_slc_8_svs_st_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_24_itm_8_1,
          alu_loop_op_5_FpCmp_8U_23U_false_slc_8_svs_st, alu_loop_op_5_FpCmp_8U_23U_true_slc_8_svs_st,
          IsNaN_8U_23U_2_land_5_lpi_1_dfm_st_1, {and_498_rgt , and_dcpl_34 , and_dcpl_36
          , and_543_rgt});
      alu_loop_op_6_FpCmp_8U_23U_false_slc_8_1_svs_st_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_26_itm_8_1,
          alu_loop_op_6_FpCmp_8U_23U_false_slc_8_1_svs_st, alu_loop_op_6_FpCmp_8U_23U_true_slc_8_1_svs_st,
          IsNaN_8U_23U_2_land_6_lpi_1_dfm_st_1, {and_498_rgt , and_dcpl_34 , and_dcpl_36
          , and_543_rgt});
      alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_st_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_28_itm_8_1,
          alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_st, alu_loop_op_7_FpCmp_8U_23U_true_slc_8_svs_st,
          IsNaN_8U_23U_2_land_7_lpi_1_dfm_st_1, {and_498_rgt , and_dcpl_34 , and_dcpl_36
          , and_543_rgt});
      alu_loop_op_9_FpCmp_8U_23U_false_slc_8_svs_st_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_32_itm_8_1,
          alu_loop_op_9_FpCmp_8U_23U_false_slc_8_svs_st, alu_loop_op_9_FpCmp_8U_23U_true_slc_8_svs_st,
          IsNaN_8U_23U_2_land_9_lpi_1_dfm_st_1, {and_498_rgt , and_dcpl_34 , and_dcpl_36
          , and_543_rgt});
      alu_loop_op_10_FpCmp_8U_23U_false_slc_8_1_svs_st_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_34_itm_8_1,
          alu_loop_op_10_FpCmp_8U_23U_false_slc_8_1_svs_st, alu_loop_op_10_FpCmp_8U_23U_true_slc_8_1_svs_st,
          IsNaN_8U_23U_2_land_10_lpi_1_dfm_st_1, {and_498_rgt , and_dcpl_34 , and_dcpl_36
          , and_543_rgt});
      alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_st_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_36_itm_8_1,
          alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_st, alu_loop_op_11_FpCmp_8U_23U_true_slc_8_svs_st,
          IsNaN_8U_23U_2_land_11_lpi_1_dfm_st_1, {and_498_rgt , and_dcpl_34 , and_dcpl_36
          , and_543_rgt});
      alu_loop_op_13_FpCmp_8U_23U_false_slc_8_svs_st_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_40_itm_8_1,
          alu_loop_op_13_FpCmp_8U_23U_false_slc_8_svs_st, alu_loop_op_13_FpCmp_8U_23U_true_slc_8_svs_st,
          IsNaN_8U_23U_2_land_13_lpi_1_dfm_st_1, {and_498_rgt , and_dcpl_34 , and_dcpl_36
          , and_543_rgt});
      alu_loop_op_14_FpCmp_8U_23U_false_slc_8_1_svs_st_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_42_itm_8_1,
          alu_loop_op_14_FpCmp_8U_23U_false_slc_8_1_svs_st, alu_loop_op_14_FpCmp_8U_23U_true_slc_8_1_svs_st,
          IsNaN_8U_23U_2_land_14_lpi_1_dfm_st_1, {and_498_rgt , and_dcpl_34 , and_dcpl_36
          , and_543_rgt});
      alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_st_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_44_itm_8_1,
          alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_st, alu_loop_op_15_FpCmp_8U_23U_true_slc_8_svs_st,
          IsNaN_8U_23U_2_land_15_lpi_1_dfm_st_1, {and_498_rgt , and_dcpl_34 , and_dcpl_36
          , and_543_rgt});
      alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_st_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_46_itm_8_1,
          alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_st, alu_loop_op_16_FpCmp_8U_23U_true_slc_8_1_svs_st,
          IsNaN_8U_23U_2_land_lpi_1_dfm_st_1, {and_498_rgt , and_dcpl_34 , and_dcpl_36
          , and_543_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_is_a_greater_oelse_FpAdd_8U_23U_is_a_greater_oelse_or_21_cse
        & (mux_18_nl) ) begin
      alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_st_2 <= MUX_s_1_2_2(alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0,
          alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_st, and_dcpl_23);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_2_FpAdd_8U_23U_is_a_greater_slc_8_1_svs_st_2 <= 1'b0;
      alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3
          <= 1'b0;
      alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3
          <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3
          <= 1'b0;
      alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3
          <= 1'b0;
      alu_loop_op_5_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3
          <= 1'b0;
      alu_loop_op_6_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3
          <= 1'b0;
      alu_loop_op_7_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3
          <= 1'b0;
      alu_loop_op_8_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3
          <= 1'b0;
      alu_loop_op_9_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3
          <= 1'b0;
      alu_loop_op_10_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3
          <= 1'b0;
      alu_loop_op_11_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3
          <= 1'b0;
      alu_loop_op_12_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3
          <= 1'b0;
      alu_loop_op_13_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3
          <= 1'b0;
      alu_loop_op_14_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3
          <= 1'b0;
      alu_loop_op_15_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3
          <= 1'b0;
      alu_loop_op_16_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3
          <= 1'b0;
      alu_loop_op_4_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm_2 <= 1'b0;
      alu_loop_op_4_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm_2 <= 1'b0;
      alu_loop_op_6_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm_2 <= 1'b0;
      alu_loop_op_6_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm_2 <= 1'b0;
      alu_loop_op_13_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_itm_2 <= 1'b0;
      alu_loop_op_13_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_itm_2 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_is_a_greater_and_17_cse ) begin
      alu_loop_op_2_FpAdd_8U_23U_is_a_greater_slc_8_1_svs_st_2 <= MUX_s_1_2_2(FpCmp_8U_23U_true_if_acc_18_itm_8_1,
          reg_alu_loop_op_2_FpAdd_8U_23U_is_a_greater_slc_8_1_svs_cse, and_dcpl_23);
      alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3
          <= MUX_s_1_2_2(alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0,
          alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st,
          and_dcpl_23);
      alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3
          <= MUX_s_1_2_2(alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0,
          alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st,
          and_dcpl_23);
      alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3
          <= MUX_s_1_2_2(alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0,
          alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st,
          and_dcpl_23);
      alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3
          <= MUX_s_1_2_2(alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0,
          alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st,
          and_dcpl_23);
      alu_loop_op_5_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3
          <= MUX_s_1_2_2(alu_loop_op_5_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0,
          alu_loop_op_5_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st,
          and_dcpl_23);
      alu_loop_op_6_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3
          <= MUX_s_1_2_2(alu_loop_op_6_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0,
          alu_loop_op_6_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st,
          and_dcpl_23);
      alu_loop_op_7_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3
          <= MUX_s_1_2_2(alu_loop_op_7_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0,
          alu_loop_op_7_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st,
          and_dcpl_23);
      alu_loop_op_8_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3
          <= MUX_s_1_2_2(alu_loop_op_8_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0,
          alu_loop_op_8_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st,
          and_dcpl_23);
      alu_loop_op_9_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3
          <= MUX_s_1_2_2(alu_loop_op_9_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0,
          alu_loop_op_9_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st,
          and_dcpl_23);
      alu_loop_op_10_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3
          <= MUX_s_1_2_2(alu_loop_op_10_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0,
          alu_loop_op_10_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st,
          and_dcpl_23);
      alu_loop_op_11_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3
          <= MUX_s_1_2_2(alu_loop_op_11_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0,
          alu_loop_op_11_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st,
          and_dcpl_23);
      alu_loop_op_12_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3
          <= MUX_s_1_2_2(alu_loop_op_12_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0,
          alu_loop_op_12_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st,
          and_dcpl_23);
      alu_loop_op_13_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3
          <= MUX_s_1_2_2(alu_loop_op_13_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0,
          alu_loop_op_13_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st,
          and_dcpl_23);
      alu_loop_op_14_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3
          <= MUX_s_1_2_2(alu_loop_op_14_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0,
          alu_loop_op_14_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st,
          and_dcpl_23);
      alu_loop_op_15_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3
          <= MUX_s_1_2_2(alu_loop_op_15_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0,
          alu_loop_op_15_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st,
          and_dcpl_23);
      alu_loop_op_16_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3
          <= MUX_s_1_2_2(alu_loop_op_16_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0,
          alu_loop_op_16_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st,
          and_dcpl_23);
      alu_loop_op_4_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm_2 <= MUX_s_1_2_2(alu_loop_op_4_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm_mx0w0,
          alu_loop_op_4_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm, and_dcpl_23);
      alu_loop_op_4_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm_2 <= MUX_s_1_2_2(alu_loop_op_4_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm_mx0w0,
          alu_loop_op_4_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm, and_dcpl_23);
      alu_loop_op_6_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm_2 <= MUX_s_1_2_2(alu_loop_op_6_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm_mx0w0,
          alu_loop_op_6_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm, and_dcpl_23);
      alu_loop_op_6_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm_2 <= MUX_s_1_2_2(alu_loop_op_6_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm_mx0w0,
          alu_loop_op_6_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm, and_dcpl_23);
      alu_loop_op_13_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_itm_2 <= MUX_s_1_2_2(alu_loop_op_13_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_itm_mx0w0,
          alu_loop_op_13_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_itm, and_dcpl_23);
      alu_loop_op_13_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_itm_2 <= MUX_s_1_2_2(alu_loop_op_13_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_itm_mx0w0,
          alu_loop_op_13_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_itm, and_dcpl_23);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_st_2 <= 1'b0;
      alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_st_2 <= 1'b0;
    end
    else if ( FpCmp_8U_23U_false_if_and_39_cse ) begin
      alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_st_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_30_itm_8_1,
          alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_st, alu_loop_op_8_FpCmp_8U_23U_true_slc_8_1_svs_st,
          IsNaN_8U_23U_2_land_8_lpi_1_dfm_st_1, {and_589_rgt , and_dcpl_34 , and_dcpl_127
          , and_543_rgt});
      alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_st_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_38_itm_8_1,
          alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_st, alu_loop_op_12_FpCmp_8U_23U_true_slc_8_1_svs_st,
          IsNaN_8U_23U_2_land_12_lpi_1_dfm_st_1, {and_589_rgt , and_dcpl_34 , and_dcpl_127
          , and_543_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_cfg_alu_algo_1_sva_st_93_cse <= 2'b0;
      reg_cfg_alu_algo_1_sva_st_157_cse <= 2'b0;
      IsNaN_8U_23U_3_land_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_4_land_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_3_land_15_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_4_land_15_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_3_land_14_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_4_land_14_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_3_land_13_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_4_land_13_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_3_land_12_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_4_land_12_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_3_land_11_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_4_land_11_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_3_land_10_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_4_land_10_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_3_land_9_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_4_land_9_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_3_land_8_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_4_land_8_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_3_land_7_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_4_land_7_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_3_land_6_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_4_land_6_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_3_land_5_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_4_land_5_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_3_land_4_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_4_land_4_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_3_land_3_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_4_land_3_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_3_land_2_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_4_land_2_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_3_land_1_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_4_land_1_lpi_1_dfm_6 <= 1'b0;
      cfg_alu_algo_1_sva_5 <= 2'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp_2 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_75_cse ) begin
      reg_cfg_alu_algo_1_sva_st_93_cse <= cfg_alu_algo_1_sva_st_92;
      reg_cfg_alu_algo_1_sva_st_157_cse <= cfg_alu_algo_1_sva_st_96;
      IsNaN_8U_23U_3_land_lpi_1_dfm_6 <= IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_4_land_lpi_1_dfm_6 <= IsNaN_8U_23U_4_land_lpi_1_dfm_4;
      IsNaN_8U_23U_3_land_15_lpi_1_dfm_6 <= IsNaN_8U_23U_3_land_15_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_4_land_15_lpi_1_dfm_6 <= IsNaN_8U_23U_4_land_15_lpi_1_dfm_4;
      IsNaN_8U_23U_3_land_14_lpi_1_dfm_6 <= IsNaN_8U_23U_3_land_14_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_4_land_14_lpi_1_dfm_6 <= IsNaN_8U_23U_4_land_14_lpi_1_dfm_4;
      IsNaN_8U_23U_3_land_13_lpi_1_dfm_6 <= IsNaN_8U_23U_3_land_13_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_4_land_13_lpi_1_dfm_6 <= IsNaN_8U_23U_4_land_13_lpi_1_dfm_4;
      IsNaN_8U_23U_3_land_12_lpi_1_dfm_6 <= IsNaN_8U_23U_3_land_12_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_4_land_12_lpi_1_dfm_6 <= IsNaN_8U_23U_4_land_12_lpi_1_dfm_4;
      IsNaN_8U_23U_3_land_11_lpi_1_dfm_6 <= IsNaN_8U_23U_3_land_11_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_4_land_11_lpi_1_dfm_6 <= IsNaN_8U_23U_4_land_11_lpi_1_dfm_4;
      IsNaN_8U_23U_3_land_10_lpi_1_dfm_6 <= IsNaN_8U_23U_3_land_10_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_4_land_10_lpi_1_dfm_6 <= IsNaN_8U_23U_4_land_10_lpi_1_dfm_4;
      IsNaN_8U_23U_3_land_9_lpi_1_dfm_6 <= IsNaN_8U_23U_3_land_9_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_4_land_9_lpi_1_dfm_6 <= IsNaN_8U_23U_4_land_9_lpi_1_dfm_4;
      IsNaN_8U_23U_3_land_8_lpi_1_dfm_6 <= IsNaN_8U_23U_3_land_8_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_4_land_8_lpi_1_dfm_6 <= IsNaN_8U_23U_4_land_8_lpi_1_dfm_4;
      IsNaN_8U_23U_3_land_7_lpi_1_dfm_6 <= IsNaN_8U_23U_3_land_7_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_4_land_7_lpi_1_dfm_6 <= IsNaN_8U_23U_4_land_7_lpi_1_dfm_4;
      IsNaN_8U_23U_3_land_6_lpi_1_dfm_6 <= IsNaN_8U_23U_3_land_6_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_4_land_6_lpi_1_dfm_6 <= IsNaN_8U_23U_4_land_6_lpi_1_dfm_4;
      IsNaN_8U_23U_3_land_5_lpi_1_dfm_6 <= IsNaN_8U_23U_3_land_5_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_4_land_5_lpi_1_dfm_6 <= IsNaN_8U_23U_4_land_5_lpi_1_dfm_4;
      IsNaN_8U_23U_3_land_4_lpi_1_dfm_6 <= IsNaN_8U_23U_3_land_4_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_4_land_4_lpi_1_dfm_6 <= IsNaN_8U_23U_4_land_4_lpi_1_dfm_4;
      IsNaN_8U_23U_3_land_3_lpi_1_dfm_6 <= IsNaN_8U_23U_3_land_3_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_4_land_3_lpi_1_dfm_6 <= IsNaN_8U_23U_4_land_3_lpi_1_dfm_4;
      IsNaN_8U_23U_3_land_2_lpi_1_dfm_6 <= IsNaN_8U_23U_3_land_2_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_4_land_2_lpi_1_dfm_6 <= IsNaN_8U_23U_4_land_2_lpi_1_dfm_4;
      IsNaN_8U_23U_3_land_1_lpi_1_dfm_6 <= IsNaN_8U_23U_3_land_1_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_4_land_1_lpi_1_dfm_6 <= IsNaN_8U_23U_4_land_1_lpi_1_dfm_4;
      cfg_alu_algo_1_sva_5 <= cfg_alu_algo_1_sva_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_15_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_93_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_22_13, {and_dcpl_1307
          , and_dcpl_1308 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_12_10, or_dcpl_14);
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp_2 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_15_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_92_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_9_0, {and_dcpl_1307
          , and_dcpl_1308 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_14_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_91_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_22_13, {and_dcpl_1289
          , and_dcpl_1290 , or_dcpl_14});
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_12_10, or_dcpl_14);
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp_2 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_14_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_90_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_9_0, {and_dcpl_1289
          , and_dcpl_1290 , or_dcpl_14});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_3 <= 1'b0;
    end
    else if ( core_wen & ((or_cse_2 & main_stage_v_2) | main_stage_v_3_mx0c1) ) begin
      main_stage_v_3 <= ~ main_stage_v_3_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
          <= 1'b0;
      reg_alu_loop_op_6_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
          <= 1'b0;
      reg_alu_loop_op_7_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
          <= 1'b0;
      reg_alu_loop_op_8_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
          <= 1'b0;
      reg_alu_loop_op_9_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
          <= 1'b0;
      reg_alu_loop_op_10_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
          <= 1'b0;
      reg_alu_loop_op_13_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
          <= 1'b0;
      reg_alu_loop_op_14_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
          <= 1'b0;
      reg_alu_loop_op_15_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
          <= 1'b0;
      reg_alu_loop_op_16_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
          <= 1'b0;
    end
    else if ( FpAdd_8U_23U_is_addition_and_cse ) begin
      reg_alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
          <= alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
      reg_alu_loop_op_6_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
          <= alu_loop_op_6_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3;
      reg_alu_loop_op_7_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
          <= alu_loop_op_7_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
      reg_alu_loop_op_8_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
          <= alu_loop_op_8_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3;
      reg_alu_loop_op_9_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
          <= alu_loop_op_9_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
      reg_alu_loop_op_10_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
          <= alu_loop_op_10_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3;
      reg_alu_loop_op_13_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
          <= alu_loop_op_13_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
      reg_alu_loop_op_14_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
          <= alu_loop_op_14_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3;
      reg_alu_loop_op_15_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
          <= alu_loop_op_15_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
      reg_alu_loop_op_16_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
          <= alu_loop_op_16_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4 <= 1'b0;
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= 1'b0;
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4 <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= 1'b0;
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= 1'b0;
      alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= 1'b0;
      alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= 1'b0;
      alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4 <= 1'b0;
      alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= 1'b0;
      alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4 <= 1'b0;
      alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= 1'b0;
      alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= 1'b0;
      alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= 1'b0;
      alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= 1'b0;
      alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= 1'b0;
      alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= 1'b0;
      alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= 1'b0;
      alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4 <= 1'b0;
      alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= 1'b0;
      alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4 <= 1'b0;
      alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= 1'b0;
    end
    else if ( IsZero_8U_23U_1_and_cse ) begin
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4 <= alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3;
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4 <= alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3;
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
      alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
      alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
      alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4 <= alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3;
      alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
      alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4 <= alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3;
      alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
      alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
      alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
      alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
      alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
      alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
      alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
      alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4 <= alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3;
      alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
      alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_4 <= alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3;
      alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_itm_2 <= 8'b0;
      alu_loop_op_1_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2
          <= 1'b0;
      alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_itm_2 <= 8'b0;
      alu_loop_op_1_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2
          <= 1'b0;
      alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_1_itm_2 <= 8'b0;
      alu_loop_op_2_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2
          <= 1'b0;
      alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_1_itm_2 <= 8'b0;
      alu_loop_op_2_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2
          <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_itm_2 <= 8'b0;
      alu_loop_op_3_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2
          <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_itm_2 <= 8'b0;
      alu_loop_op_3_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2
          <= 1'b0;
      alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_1_itm_2 <= 8'b0;
      alu_loop_op_4_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2
          <= 1'b0;
      alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_1_itm_2 <= 8'b0;
      alu_loop_op_4_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2
          <= 1'b0;
      alu_loop_op_5_FpAdd_8U_23U_b_left_shift_acc_itm_2 <= 8'b0;
      alu_loop_op_5_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2
          <= 1'b0;
      alu_loop_op_5_FpAdd_8U_23U_a_left_shift_acc_itm_2 <= 8'b0;
      alu_loop_op_5_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2
          <= 1'b0;
      alu_loop_op_6_FpAdd_8U_23U_b_left_shift_acc_1_itm_2 <= 8'b0;
      alu_loop_op_6_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2
          <= 1'b0;
      alu_loop_op_6_FpAdd_8U_23U_a_left_shift_acc_1_itm_2 <= 8'b0;
      alu_loop_op_6_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2
          <= 1'b0;
      alu_loop_op_7_FpAdd_8U_23U_b_left_shift_acc_itm_2 <= 8'b0;
      alu_loop_op_7_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2
          <= 1'b0;
      alu_loop_op_7_FpAdd_8U_23U_a_left_shift_acc_itm_2 <= 8'b0;
      alu_loop_op_7_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2
          <= 1'b0;
      alu_loop_op_8_FpAdd_8U_23U_b_left_shift_acc_1_itm_2 <= 8'b0;
      alu_loop_op_8_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2
          <= 1'b0;
      alu_loop_op_8_FpAdd_8U_23U_a_left_shift_acc_1_itm_2 <= 8'b0;
      alu_loop_op_8_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2
          <= 1'b0;
      alu_loop_op_9_FpAdd_8U_23U_b_left_shift_acc_itm_2 <= 8'b0;
      alu_loop_op_9_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2
          <= 1'b0;
      alu_loop_op_9_FpAdd_8U_23U_a_left_shift_acc_itm_2 <= 8'b0;
      alu_loop_op_9_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2
          <= 1'b0;
      alu_loop_op_10_FpAdd_8U_23U_b_left_shift_acc_1_itm_2 <= 8'b0;
      alu_loop_op_10_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2
          <= 1'b0;
      alu_loop_op_10_FpAdd_8U_23U_a_left_shift_acc_1_itm_2 <= 8'b0;
      alu_loop_op_10_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2
          <= 1'b0;
      alu_loop_op_11_FpAdd_8U_23U_b_left_shift_acc_itm_2 <= 8'b0;
      alu_loop_op_11_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2
          <= 1'b0;
      alu_loop_op_11_FpAdd_8U_23U_a_left_shift_acc_itm_2 <= 8'b0;
      alu_loop_op_11_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2
          <= 1'b0;
      alu_loop_op_12_FpAdd_8U_23U_b_left_shift_acc_1_itm_2 <= 8'b0;
      alu_loop_op_12_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2
          <= 1'b0;
      alu_loop_op_12_FpAdd_8U_23U_a_left_shift_acc_1_itm_2 <= 8'b0;
      alu_loop_op_12_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2
          <= 1'b0;
      alu_loop_op_13_FpAdd_8U_23U_b_left_shift_acc_itm_2 <= 8'b0;
      alu_loop_op_13_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2
          <= 1'b0;
      alu_loop_op_13_FpAdd_8U_23U_a_left_shift_acc_itm_2 <= 8'b0;
      alu_loop_op_13_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2
          <= 1'b0;
      alu_loop_op_14_FpAdd_8U_23U_b_left_shift_acc_1_itm_2 <= 8'b0;
      alu_loop_op_14_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2
          <= 1'b0;
      alu_loop_op_14_FpAdd_8U_23U_a_left_shift_acc_1_itm_2 <= 8'b0;
      alu_loop_op_14_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2
          <= 1'b0;
      alu_loop_op_15_FpAdd_8U_23U_b_left_shift_acc_itm_2 <= 8'b0;
      alu_loop_op_15_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2
          <= 1'b0;
      alu_loop_op_15_FpAdd_8U_23U_a_left_shift_acc_itm_2 <= 8'b0;
      alu_loop_op_15_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2
          <= 1'b0;
      alu_loop_op_16_FpAdd_8U_23U_b_left_shift_acc_1_itm_2 <= 8'b0;
      alu_loop_op_16_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2
          <= 1'b0;
      alu_loop_op_16_FpAdd_8U_23U_a_left_shift_acc_1_itm_2 <= 8'b0;
      alu_loop_op_16_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2
          <= 1'b0;
    end
    else if ( FpAdd_8U_23U_b_left_shift_and_32_cse ) begin
      alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_itm_2 <= MUX_v_8_2_2(alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0,
          alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_itm, and_dcpl_241);
      alu_loop_op_1_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm[0]), alu_loop_op_1_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm,
          and_dcpl_241);
      alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_itm_2 <= MUX_v_8_2_2(alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0,
          alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_itm, and_dcpl_241);
      alu_loop_op_1_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm[0]), alu_loop_op_1_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm,
          and_dcpl_241);
      alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_1_itm_2 <= MUX_v_8_2_2(alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0,
          alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_1_itm, and_dcpl_241);
      alu_loop_op_2_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm[0]), alu_loop_op_2_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm,
          and_dcpl_241);
      alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_1_itm_2 <= MUX_v_8_2_2(alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0,
          alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_1_itm, and_dcpl_241);
      alu_loop_op_2_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm[0]), alu_loop_op_2_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm,
          and_dcpl_241);
      alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_itm_2 <= MUX_v_8_2_2(alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0,
          alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_itm, and_dcpl_241);
      alu_loop_op_3_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm[0]), alu_loop_op_3_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm,
          and_dcpl_241);
      alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_itm_2 <= MUX_v_8_2_2(alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0,
          alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_itm, and_dcpl_241);
      alu_loop_op_3_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm[0]), alu_loop_op_3_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm,
          and_dcpl_241);
      alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_1_itm_2 <= MUX_v_8_2_2(alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0,
          alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_1_itm, and_dcpl_241);
      alu_loop_op_4_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_b_right_shift_qr_4_lpi_1_dfm[0]), alu_loop_op_4_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm,
          and_dcpl_241);
      alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_1_itm_2 <= MUX_v_8_2_2(alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0,
          alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_1_itm, and_dcpl_241);
      alu_loop_op_4_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_a_right_shift_qr_4_lpi_1_dfm[0]), alu_loop_op_4_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm,
          and_dcpl_241);
      alu_loop_op_5_FpAdd_8U_23U_b_left_shift_acc_itm_2 <= MUX_v_8_2_2(alu_loop_op_5_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0,
          alu_loop_op_5_FpAdd_8U_23U_b_left_shift_acc_itm, and_dcpl_241);
      alu_loop_op_5_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_b_right_shift_qr_5_lpi_1_dfm[0]), alu_loop_op_5_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm,
          and_dcpl_241);
      alu_loop_op_5_FpAdd_8U_23U_a_left_shift_acc_itm_2 <= MUX_v_8_2_2(alu_loop_op_5_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0,
          alu_loop_op_5_FpAdd_8U_23U_a_left_shift_acc_itm, and_dcpl_241);
      alu_loop_op_5_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_a_right_shift_qr_5_lpi_1_dfm[0]), alu_loop_op_5_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm,
          and_dcpl_241);
      alu_loop_op_6_FpAdd_8U_23U_b_left_shift_acc_1_itm_2 <= MUX_v_8_2_2(alu_loop_op_6_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0,
          alu_loop_op_6_FpAdd_8U_23U_b_left_shift_acc_1_itm, and_dcpl_241);
      alu_loop_op_6_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_b_right_shift_qr_6_lpi_1_dfm[0]), alu_loop_op_6_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm,
          and_dcpl_241);
      alu_loop_op_6_FpAdd_8U_23U_a_left_shift_acc_1_itm_2 <= MUX_v_8_2_2(alu_loop_op_6_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0,
          alu_loop_op_6_FpAdd_8U_23U_a_left_shift_acc_1_itm, and_dcpl_241);
      alu_loop_op_6_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_a_right_shift_qr_6_lpi_1_dfm[0]), alu_loop_op_6_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm,
          and_dcpl_241);
      alu_loop_op_7_FpAdd_8U_23U_b_left_shift_acc_itm_2 <= MUX_v_8_2_2(alu_loop_op_7_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0,
          alu_loop_op_7_FpAdd_8U_23U_b_left_shift_acc_itm, and_dcpl_241);
      alu_loop_op_7_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_b_right_shift_qr_7_lpi_1_dfm[0]), alu_loop_op_7_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm,
          and_dcpl_241);
      alu_loop_op_7_FpAdd_8U_23U_a_left_shift_acc_itm_2 <= MUX_v_8_2_2(alu_loop_op_7_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0,
          alu_loop_op_7_FpAdd_8U_23U_a_left_shift_acc_itm, and_dcpl_241);
      alu_loop_op_7_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_a_right_shift_qr_7_lpi_1_dfm[0]), alu_loop_op_7_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm,
          and_dcpl_241);
      alu_loop_op_8_FpAdd_8U_23U_b_left_shift_acc_1_itm_2 <= MUX_v_8_2_2(alu_loop_op_8_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0,
          alu_loop_op_8_FpAdd_8U_23U_b_left_shift_acc_1_itm, and_dcpl_241);
      alu_loop_op_8_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_b_right_shift_qr_8_lpi_1_dfm[0]), alu_loop_op_8_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm,
          and_dcpl_241);
      alu_loop_op_8_FpAdd_8U_23U_a_left_shift_acc_1_itm_2 <= MUX_v_8_2_2(alu_loop_op_8_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0,
          alu_loop_op_8_FpAdd_8U_23U_a_left_shift_acc_1_itm, and_dcpl_241);
      alu_loop_op_8_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_a_right_shift_qr_8_lpi_1_dfm[0]), alu_loop_op_8_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm,
          and_dcpl_241);
      alu_loop_op_9_FpAdd_8U_23U_b_left_shift_acc_itm_2 <= MUX_v_8_2_2(alu_loop_op_9_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0,
          alu_loop_op_9_FpAdd_8U_23U_b_left_shift_acc_itm, and_dcpl_241);
      alu_loop_op_9_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_b_right_shift_qr_9_lpi_1_dfm[0]), alu_loop_op_9_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm,
          and_dcpl_241);
      alu_loop_op_9_FpAdd_8U_23U_a_left_shift_acc_itm_2 <= MUX_v_8_2_2(alu_loop_op_9_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0,
          alu_loop_op_9_FpAdd_8U_23U_a_left_shift_acc_itm, and_dcpl_241);
      alu_loop_op_9_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_a_right_shift_qr_9_lpi_1_dfm[0]), alu_loop_op_9_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm,
          and_dcpl_241);
      alu_loop_op_10_FpAdd_8U_23U_b_left_shift_acc_1_itm_2 <= MUX_v_8_2_2(alu_loop_op_10_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0,
          alu_loop_op_10_FpAdd_8U_23U_b_left_shift_acc_1_itm, and_dcpl_241);
      alu_loop_op_10_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_b_right_shift_qr_10_lpi_1_dfm[0]), alu_loop_op_10_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm,
          and_dcpl_241);
      alu_loop_op_10_FpAdd_8U_23U_a_left_shift_acc_1_itm_2 <= MUX_v_8_2_2(alu_loop_op_10_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0,
          alu_loop_op_10_FpAdd_8U_23U_a_left_shift_acc_1_itm, and_dcpl_241);
      alu_loop_op_10_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_a_right_shift_qr_10_lpi_1_dfm[0]), alu_loop_op_10_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm,
          and_dcpl_241);
      alu_loop_op_11_FpAdd_8U_23U_b_left_shift_acc_itm_2 <= MUX_v_8_2_2(alu_loop_op_11_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0,
          alu_loop_op_11_FpAdd_8U_23U_b_left_shift_acc_itm, and_dcpl_241);
      alu_loop_op_11_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_b_right_shift_qr_11_lpi_1_dfm[0]), alu_loop_op_11_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm,
          and_dcpl_241);
      alu_loop_op_11_FpAdd_8U_23U_a_left_shift_acc_itm_2 <= MUX_v_8_2_2(alu_loop_op_11_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0,
          alu_loop_op_11_FpAdd_8U_23U_a_left_shift_acc_itm, and_dcpl_241);
      alu_loop_op_11_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_a_right_shift_qr_11_lpi_1_dfm[0]), alu_loop_op_11_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm,
          and_dcpl_241);
      alu_loop_op_12_FpAdd_8U_23U_b_left_shift_acc_1_itm_2 <= MUX_v_8_2_2(alu_loop_op_12_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0,
          alu_loop_op_12_FpAdd_8U_23U_b_left_shift_acc_1_itm, and_dcpl_241);
      alu_loop_op_12_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_b_right_shift_qr_12_lpi_1_dfm[0]), alu_loop_op_12_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm,
          and_dcpl_241);
      alu_loop_op_12_FpAdd_8U_23U_a_left_shift_acc_1_itm_2 <= MUX_v_8_2_2(alu_loop_op_12_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0,
          alu_loop_op_12_FpAdd_8U_23U_a_left_shift_acc_1_itm, and_dcpl_241);
      alu_loop_op_12_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_a_right_shift_qr_12_lpi_1_dfm[0]), alu_loop_op_12_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm,
          and_dcpl_241);
      alu_loop_op_13_FpAdd_8U_23U_b_left_shift_acc_itm_2 <= MUX_v_8_2_2(alu_loop_op_13_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0,
          alu_loop_op_13_FpAdd_8U_23U_b_left_shift_acc_itm, and_dcpl_241);
      alu_loop_op_13_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_b_right_shift_qr_13_lpi_1_dfm[0]), alu_loop_op_13_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm,
          and_dcpl_241);
      alu_loop_op_13_FpAdd_8U_23U_a_left_shift_acc_itm_2 <= MUX_v_8_2_2(alu_loop_op_13_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0,
          alu_loop_op_13_FpAdd_8U_23U_a_left_shift_acc_itm, and_dcpl_241);
      alu_loop_op_13_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_a_right_shift_qr_13_lpi_1_dfm[0]), alu_loop_op_13_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm,
          and_dcpl_241);
      alu_loop_op_14_FpAdd_8U_23U_b_left_shift_acc_1_itm_2 <= MUX_v_8_2_2(alu_loop_op_14_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0,
          alu_loop_op_14_FpAdd_8U_23U_b_left_shift_acc_1_itm, and_dcpl_241);
      alu_loop_op_14_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_b_right_shift_qr_14_lpi_1_dfm[0]), alu_loop_op_14_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm,
          and_dcpl_241);
      alu_loop_op_14_FpAdd_8U_23U_a_left_shift_acc_1_itm_2 <= MUX_v_8_2_2(alu_loop_op_14_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0,
          alu_loop_op_14_FpAdd_8U_23U_a_left_shift_acc_1_itm, and_dcpl_241);
      alu_loop_op_14_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_a_right_shift_qr_14_lpi_1_dfm[0]), alu_loop_op_14_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm,
          and_dcpl_241);
      alu_loop_op_15_FpAdd_8U_23U_b_left_shift_acc_itm_2 <= MUX_v_8_2_2(alu_loop_op_15_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0,
          alu_loop_op_15_FpAdd_8U_23U_b_left_shift_acc_itm, and_dcpl_241);
      alu_loop_op_15_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_b_right_shift_qr_15_lpi_1_dfm[0]), alu_loop_op_15_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm,
          and_dcpl_241);
      alu_loop_op_15_FpAdd_8U_23U_a_left_shift_acc_itm_2 <= MUX_v_8_2_2(alu_loop_op_15_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0,
          alu_loop_op_15_FpAdd_8U_23U_a_left_shift_acc_itm, and_dcpl_241);
      alu_loop_op_15_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_a_right_shift_qr_15_lpi_1_dfm[0]), alu_loop_op_15_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm,
          and_dcpl_241);
      alu_loop_op_16_FpAdd_8U_23U_b_left_shift_acc_1_itm_2 <= MUX_v_8_2_2(alu_loop_op_16_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0,
          alu_loop_op_16_FpAdd_8U_23U_b_left_shift_acc_1_itm, and_dcpl_241);
      alu_loop_op_16_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm[0]), alu_loop_op_16_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm,
          and_dcpl_241);
      alu_loop_op_16_FpAdd_8U_23U_a_left_shift_acc_1_itm_2 <= MUX_v_8_2_2(alu_loop_op_16_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0,
          alu_loop_op_16_FpAdd_8U_23U_a_left_shift_acc_1_itm, and_dcpl_241);
      alu_loop_op_16_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm_2
          <= MUX_s_1_2_2((FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm[0]), alu_loop_op_16_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm,
          and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      AluIn_data_sva_502 <= 512'b0;
      io_read_cfg_alu_bypass_rsc_svs_st_6 <= 1'b0;
      alu_loop_op_else_nor_tmp_81 <= 1'b0;
    end
    else if ( AluIn_data_and_2_cse ) begin
      AluIn_data_sva_502 <= AluIn_data_sva_501;
      io_read_cfg_alu_bypass_rsc_svs_st_6 <= io_read_cfg_alu_bypass_rsc_svs_st_5;
      alu_loop_op_else_nor_tmp_81 <= alu_loop_op_else_nor_tmp_80;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
          <= 1'b0;
      reg_alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
          <= 1'b0;
      reg_alu_loop_op_5_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
          <= 1'b0;
      reg_alu_loop_op_11_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
          <= 1'b0;
      reg_alu_loop_op_12_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
          <= 1'b0;
    end
    else if ( FpAdd_8U_23U_is_addition_and_33_cse ) begin
      reg_alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
          <= alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3;
      reg_alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
          <= alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3;
      reg_alu_loop_op_5_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
          <= alu_loop_op_5_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
      reg_alu_loop_op_11_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
          <= alu_loop_op_11_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
      reg_alu_loop_op_12_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_2_cse
          <= alu_loop_op_12_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (~ (mux_172_nl)) ) begin
      reg_alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_2_cse
          <= alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_algo_1_sva_st_204 <= 2'b0;
      reg_cfg_alu_algo_1_sva_st_110_cse <= 2'b0;
      cfg_alu_algo_1_sva_6 <= 2'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp_2 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_78_cse ) begin
      cfg_alu_algo_1_sva_st_204 <= reg_cfg_alu_algo_1_sva_st_93_cse;
      reg_cfg_alu_algo_1_sva_st_110_cse <= reg_cfg_alu_algo_1_sva_st_157_cse;
      cfg_alu_algo_1_sva_6 <= cfg_alu_algo_1_sva_5;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp_2;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_4 <= 1'b0;
    end
    else if ( core_wen & ((or_cse_2 & main_stage_v_3) | main_stage_v_4_mx0c1) ) begin
      main_stage_v_4 <= ~ main_stage_v_4_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_22_0_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((((FpCmp_8U_23U_false_is_a_greater_lpi_1_dfm_7 & (~ IsNaN_8U_23U_3_land_lpi_1_dfm_7))
        | IsNaN_8U_23U_1_land_lpi_1_dfm_8) & or_cse_2) | and_715_rgt) & mux_250_cse
        ) begin
      FpCmp_8U_23U_true_o_22_0_lpi_1_dfm_6 <= MUX_v_23_2_2((AluIn_data_sva_502[502:480]),
          ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp_2}), and_715_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_22_0_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((or_cse_2 & (FpCmp_8U_23U_false_is_a_greater_lpi_1_dfm_7
        | IsNaN_8U_23U_3_land_lpi_1_dfm_7) & (~ IsNaN_8U_23U_1_land_lpi_1_dfm_8))
        | and_719_rgt) & mux_251_cse ) begin
      FpCmp_8U_23U_false_o_22_0_lpi_1_dfm_6 <= MUX_v_23_2_2(({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp_2}),
          (AluIn_data_sva_502[502:480]), and_719_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_22_0_15_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & (((((~ IsNaN_8U_23U_3_land_15_lpi_1_dfm_7) & FpCmp_8U_23U_false_is_a_greater_15_lpi_1_dfm_7)
        | IsNaN_8U_23U_1_land_15_lpi_1_dfm_8) & or_cse_2) | and_723_rgt) & mux_250_cse
        ) begin
      FpCmp_8U_23U_true_o_22_0_15_lpi_1_dfm_6 <= MUX_v_23_2_2((AluIn_data_sva_502[470:448]),
          ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp_2}), and_723_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_22_0_15_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((and_dcpl_256 & (IsNaN_8U_23U_3_land_15_lpi_1_dfm_7 | FpCmp_8U_23U_false_is_a_greater_15_lpi_1_dfm_7))
        | and_726_rgt) & mux_251_cse ) begin
      FpCmp_8U_23U_false_o_22_0_15_lpi_1_dfm_6 <= MUX_v_23_2_2(({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp_2}),
          (AluIn_data_sva_502[470:448]), and_726_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_22_0_14_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((((FpCmp_8U_23U_false_is_a_greater_14_lpi_1_dfm_7 & (~
        IsNaN_8U_23U_3_land_14_lpi_1_dfm_7)) | IsNaN_8U_23U_2_land_14_lpi_1_dfm_8)
        & or_cse_2) | and_730_rgt) & mux_250_cse ) begin
      FpCmp_8U_23U_true_o_22_0_14_lpi_1_dfm_6 <= MUX_v_23_2_2((AluIn_data_sva_502[438:416]),
          ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp_2}), and_730_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_22_0_14_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((and_dcpl_263 & (FpCmp_8U_23U_false_is_a_greater_14_lpi_1_dfm_7
        | IsNaN_8U_23U_3_land_14_lpi_1_dfm_7)) | and_733_rgt) & mux_251_cse ) begin
      FpCmp_8U_23U_false_o_22_0_14_lpi_1_dfm_6 <= MUX_v_23_2_2(({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp_2}),
          (AluIn_data_sva_502[438:416]), and_733_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_22_0_13_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((((FpCmp_8U_23U_false_is_a_greater_13_lpi_1_dfm_7 & (~
        IsNaN_8U_23U_3_land_13_lpi_1_dfm_7)) | IsNaN_8U_23U_2_land_13_lpi_1_dfm_8)
        & or_cse_2) | and_737_rgt) & mux_250_cse ) begin
      FpCmp_8U_23U_true_o_22_0_13_lpi_1_dfm_6 <= MUX_v_23_2_2((AluIn_data_sva_502[406:384]),
          ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp_2}), and_737_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_22_0_13_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((or_cse_2 & (FpCmp_8U_23U_false_is_a_greater_13_lpi_1_dfm_7
        | IsNaN_8U_23U_3_land_13_lpi_1_dfm_7) & (~ IsNaN_8U_23U_2_land_13_lpi_1_dfm_8))
        | and_741_rgt) & mux_251_cse ) begin
      FpCmp_8U_23U_false_o_22_0_13_lpi_1_dfm_6 <= MUX_v_23_2_2(({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp_2}),
          (AluIn_data_sva_502[406:384]), and_741_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_22_0_12_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & (((((~ IsNaN_8U_23U_3_land_12_lpi_1_dfm_7) & FpCmp_8U_23U_false_is_a_greater_12_lpi_1_dfm_7)
        | IsNaN_8U_23U_2_land_12_lpi_1_dfm_8) & or_cse_2) | and_745_rgt) & mux_250_cse
        ) begin
      FpCmp_8U_23U_true_o_22_0_12_lpi_1_dfm_6 <= MUX_v_23_2_2((AluIn_data_sva_502[374:352]),
          ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp_2}), and_745_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_22_0_12_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((or_cse_2 & (IsNaN_8U_23U_3_land_12_lpi_1_dfm_7 | FpCmp_8U_23U_false_is_a_greater_12_lpi_1_dfm_7)
        & (~ IsNaN_8U_23U_2_land_12_lpi_1_dfm_8)) | and_749_rgt) & mux_251_cse )
        begin
      FpCmp_8U_23U_false_o_22_0_12_lpi_1_dfm_6 <= MUX_v_23_2_2(({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp_2}),
          (AluIn_data_sva_502[374:352]), and_749_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_22_0_11_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((((FpCmp_8U_23U_false_is_a_greater_11_lpi_1_dfm_7 & (~
        IsNaN_8U_23U_3_land_11_lpi_1_dfm_7)) | IsNaN_8U_23U_2_land_11_lpi_1_dfm_8)
        & or_cse_2) | and_753_rgt) & mux_250_cse ) begin
      FpCmp_8U_23U_true_o_22_0_11_lpi_1_dfm_6 <= MUX_v_23_2_2((AluIn_data_sva_502[342:320]),
          ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp_2}), and_753_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_22_0_11_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((or_cse_2 & (FpCmp_8U_23U_false_is_a_greater_11_lpi_1_dfm_7
        | IsNaN_8U_23U_3_land_11_lpi_1_dfm_7) & (~ IsNaN_8U_23U_2_land_11_lpi_1_dfm_8))
        | and_757_rgt) & mux_251_cse ) begin
      FpCmp_8U_23U_false_o_22_0_11_lpi_1_dfm_6 <= MUX_v_23_2_2(({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp_2}),
          (AluIn_data_sva_502[342:320]), and_757_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_22_0_10_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & (((((~ IsNaN_8U_23U_3_land_10_lpi_1_dfm_7) & FpCmp_8U_23U_false_is_a_greater_10_lpi_1_dfm_7)
        | IsNaN_8U_23U_2_land_10_lpi_1_dfm_8) & or_cse_2) | and_761_rgt) & mux_250_cse
        ) begin
      FpCmp_8U_23U_true_o_22_0_10_lpi_1_dfm_6 <= MUX_v_23_2_2((AluIn_data_sva_502[310:288]),
          ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp_2}), and_761_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_22_0_10_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((and_dcpl_294 & (IsNaN_8U_23U_3_land_10_lpi_1_dfm_7 | FpCmp_8U_23U_false_is_a_greater_10_lpi_1_dfm_7))
        | and_764_rgt) & mux_251_cse ) begin
      FpCmp_8U_23U_false_o_22_0_10_lpi_1_dfm_6 <= MUX_v_23_2_2(({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp_2}),
          (AluIn_data_sva_502[310:288]), and_764_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_22_0_9_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((((FpCmp_8U_23U_false_is_a_greater_9_lpi_1_dfm_7 & (~ IsNaN_8U_23U_3_land_9_lpi_1_dfm_7))
        | IsNaN_8U_23U_2_land_9_lpi_1_dfm_8) & or_cse_2) | and_768_rgt) & mux_250_cse
        ) begin
      FpCmp_8U_23U_true_o_22_0_9_lpi_1_dfm_6 <= MUX_v_23_2_2((AluIn_data_sva_502[278:256]),
          ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp_2}), and_768_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_22_0_9_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((or_cse_2 & (FpCmp_8U_23U_false_is_a_greater_9_lpi_1_dfm_7
        | IsNaN_8U_23U_3_land_9_lpi_1_dfm_7) & (~ IsNaN_8U_23U_2_land_9_lpi_1_dfm_8))
        | and_772_rgt) & mux_251_cse ) begin
      FpCmp_8U_23U_false_o_22_0_9_lpi_1_dfm_6 <= MUX_v_23_2_2(({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp_2}),
          (AluIn_data_sva_502[278:256]), and_772_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_22_0_8_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((((FpCmp_8U_23U_false_is_a_greater_8_lpi_1_dfm_7 & (~ IsNaN_8U_23U_3_land_8_lpi_1_dfm_7))
        | IsNaN_8U_23U_1_land_8_lpi_1_dfm_8) & or_cse_2) | and_776_rgt) & mux_250_cse
        ) begin
      FpCmp_8U_23U_true_o_22_0_8_lpi_1_dfm_6 <= MUX_v_23_2_2((AluIn_data_sva_502[246:224]),
          ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp_2}), and_776_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_22_0_8_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((and_dcpl_309 & (FpCmp_8U_23U_false_is_a_greater_8_lpi_1_dfm_7
        | IsNaN_8U_23U_3_land_8_lpi_1_dfm_7)) | and_779_rgt) & mux_251_cse ) begin
      FpCmp_8U_23U_false_o_22_0_8_lpi_1_dfm_6 <= MUX_v_23_2_2(({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp_2}),
          (AluIn_data_sva_502[246:224]), and_779_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_22_0_7_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & (((((~ IsNaN_8U_23U_3_land_7_lpi_1_dfm_7) & FpCmp_8U_23U_false_is_a_greater_7_lpi_1_dfm_7)
        | IsNaN_8U_23U_1_land_7_lpi_1_dfm_8) & or_cse_2) | and_783_rgt) & mux_250_cse
        ) begin
      FpCmp_8U_23U_true_o_22_0_7_lpi_1_dfm_6 <= MUX_v_23_2_2((AluIn_data_sva_502[214:192]),
          ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp_2}), and_783_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_22_0_7_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((and_dcpl_316 & (IsNaN_8U_23U_3_land_7_lpi_1_dfm_7 | FpCmp_8U_23U_false_is_a_greater_7_lpi_1_dfm_7))
        | and_786_rgt) & mux_251_cse ) begin
      FpCmp_8U_23U_false_o_22_0_7_lpi_1_dfm_6 <= MUX_v_23_2_2(({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp_2}),
          (AluIn_data_sva_502[214:192]), and_786_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_22_0_6_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & (((((~ IsNaN_8U_23U_3_land_6_lpi_1_dfm_7) & FpCmp_8U_23U_false_is_a_greater_6_lpi_1_dfm_7)
        | IsNaN_8U_23U_2_land_6_lpi_1_dfm_8) & or_cse_2) | and_790_rgt) & mux_250_cse
        ) begin
      FpCmp_8U_23U_true_o_22_0_6_lpi_1_dfm_6 <= MUX_v_23_2_2((AluIn_data_sva_502[182:160]),
          ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp_2}), and_790_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_22_0_6_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((or_cse_2 & (IsNaN_8U_23U_3_land_6_lpi_1_dfm_7 | FpCmp_8U_23U_false_is_a_greater_6_lpi_1_dfm_7)
        & (~ IsNaN_8U_23U_2_land_6_lpi_1_dfm_8)) | and_794_rgt) & mux_251_cse ) begin
      FpCmp_8U_23U_false_o_22_0_6_lpi_1_dfm_6 <= MUX_v_23_2_2(({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp_2}),
          (AluIn_data_sva_502[182:160]), and_794_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_22_0_5_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & (((((~ IsNaN_8U_23U_3_land_5_lpi_1_dfm_7) & FpCmp_8U_23U_false_is_a_greater_5_lpi_1_dfm_7)
        | IsNaN_8U_23U_2_land_5_lpi_1_dfm_8) & or_cse_2) | and_798_rgt) & mux_250_cse
        ) begin
      FpCmp_8U_23U_true_o_22_0_5_lpi_1_dfm_6 <= MUX_v_23_2_2((AluIn_data_sva_502[150:128]),
          ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp_2}), and_798_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_22_0_5_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((or_cse_2 & (IsNaN_8U_23U_3_land_5_lpi_1_dfm_7 | FpCmp_8U_23U_false_is_a_greater_5_lpi_1_dfm_7)
        & (~ IsNaN_8U_23U_2_land_5_lpi_1_dfm_8)) | and_802_rgt) & mux_251_cse ) begin
      FpCmp_8U_23U_false_o_22_0_5_lpi_1_dfm_6 <= MUX_v_23_2_2(({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp_2}),
          (AluIn_data_sva_502[150:128]), and_802_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_22_0_4_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((((FpCmp_8U_23U_false_is_a_greater_4_lpi_1_dfm_7 & (~ IsNaN_8U_23U_3_land_4_lpi_1_dfm_7))
        | IsNaN_8U_23U_2_land_4_lpi_1_dfm_8) & or_cse_2) | and_806_rgt) & mux_250_cse
        ) begin
      FpCmp_8U_23U_true_o_22_0_4_lpi_1_dfm_6 <= MUX_v_23_2_2((AluIn_data_sva_502[118:96]),
          ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp_2}), and_806_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_22_0_4_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((or_cse_2 & (FpCmp_8U_23U_false_is_a_greater_4_lpi_1_dfm_7
        | IsNaN_8U_23U_3_land_4_lpi_1_dfm_7) & (~ IsNaN_8U_23U_2_land_4_lpi_1_dfm_8))
        | and_810_rgt) & mux_251_cse ) begin
      FpCmp_8U_23U_false_o_22_0_4_lpi_1_dfm_6 <= MUX_v_23_2_2(({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp_2}),
          (AluIn_data_sva_502[118:96]), and_810_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_22_0_3_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & (((((~ IsNaN_8U_23U_3_land_3_lpi_1_dfm_7) & FpCmp_8U_23U_false_is_a_greater_3_lpi_1_dfm_7)
        | IsNaN_8U_23U_1_land_3_lpi_1_dfm_8) & or_cse_2) | and_814_rgt) & mux_250_cse
        ) begin
      FpCmp_8U_23U_true_o_22_0_3_lpi_1_dfm_6 <= MUX_v_23_2_2((AluIn_data_sva_502[86:64]),
          ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp_2}), and_814_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_22_0_3_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((and_dcpl_347 & (IsNaN_8U_23U_3_land_3_lpi_1_dfm_7 | FpCmp_8U_23U_false_is_a_greater_3_lpi_1_dfm_7))
        | and_817_rgt) & mux_251_cse ) begin
      FpCmp_8U_23U_false_o_22_0_3_lpi_1_dfm_6 <= MUX_v_23_2_2(({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp_2}),
          (AluIn_data_sva_502[86:64]), and_817_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_22_0_2_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((((FpCmp_8U_23U_false_is_a_greater_2_lpi_1_dfm_7 & (~ IsNaN_8U_23U_3_land_2_lpi_1_dfm_7))
        | IsNaN_8U_23U_2_land_2_lpi_1_dfm_8) & or_cse_2) | and_821_rgt) & mux_250_cse
        ) begin
      FpCmp_8U_23U_true_o_22_0_2_lpi_1_dfm_6 <= MUX_v_23_2_2((AluIn_data_sva_502[54:32]),
          ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp_2}), and_821_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_22_0_2_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((and_dcpl_354 & (FpCmp_8U_23U_false_is_a_greater_2_lpi_1_dfm_7
        | IsNaN_8U_23U_3_land_2_lpi_1_dfm_7)) | and_824_rgt) & mux_251_cse ) begin
      FpCmp_8U_23U_false_o_22_0_2_lpi_1_dfm_6 <= MUX_v_23_2_2(({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp_2}),
          (AluIn_data_sva_502[54:32]), and_824_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_22_0_1_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & (((((~ IsNaN_8U_23U_3_land_1_lpi_1_dfm_7) & FpCmp_8U_23U_false_is_a_greater_1_lpi_1_dfm_7)
        | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8) & or_cse_2) | and_828_rgt) & mux_250_cse
        ) begin
      FpCmp_8U_23U_true_o_22_0_1_lpi_1_dfm_6 <= MUX_v_23_2_2((AluIn_data_sva_502[22:0]),
          ({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp_2}), and_828_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_22_0_1_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((and_dcpl_361 & (IsNaN_8U_23U_3_land_1_lpi_1_dfm_7 | FpCmp_8U_23U_false_is_a_greater_1_lpi_1_dfm_7))
        | and_831_rgt) & mux_251_cse ) begin
      FpCmp_8U_23U_false_o_22_0_1_lpi_1_dfm_6 <= MUX_v_23_2_2(({reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp_1 , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp_2}),
          (AluIn_data_sva_502[22:0]), and_831_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_45_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_47_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_46_itm_4 <= 30'b0;
      alu_loop_op_else_else_if_mux_42_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_44_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_43_itm_4 <= 30'b0;
      alu_loop_op_else_else_if_mux_39_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_41_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_40_itm_4 <= 30'b0;
      alu_loop_op_else_else_if_mux_6_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_8_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_7_itm_4 <= 30'b0;
      alu_loop_op_else_else_if_mux_36_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_38_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_37_itm_4 <= 30'b0;
      alu_loop_op_else_else_if_mux_33_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_35_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_34_itm_4 <= 30'b0;
      alu_loop_op_else_else_if_mux_12_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_14_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_13_itm_4 <= 30'b0;
      alu_loop_op_else_else_if_mux_30_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_32_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_31_itm_4 <= 30'b0;
      alu_loop_op_else_else_if_mux_15_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_17_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_16_itm_4 <= 30'b0;
      alu_loop_op_else_else_if_mux_27_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_29_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_28_itm_4 <= 30'b0;
      alu_loop_op_else_else_if_mux_18_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_20_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_19_itm_4 <= 30'b0;
      alu_loop_op_else_else_if_mux_24_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_26_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_25_itm_4 <= 30'b0;
      alu_loop_op_else_else_if_mux_21_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_23_itm_4 <= 1'b0;
      alu_loop_op_else_else_if_mux_22_itm_4 <= 30'b0;
    end
    else if ( alu_loop_op_else_else_if_and_57_cse ) begin
      alu_loop_op_else_else_if_mux_45_itm_4 <= alu_loop_op_else_else_if_mux_45_itm_3;
      alu_loop_op_else_else_if_mux_47_itm_4 <= alu_loop_op_else_else_if_mux_47_itm_3;
      alu_loop_op_else_else_if_mux_46_itm_4 <= alu_loop_op_else_else_if_mux_46_itm_3;
      alu_loop_op_else_else_if_mux_42_itm_4 <= alu_loop_op_else_else_if_mux_42_itm_3;
      alu_loop_op_else_else_if_mux_44_itm_4 <= alu_loop_op_else_else_if_mux_44_itm_3;
      alu_loop_op_else_else_if_mux_43_itm_4 <= alu_loop_op_else_else_if_mux_43_itm_3;
      alu_loop_op_else_else_if_mux_39_itm_4 <= alu_loop_op_else_else_if_mux_39_itm_3;
      alu_loop_op_else_else_if_mux_41_itm_4 <= alu_loop_op_else_else_if_mux_41_itm_3;
      alu_loop_op_else_else_if_mux_40_itm_4 <= alu_loop_op_else_else_if_mux_40_itm_3;
      alu_loop_op_else_else_if_mux_6_itm_4 <= alu_loop_op_else_else_if_mux_6_itm_3;
      alu_loop_op_else_else_if_mux_8_itm_4 <= alu_loop_op_else_else_if_mux_8_itm_3;
      alu_loop_op_else_else_if_mux_7_itm_4 <= alu_loop_op_else_else_if_mux_7_itm_3;
      alu_loop_op_else_else_if_mux_36_itm_4 <= alu_loop_op_else_else_if_mux_36_itm_3;
      alu_loop_op_else_else_if_mux_38_itm_4 <= alu_loop_op_else_else_if_mux_38_itm_3;
      alu_loop_op_else_else_if_mux_37_itm_4 <= alu_loop_op_else_else_if_mux_37_itm_3;
      alu_loop_op_else_else_if_mux_33_itm_4 <= alu_loop_op_else_else_if_mux_33_itm_3;
      alu_loop_op_else_else_if_mux_35_itm_4 <= alu_loop_op_else_else_if_mux_35_itm_3;
      alu_loop_op_else_else_if_mux_34_itm_4 <= alu_loop_op_else_else_if_mux_34_itm_3;
      alu_loop_op_else_else_if_mux_12_itm_4 <= alu_loop_op_else_else_if_mux_12_itm_3;
      alu_loop_op_else_else_if_mux_14_itm_4 <= alu_loop_op_else_else_if_mux_14_itm_3;
      alu_loop_op_else_else_if_mux_13_itm_4 <= alu_loop_op_else_else_if_mux_13_itm_3;
      alu_loop_op_else_else_if_mux_30_itm_4 <= alu_loop_op_else_else_if_mux_30_itm_3;
      alu_loop_op_else_else_if_mux_32_itm_4 <= alu_loop_op_else_else_if_mux_32_itm_3;
      alu_loop_op_else_else_if_mux_31_itm_4 <= alu_loop_op_else_else_if_mux_31_itm_3;
      alu_loop_op_else_else_if_mux_15_itm_4 <= alu_loop_op_else_else_if_mux_15_itm_3;
      alu_loop_op_else_else_if_mux_17_itm_4 <= alu_loop_op_else_else_if_mux_17_itm_3;
      alu_loop_op_else_else_if_mux_16_itm_4 <= alu_loop_op_else_else_if_mux_16_itm_3;
      alu_loop_op_else_else_if_mux_27_itm_4 <= alu_loop_op_else_else_if_mux_27_itm_3;
      alu_loop_op_else_else_if_mux_29_itm_4 <= alu_loop_op_else_else_if_mux_29_itm_3;
      alu_loop_op_else_else_if_mux_28_itm_4 <= alu_loop_op_else_else_if_mux_28_itm_3;
      alu_loop_op_else_else_if_mux_18_itm_4 <= alu_loop_op_else_else_if_mux_18_itm_3;
      alu_loop_op_else_else_if_mux_20_itm_4 <= alu_loop_op_else_else_if_mux_20_itm_3;
      alu_loop_op_else_else_if_mux_19_itm_4 <= alu_loop_op_else_else_if_mux_19_itm_3;
      alu_loop_op_else_else_if_mux_24_itm_4 <= alu_loop_op_else_else_if_mux_24_itm_3;
      alu_loop_op_else_else_if_mux_26_itm_4 <= alu_loop_op_else_else_if_mux_26_itm_3;
      alu_loop_op_else_else_if_mux_25_itm_4 <= alu_loop_op_else_else_if_mux_25_itm_3;
      alu_loop_op_else_else_if_mux_21_itm_4 <= alu_loop_op_else_else_if_mux_21_itm_3;
      alu_loop_op_else_else_if_mux_23_itm_4 <= alu_loop_op_else_else_if_mux_23_itm_3;
      alu_loop_op_else_else_if_mux_22_itm_4 <= alu_loop_op_else_else_if_mux_22_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_else_else_if_conc_itm_1_31_1 <= 1'b0;
      alu_loop_op_1_else_else_if_conc_itm_1_0_1 <= 1'b0;
      alu_loop_op_1_else_else_if_conc_itm_1_30_1_1 <= 30'b0;
    end
    else if ( alu_loop_op_else_else_if_and_60_cse ) begin
      alu_loop_op_1_else_else_if_conc_itm_1_31_1 <= MUX1HOT_s_1_3_2(alu_loop_op_else_else_if_mux_itm_2,
          alu_loop_op_1_else_else_if_conc_itm_31, alu_loop_op_1_else_if_conc_itm_31,
          {and_dcpl_369 , and_dcpl_372 , and_dcpl_375});
      alu_loop_op_1_else_else_if_conc_itm_1_0_1 <= MUX1HOT_s_1_3_2(alu_loop_op_else_else_if_mux_2_itm_2,
          alu_loop_op_1_else_else_if_conc_itm_0, alu_loop_op_1_else_if_conc_itm_0,
          {and_dcpl_369 , and_dcpl_372 , and_dcpl_375});
      alu_loop_op_1_else_else_if_conc_itm_1_30_1_1 <= MUX1HOT_v_30_3_2(alu_loop_op_else_else_if_mux_1_itm_2,
          alu_loop_op_1_else_else_if_conc_itm_30_1, alu_loop_op_1_else_if_conc_itm_30_1,
          {and_dcpl_369 , and_dcpl_372 , and_dcpl_375});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_2_else_else_if_conc_1_itm_1_31_1 <= 1'b0;
      alu_loop_op_2_else_else_if_conc_1_itm_1_0_1 <= 1'b0;
      alu_loop_op_2_else_else_if_conc_1_itm_1_30_1_1 <= 30'b0;
      alu_loop_op_4_else_else_if_conc_1_itm_1_31_1 <= 1'b0;
      alu_loop_op_4_else_else_if_conc_1_itm_1_0_1 <= 1'b0;
      alu_loop_op_4_else_else_if_conc_1_itm_1_30_1_1 <= 30'b0;
    end
    else if ( alu_loop_op_else_else_if_and_66_cse ) begin
      alu_loop_op_2_else_else_if_conc_1_itm_1_31_1 <= MUX1HOT_s_1_3_2(alu_loop_op_else_else_if_mux_3_itm_2,
          alu_loop_op_2_else_else_if_conc_1_itm_31, alu_loop_op_2_else_if_conc_1_itm_31,
          {and_dcpl_379 , and_dcpl_372 , and_dcpl_375});
      alu_loop_op_2_else_else_if_conc_1_itm_1_0_1 <= MUX1HOT_s_1_3_2(alu_loop_op_else_else_if_mux_5_itm_2,
          alu_loop_op_2_else_else_if_conc_1_itm_0, alu_loop_op_2_else_if_conc_1_itm_0,
          {and_dcpl_379 , and_dcpl_372 , and_dcpl_375});
      alu_loop_op_2_else_else_if_conc_1_itm_1_30_1_1 <= MUX1HOT_v_30_3_2(alu_loop_op_else_else_if_mux_4_itm_2,
          alu_loop_op_2_else_else_if_conc_1_itm_30_1, alu_loop_op_2_else_if_conc_1_itm_30_1,
          {and_dcpl_379 , and_dcpl_372 , and_dcpl_375});
      alu_loop_op_4_else_else_if_conc_1_itm_1_31_1 <= MUX1HOT_s_1_3_2(alu_loop_op_else_else_if_mux_9_itm_2,
          alu_loop_op_4_else_else_if_conc_1_itm_31, alu_loop_op_4_else_if_conc_1_itm_31,
          {and_dcpl_379 , and_dcpl_372 , and_dcpl_375});
      alu_loop_op_4_else_else_if_conc_1_itm_1_0_1 <= MUX1HOT_s_1_3_2(alu_loop_op_else_else_if_mux_11_itm_2,
          alu_loop_op_4_else_else_if_conc_1_itm_0, alu_loop_op_4_else_if_conc_1_itm_0,
          {and_dcpl_379 , and_dcpl_372 , and_dcpl_375});
      alu_loop_op_4_else_else_if_conc_1_itm_1_30_1_1 <= MUX1HOT_v_30_3_2(alu_loop_op_else_else_if_mux_10_itm_2,
          alu_loop_op_4_else_else_if_conc_1_itm_30_1, alu_loop_op_4_else_if_conc_1_itm_30_1,
          {and_dcpl_379 , and_dcpl_372 , and_dcpl_375});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_and_60_itm_4 <= 1'b0;
      FpAlu_8U_23U_and_itm_4 <= 1'b0;
      FpAlu_8U_23U_and_56_itm_4 <= 1'b0;
      FpAlu_8U_23U_and_4_itm_4 <= 1'b0;
      FpAlu_8U_23U_and_52_itm_4 <= 1'b0;
      FpAlu_8U_23U_and_8_itm_4 <= 1'b0;
      FpAlu_8U_23U_and_48_itm_4 <= 1'b0;
      FpAlu_8U_23U_and_12_itm_4 <= 1'b0;
      FpAlu_8U_23U_and_44_itm_4 <= 1'b0;
      FpAlu_8U_23U_and_16_itm_4 <= 1'b0;
      FpAlu_8U_23U_and_40_itm_4 <= 1'b0;
      FpAlu_8U_23U_and_20_itm_4 <= 1'b0;
      FpAlu_8U_23U_and_36_itm_4 <= 1'b0;
      FpAlu_8U_23U_and_24_itm_4 <= 1'b0;
      FpAlu_8U_23U_and_32_itm_4 <= 1'b0;
      FpAlu_8U_23U_and_28_itm_4 <= 1'b0;
    end
    else if ( FpAlu_8U_23U_and_832_cse ) begin
      FpAlu_8U_23U_and_60_itm_4 <= FpAlu_8U_23U_and_60_itm_3;
      FpAlu_8U_23U_and_itm_4 <= FpAlu_8U_23U_and_itm_3;
      FpAlu_8U_23U_and_56_itm_4 <= FpAlu_8U_23U_and_56_itm_3;
      FpAlu_8U_23U_and_4_itm_4 <= FpAlu_8U_23U_and_4_itm_3;
      FpAlu_8U_23U_and_52_itm_4 <= FpAlu_8U_23U_and_52_itm_3;
      FpAlu_8U_23U_and_8_itm_4 <= FpAlu_8U_23U_and_8_itm_3;
      FpAlu_8U_23U_and_48_itm_4 <= FpAlu_8U_23U_and_48_itm_3;
      FpAlu_8U_23U_and_12_itm_4 <= FpAlu_8U_23U_and_12_itm_3;
      FpAlu_8U_23U_and_44_itm_4 <= FpAlu_8U_23U_and_44_itm_3;
      FpAlu_8U_23U_and_16_itm_4 <= FpAlu_8U_23U_and_16_itm_3;
      FpAlu_8U_23U_and_40_itm_4 <= FpAlu_8U_23U_and_40_itm_3;
      FpAlu_8U_23U_and_20_itm_4 <= FpAlu_8U_23U_and_20_itm_3;
      FpAlu_8U_23U_and_36_itm_4 <= FpAlu_8U_23U_and_36_itm_3;
      FpAlu_8U_23U_and_24_itm_4 <= FpAlu_8U_23U_and_24_itm_3;
      FpAlu_8U_23U_and_32_itm_4 <= FpAlu_8U_23U_and_32_itm_3;
      FpAlu_8U_23U_and_28_itm_4 <= FpAlu_8U_23U_and_28_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      AluOut_data_15_sva_8 <= 33'b0;
      AluOut_data_0_sva_8 <= 33'b0;
      AluOut_data_14_sva_8 <= 33'b0;
      AluOut_data_1_sva_8 <= 33'b0;
      AluOut_data_13_sva_8 <= 33'b0;
      AluOut_data_2_sva_8 <= 33'b0;
      AluOut_data_12_sva_8 <= 33'b0;
      AluOut_data_3_sva_8 <= 33'b0;
      AluOut_data_11_sva_8 <= 33'b0;
      AluOut_data_4_sva_8 <= 33'b0;
      AluOut_data_10_sva_8 <= 33'b0;
      AluOut_data_5_sva_8 <= 33'b0;
      AluOut_data_9_sva_8 <= 33'b0;
      AluOut_data_6_sva_8 <= 33'b0;
      AluOut_data_8_sva_8 <= 33'b0;
      AluOut_data_7_sva_8 <= 33'b0;
    end
    else if ( AluOut_data_and_cse ) begin
      AluOut_data_15_sva_8 <= AluOut_data_15_sva_7;
      AluOut_data_0_sva_8 <= AluOut_data_0_sva_7;
      AluOut_data_14_sva_8 <= AluOut_data_14_sva_7;
      AluOut_data_1_sva_8 <= AluOut_data_1_sva_7;
      AluOut_data_13_sva_8 <= AluOut_data_13_sva_7;
      AluOut_data_2_sva_8 <= AluOut_data_2_sva_7;
      AluOut_data_12_sva_8 <= AluOut_data_12_sva_7;
      AluOut_data_3_sva_8 <= AluOut_data_3_sva_7;
      AluOut_data_11_sva_8 <= AluOut_data_11_sva_7;
      AluOut_data_4_sva_8 <= AluOut_data_4_sva_7;
      AluOut_data_10_sva_8 <= AluOut_data_10_sva_7;
      AluOut_data_5_sva_8 <= AluOut_data_5_sva_7;
      AluOut_data_9_sva_8 <= AluOut_data_9_sva_7;
      AluOut_data_6_sva_8 <= AluOut_data_6_sva_7;
      AluOut_data_8_sva_8 <= AluOut_data_8_sva_7;
      AluOut_data_7_sva_8 <= AluOut_data_7_sva_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_o_0_sva_7 <= 1'b0;
      FpAlu_8U_23U_o_0_1_sva_7 <= 1'b0;
      FpAlu_8U_23U_o_0_15_sva_7 <= 1'b0;
      FpAlu_8U_23U_o_0_2_sva_7 <= 1'b0;
      FpAlu_8U_23U_o_0_14_sva_7 <= 1'b0;
      FpAlu_8U_23U_o_0_3_sva_7 <= 1'b0;
      FpAlu_8U_23U_o_0_13_sva_7 <= 1'b0;
      FpAlu_8U_23U_o_0_4_sva_7 <= 1'b0;
      FpAlu_8U_23U_o_0_12_sva_7 <= 1'b0;
      FpAlu_8U_23U_o_0_5_sva_7 <= 1'b0;
      FpAlu_8U_23U_o_0_11_sva_7 <= 1'b0;
      FpAlu_8U_23U_o_0_6_sva_7 <= 1'b0;
      FpAlu_8U_23U_o_0_10_sva_7 <= 1'b0;
      FpAlu_8U_23U_o_0_7_sva_7 <= 1'b0;
      FpAlu_8U_23U_o_0_9_sva_7 <= 1'b0;
      FpAlu_8U_23U_o_0_8_sva_7 <= 1'b0;
    end
    else if ( FpAlu_8U_23U_o_and_cse ) begin
      FpAlu_8U_23U_o_0_sva_7 <= FpAlu_8U_23U_o_0_sva_6;
      FpAlu_8U_23U_o_0_1_sva_7 <= FpAlu_8U_23U_o_0_1_sva_6;
      FpAlu_8U_23U_o_0_15_sva_7 <= FpAlu_8U_23U_o_0_15_sva_6;
      FpAlu_8U_23U_o_0_2_sva_7 <= FpAlu_8U_23U_o_0_2_sva_6;
      FpAlu_8U_23U_o_0_14_sva_7 <= FpAlu_8U_23U_o_0_14_sva_6;
      FpAlu_8U_23U_o_0_3_sva_7 <= FpAlu_8U_23U_o_0_3_sva_6;
      FpAlu_8U_23U_o_0_13_sva_7 <= FpAlu_8U_23U_o_0_13_sva_6;
      FpAlu_8U_23U_o_0_4_sva_7 <= FpAlu_8U_23U_o_0_4_sva_6;
      FpAlu_8U_23U_o_0_12_sva_7 <= FpAlu_8U_23U_o_0_12_sva_6;
      FpAlu_8U_23U_o_0_5_sva_7 <= FpAlu_8U_23U_o_0_5_sva_6;
      FpAlu_8U_23U_o_0_11_sva_7 <= FpAlu_8U_23U_o_0_11_sva_6;
      FpAlu_8U_23U_o_0_6_sva_7 <= FpAlu_8U_23U_o_0_6_sva_6;
      FpAlu_8U_23U_o_0_10_sva_7 <= FpAlu_8U_23U_o_0_10_sva_6;
      FpAlu_8U_23U_o_0_7_sva_7 <= FpAlu_8U_23U_o_0_7_sva_6;
      FpAlu_8U_23U_o_0_9_sva_7 <= FpAlu_8U_23U_o_0_9_sva_6;
      FpAlu_8U_23U_o_0_8_sva_7 <= FpAlu_8U_23U_o_0_8_sva_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_386_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_2_lpi_1_dfm_5_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_2_lpi_1_dfm_5_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_176_cse ) begin
      FpAdd_8U_23U_qr_2_lpi_1_dfm_5_7_4_1 <= FpAdd_8U_23U_qr_2_lpi_1_dfm_4_7_4_1;
      FpAdd_8U_23U_qr_2_lpi_1_dfm_5_3_0_1 <= FpAdd_8U_23U_qr_2_lpi_1_dfm_4_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
        & (mux_390_nl) ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_st_3 <= MUX_s_1_2_2(alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_itm_7,
          FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_st_2, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5 <= 50'b0;
      alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 <= 1'b0;
      FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5 <= 50'b0;
      alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 <= 1'b0;
      FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_5 <= 50'b0;
      alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 <= 1'b0;
      FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_5 <= 50'b0;
      alu_loop_op_9_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 <= 1'b0;
      FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_5 <= 50'b0;
      alu_loop_op_13_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_int_mant_p1_and_16_cse ) begin
      FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5 <= MUX_v_50_2_2(FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_mx1,
          FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm, and_dcpl_241);
      alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 <= MUX_s_1_2_2((FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_mx2[49]),
          alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm, and_dcpl_241);
      FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5 <= MUX_v_50_2_2(FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_mx1,
          FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm, and_dcpl_241);
      alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 <= MUX_s_1_2_2((FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_mx2[49]),
          alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm, and_dcpl_241);
      FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_5 <= MUX_v_50_2_2(FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_mx1,
          FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm, and_dcpl_241);
      alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 <= MUX_s_1_2_2((FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_mx2[49]),
          alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm, and_dcpl_241);
      FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_5 <= MUX_v_50_2_2(FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_mx1,
          FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm, and_dcpl_241);
      alu_loop_op_9_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 <= MUX_s_1_2_2((FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_mx2[49]),
          alu_loop_op_9_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm, and_dcpl_241);
      FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_5 <= MUX_v_50_2_2(FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_mx1,
          FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm, and_dcpl_241);
      alu_loop_op_13_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 <= MUX_s_1_2_2((FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_mx2[49]),
          alu_loop_op_13_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_1_sva_2 <= 6'b0;
      FpNormalize_8U_49U_if_or_itm_2 <= 1'b0;
    end
    else if ( IntLeadZero_49U_leading_sign_49_0_rtn_and_cse ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_1_sva_2 <= MUX_v_6_2_2(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_16,
          IntLeadZero_49U_leading_sign_49_0_rtn_1_sva, and_dcpl_241);
      FpNormalize_8U_49U_if_or_itm_2 <= MUX_s_1_2_2(FpNormalize_8U_49U_if_or_itm_mx0w0,
          FpNormalize_8U_49U_if_or_itm, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_397_nl) ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      AluIn_data_sva_503 <= 512'b0;
      FpAlu_8U_23U_nor_dfs_79 <= 1'b0;
      FpAlu_8U_23U_equal_tmp_237 <= 1'b0;
      FpAlu_8U_23U_equal_tmp_235 <= 1'b0;
      FpAlu_8U_23U_equal_tmp_239 <= 1'b0;
      io_read_cfg_alu_bypass_rsc_svs_7 <= 1'b0;
      alu_loop_op_else_nor_tmp_82 <= 1'b0;
    end
    else if ( AluIn_data_and_3_cse ) begin
      AluIn_data_sva_503 <= AluIn_data_sva_502;
      FpAlu_8U_23U_nor_dfs_79 <= FpAlu_8U_23U_nor_dfs_48;
      FpAlu_8U_23U_equal_tmp_237 <= FpAlu_8U_23U_equal_tmp_146;
      FpAlu_8U_23U_equal_tmp_235 <= FpAlu_8U_23U_equal_tmp_144;
      FpAlu_8U_23U_equal_tmp_239 <= FpAlu_8U_23U_equal_tmp_148;
      io_read_cfg_alu_bypass_rsc_svs_7 <= io_read_cfg_alu_bypass_rsc_svs_st_6;
      alu_loop_op_else_nor_tmp_82 <= alu_loop_op_else_nor_tmp_81;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_1_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_4_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_5_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_6_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_7_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_8_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_9_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_10_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_11_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_12_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_13_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_14_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_15_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_10 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_cse ) begin
      IsNaN_8U_23U_land_1_lpi_1_dfm_10 <= IsNaN_8U_23U_land_1_lpi_1_dfm_9;
      IsNaN_8U_23U_land_2_lpi_1_dfm_10 <= IsNaN_8U_23U_land_2_lpi_1_dfm_9;
      IsNaN_8U_23U_land_3_lpi_1_dfm_10 <= IsNaN_8U_23U_land_3_lpi_1_dfm_9;
      IsNaN_8U_23U_land_4_lpi_1_dfm_10 <= IsNaN_8U_23U_land_4_lpi_1_dfm_9;
      IsNaN_8U_23U_land_5_lpi_1_dfm_10 <= IsNaN_8U_23U_land_5_lpi_1_dfm_9;
      IsNaN_8U_23U_land_6_lpi_1_dfm_10 <= IsNaN_8U_23U_land_6_lpi_1_dfm_9;
      IsNaN_8U_23U_land_7_lpi_1_dfm_10 <= IsNaN_8U_23U_land_7_lpi_1_dfm_9;
      IsNaN_8U_23U_land_8_lpi_1_dfm_10 <= IsNaN_8U_23U_land_8_lpi_1_dfm_9;
      IsNaN_8U_23U_land_9_lpi_1_dfm_10 <= IsNaN_8U_23U_land_9_lpi_1_dfm_9;
      IsNaN_8U_23U_land_10_lpi_1_dfm_10 <= IsNaN_8U_23U_land_10_lpi_1_dfm_9;
      IsNaN_8U_23U_land_11_lpi_1_dfm_10 <= IsNaN_8U_23U_land_11_lpi_1_dfm_9;
      IsNaN_8U_23U_land_12_lpi_1_dfm_10 <= IsNaN_8U_23U_land_12_lpi_1_dfm_9;
      IsNaN_8U_23U_land_13_lpi_1_dfm_10 <= IsNaN_8U_23U_land_13_lpi_1_dfm_9;
      IsNaN_8U_23U_land_14_lpi_1_dfm_10 <= IsNaN_8U_23U_land_14_lpi_1_dfm_9;
      IsNaN_8U_23U_land_15_lpi_1_dfm_10 <= IsNaN_8U_23U_land_15_lpi_1_dfm_9;
      IsNaN_8U_23U_land_lpi_1_dfm_10 <= IsNaN_8U_23U_land_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_404_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_5 <= 1'b0;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_2 <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_5 <= 1'b0;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_2 <= 1'b0;
      IsNaN_8U_23U_land_4_lpi_1_dfm_st_5 <= 1'b0;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_4_sva_2 <= 1'b0;
      IsNaN_8U_23U_land_9_lpi_1_dfm_st_5 <= 1'b0;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_9_sva_2 <= 1'b0;
      IsNaN_8U_23U_land_13_lpi_1_dfm_st_5 <= 1'b0;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_13_sva_2 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_16_cse ) begin
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_5 <= IsNaN_8U_23U_3_land_1_lpi_1_dfm_7;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_2 <= alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_5 <= IsNaN_8U_23U_3_land_3_lpi_1_dfm_7;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_2 <= alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
      IsNaN_8U_23U_land_4_lpi_1_dfm_st_5 <= IsNaN_8U_23U_2_land_4_lpi_1_dfm_8;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_4_sva_2 <= alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
      IsNaN_8U_23U_land_9_lpi_1_dfm_st_5 <= IsNaN_8U_23U_2_land_9_lpi_1_dfm_8;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_9_sva_2 <= alu_loop_op_9_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
      IsNaN_8U_23U_land_13_lpi_1_dfm_st_5 <= IsNaN_8U_23U_2_land_13_lpi_1_dfm_8;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_13_sva_2 <= alu_loop_op_13_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_409_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_3_lpi_1_dfm_5_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_3_lpi_1_dfm_5_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_178_cse ) begin
      FpAdd_8U_23U_qr_3_lpi_1_dfm_5_7_4_1 <= FpAdd_8U_23U_qr_3_lpi_1_dfm_4_7_4_1;
      FpAdd_8U_23U_qr_3_lpi_1_dfm_5_3_0_1 <= FpAdd_8U_23U_qr_3_lpi_1_dfm_4_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
        & (mux_413_nl) ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_st_3 <= MUX_s_1_2_2(alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_2_itm_7,
          FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_st_2, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5 <= 50'b0;
      alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 <= 1'b0;
      FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_5 <= 50'b0;
      alu_loop_op_6_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 <= 1'b0;
      FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_5 <= 50'b0;
      alu_loop_op_7_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 <= 1'b0;
      FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_5 <= 50'b0;
      alu_loop_op_8_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 <= 1'b0;
      FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_5 <= 50'b0;
      alu_loop_op_10_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 <= 1'b0;
      FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_5 <= 50'b0;
      alu_loop_op_12_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 <= 1'b0;
      FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_5 <= 50'b0;
      alu_loop_op_14_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 <= 1'b0;
      FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_5 <= 50'b0;
      alu_loop_op_15_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 <= 1'b0;
      FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5 <= 50'b0;
      alu_loop_op_16_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_int_mant_p1_and_17_cse ) begin
      FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5 <= MUX_v_50_2_2(FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_mx1,
          FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm, and_dcpl_241);
      alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 <= MUX_s_1_2_2((FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_mx2[49]),
          alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm, and_dcpl_241);
      FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_5 <= MUX_v_50_2_2(FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_mx1,
          FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm, and_dcpl_241);
      alu_loop_op_6_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 <= MUX_s_1_2_2((FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_mx2[49]),
          alu_loop_op_6_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm, and_dcpl_241);
      FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_5 <= MUX_v_50_2_2(FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_mx1,
          FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm, and_dcpl_241);
      alu_loop_op_7_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 <= MUX_s_1_2_2((FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_mx2[49]),
          alu_loop_op_7_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm, and_dcpl_241);
      FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_5 <= MUX_v_50_2_2(FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_mx1,
          FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm, and_dcpl_241);
      alu_loop_op_8_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 <= MUX_s_1_2_2((FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_mx2[49]),
          alu_loop_op_8_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm, and_dcpl_241);
      FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_5 <= MUX_v_50_2_2(FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_mx1,
          FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm, and_dcpl_241);
      alu_loop_op_10_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 <= MUX_s_1_2_2((FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_mx2[49]),
          alu_loop_op_10_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm, and_dcpl_241);
      FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_5 <= MUX_v_50_2_2(FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_mx1,
          FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm, and_dcpl_241);
      alu_loop_op_12_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 <= MUX_s_1_2_2((FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_mx2[49]),
          alu_loop_op_12_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm, and_dcpl_241);
      FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_5 <= MUX_v_50_2_2(FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_mx1,
          FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm, and_dcpl_241);
      alu_loop_op_14_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 <= MUX_s_1_2_2((FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_mx2[49]),
          alu_loop_op_14_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm, and_dcpl_241);
      FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_5 <= MUX_v_50_2_2(FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_mx1,
          FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm, and_dcpl_241);
      alu_loop_op_15_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 <= MUX_s_1_2_2((FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_mx2[49]),
          alu_loop_op_15_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm, and_dcpl_241);
      FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5 <= MUX_v_50_2_2(FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_mx1,
          FpAdd_8U_23U_int_mant_p1_lpi_1_dfm, and_dcpl_241);
      alu_loop_op_16_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 <= MUX_s_1_2_2((FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_mx2[49]),
          alu_loop_op_16_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_2_sva_2 <= 6'b0;
      FpNormalize_8U_49U_if_or_1_itm_2 <= 1'b0;
    end
    else if ( IntLeadZero_49U_leading_sign_49_0_rtn_and_16_cse ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_2_sva_2 <= MUX_v_6_2_2(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_17,
          IntLeadZero_49U_leading_sign_49_0_rtn_2_sva, and_dcpl_241);
      FpNormalize_8U_49U_if_or_1_itm_2 <= MUX_s_1_2_2(FpNormalize_8U_49U_if_or_1_itm_mx0w0,
          FpNormalize_8U_49U_if_or_1_itm, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_419_nl) ) begin
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_425_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_5 <= 1'b0;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_2 <= 1'b0;
      IsNaN_8U_23U_land_6_lpi_1_dfm_st_5 <= 1'b0;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_6_sva_2 <= 1'b0;
      IsNaN_8U_23U_land_7_lpi_1_dfm_st_5 <= 1'b0;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_7_sva_2 <= 1'b0;
      IsNaN_8U_23U_land_8_lpi_1_dfm_st_5 <= 1'b0;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_8_sva_2 <= 1'b0;
      IsNaN_8U_23U_land_10_lpi_1_dfm_st_5 <= 1'b0;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_10_sva_2 <= 1'b0;
      IsNaN_8U_23U_land_12_lpi_1_dfm_st_5 <= 1'b0;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_12_sva_2 <= 1'b0;
      IsNaN_8U_23U_land_14_lpi_1_dfm_st_5 <= 1'b0;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_14_sva_2 <= 1'b0;
      IsNaN_8U_23U_land_15_lpi_1_dfm_st_5 <= 1'b0;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_15_sva_2 <= 1'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_st_5 <= 1'b0;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_2 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_18_cse ) begin
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_5 <= IsNaN_8U_23U_2_land_2_lpi_1_dfm_8;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_2 <= alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
      IsNaN_8U_23U_land_6_lpi_1_dfm_st_5 <= IsNaN_8U_23U_2_land_6_lpi_1_dfm_8;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_6_sva_2 <= alu_loop_op_6_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
      IsNaN_8U_23U_land_7_lpi_1_dfm_st_5 <= IsNaN_8U_23U_3_land_7_lpi_1_dfm_7;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_7_sva_2 <= alu_loop_op_7_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
      IsNaN_8U_23U_land_8_lpi_1_dfm_st_5 <= IsNaN_8U_23U_3_land_8_lpi_1_dfm_7;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_8_sva_2 <= alu_loop_op_8_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
      IsNaN_8U_23U_land_10_lpi_1_dfm_st_5 <= IsNaN_8U_23U_2_land_10_lpi_1_dfm_8;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_10_sva_2 <= alu_loop_op_10_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
      IsNaN_8U_23U_land_12_lpi_1_dfm_st_5 <= IsNaN_8U_23U_2_land_12_lpi_1_dfm_8;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_12_sva_2 <= alu_loop_op_12_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
      IsNaN_8U_23U_land_14_lpi_1_dfm_st_5 <= IsNaN_8U_23U_2_land_14_lpi_1_dfm_8;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_14_sva_2 <= alu_loop_op_14_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
      IsNaN_8U_23U_land_15_lpi_1_dfm_st_5 <= IsNaN_8U_23U_3_land_15_lpi_1_dfm_7;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_15_sva_2 <= alu_loop_op_15_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
      IsNaN_8U_23U_land_lpi_1_dfm_st_5 <= IsNaN_8U_23U_3_land_lpi_1_dfm_7;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_2 <= alu_loop_op_16_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_430_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_4_lpi_1_dfm_5_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_4_lpi_1_dfm_5_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_180_cse ) begin
      FpAdd_8U_23U_qr_4_lpi_1_dfm_5_7_4_1 <= FpAdd_8U_23U_qr_4_lpi_1_dfm_4_7_4_1;
      FpAdd_8U_23U_qr_4_lpi_1_dfm_5_3_0_1 <= FpAdd_8U_23U_qr_4_lpi_1_dfm_4_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
        & (mux_434_nl) ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_st_3 <= MUX_s_1_2_2(alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_1_itm_7,
          FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_st_2, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_3_sva_2 <= 6'b0;
      FpNormalize_8U_49U_if_or_2_itm_2 <= 1'b0;
    end
    else if ( IntLeadZero_49U_leading_sign_49_0_rtn_and_17_cse ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_3_sva_2 <= MUX_v_6_2_2(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_18,
          IntLeadZero_49U_leading_sign_49_0_rtn_3_sva, and_dcpl_241);
      FpNormalize_8U_49U_if_or_2_itm_2 <= MUX_s_1_2_2(FpNormalize_8U_49U_if_or_2_itm_mx0w0,
          FpNormalize_8U_49U_if_or_2_itm, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_440_nl) ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_446_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_451_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_5_lpi_1_dfm_5_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_5_lpi_1_dfm_5_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_182_cse ) begin
      FpAdd_8U_23U_qr_5_lpi_1_dfm_5_7_4_1 <= FpAdd_8U_23U_qr_5_lpi_1_dfm_4_7_4_1;
      FpAdd_8U_23U_qr_5_lpi_1_dfm_5_3_0_1 <= FpAdd_8U_23U_qr_5_lpi_1_dfm_4_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_4_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
        & (mux_455_nl) ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_4_sva_st_3 <= MUX_s_1_2_2(alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_2_itm_7,
          FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_4_sva_st_2, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_4_sva_2 <= 6'b0;
      FpNormalize_8U_49U_if_or_3_itm_2 <= 1'b0;
    end
    else if ( IntLeadZero_49U_leading_sign_49_0_rtn_and_18_cse ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_4_sva_2 <= MUX_v_6_2_2(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_19,
          IntLeadZero_49U_leading_sign_49_0_rtn_4_sva, and_dcpl_241);
      FpNormalize_8U_49U_if_or_3_itm_2 <= MUX_s_1_2_2(FpNormalize_8U_49U_if_or_3_itm_mx0w0,
          FpNormalize_8U_49U_if_or_3_itm, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_4_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_461_nl) ) begin
      IsNaN_8U_23U_1_land_4_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_4_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_467_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_472_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_6_lpi_1_dfm_5_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_6_lpi_1_dfm_5_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_184_cse ) begin
      FpAdd_8U_23U_qr_6_lpi_1_dfm_5_7_4_1 <= FpAdd_8U_23U_qr_6_lpi_1_dfm_4_7_4_1;
      FpAdd_8U_23U_qr_6_lpi_1_dfm_5_3_0_1 <= FpAdd_8U_23U_qr_6_lpi_1_dfm_4_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_5_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
        & (mux_476_nl) ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_5_sva_st_3 <= MUX_s_1_2_2(alu_loop_op_5_FpAdd_8U_23U_if_3_if_acc_1_itm_7,
          FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_5_sva_st_2, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_5 <= 50'b0;
      alu_loop_op_5_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_int_mant_p1_and_20_cse ) begin
      FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_5 <= MUX_v_50_2_2(FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_mx1,
          FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm, and_dcpl_241);
      alu_loop_op_5_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 <= MUX_s_1_2_2((FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_mx2[49]),
          alu_loop_op_5_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_5_sva_2 <= 6'b0;
      FpNormalize_8U_49U_if_or_4_itm_2 <= 1'b0;
    end
    else if ( IntLeadZero_49U_leading_sign_49_0_rtn_and_19_cse ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_5_sva_2 <= MUX_v_6_2_2(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_20,
          IntLeadZero_49U_leading_sign_49_0_rtn_5_sva, and_dcpl_241);
      FpNormalize_8U_49U_if_or_4_itm_2 <= MUX_s_1_2_2(FpNormalize_8U_49U_if_or_4_itm_mx0w0,
          FpNormalize_8U_49U_if_or_4_itm, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_5_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_482_nl) ) begin
      IsNaN_8U_23U_1_land_5_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_5_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_488_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_5_lpi_1_dfm_st_5 <= 1'b0;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_5_sva_2 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_24_cse ) begin
      IsNaN_8U_23U_land_5_lpi_1_dfm_st_5 <= IsNaN_8U_23U_2_land_5_lpi_1_dfm_8;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_5_sva_2 <= alu_loop_op_5_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_493_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_7_lpi_1_dfm_5_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_7_lpi_1_dfm_5_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_186_cse ) begin
      FpAdd_8U_23U_qr_7_lpi_1_dfm_5_7_4_1 <= FpAdd_8U_23U_qr_7_lpi_1_dfm_4_7_4_1;
      FpAdd_8U_23U_qr_7_lpi_1_dfm_5_3_0_1 <= FpAdd_8U_23U_qr_7_lpi_1_dfm_4_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_6_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
        & (mux_497_nl) ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_6_sva_st_3 <= MUX_s_1_2_2(alu_loop_op_6_FpAdd_8U_23U_if_3_if_acc_2_itm_7,
          FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_6_sva_st_2, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_6_sva_2 <= 6'b0;
      FpNormalize_8U_49U_if_or_5_itm_2 <= 1'b0;
    end
    else if ( IntLeadZero_49U_leading_sign_49_0_rtn_and_20_cse ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_6_sva_2 <= MUX_v_6_2_2(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_21,
          IntLeadZero_49U_leading_sign_49_0_rtn_6_sva, and_dcpl_241);
      FpNormalize_8U_49U_if_or_5_itm_2 <= MUX_s_1_2_2(FpNormalize_8U_49U_if_or_5_itm_mx0w0,
          FpNormalize_8U_49U_if_or_5_itm, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_6_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_503_nl) ) begin
      IsNaN_8U_23U_1_land_6_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_6_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_509_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_514_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_8_lpi_1_dfm_5_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_8_lpi_1_dfm_5_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_188_cse ) begin
      FpAdd_8U_23U_qr_8_lpi_1_dfm_5_7_4_1 <= FpAdd_8U_23U_qr_8_lpi_1_dfm_4_7_4_1;
      FpAdd_8U_23U_qr_8_lpi_1_dfm_5_3_0_1 <= FpAdd_8U_23U_qr_8_lpi_1_dfm_4_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_7_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
        & (mux_518_nl) ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_7_sva_st_3 <= MUX_s_1_2_2(alu_loop_op_7_FpAdd_8U_23U_if_3_if_acc_1_itm_7,
          FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_7_sva_st_2, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_7_sva_2 <= 6'b0;
      FpNormalize_8U_49U_if_or_6_itm_2 <= 1'b0;
    end
    else if ( IntLeadZero_49U_leading_sign_49_0_rtn_and_21_cse ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_7_sva_2 <= MUX_v_6_2_2(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_22,
          IntLeadZero_49U_leading_sign_49_0_rtn_7_sva, and_dcpl_241);
      FpNormalize_8U_49U_if_or_6_itm_2 <= MUX_s_1_2_2(FpNormalize_8U_49U_if_or_6_itm_mx0w0,
          FpNormalize_8U_49U_if_or_6_itm, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_7_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_524_nl) ) begin
      IsNaN_8U_23U_1_land_7_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_7_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_530_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_535_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_9_lpi_1_dfm_5_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_9_lpi_1_dfm_5_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_190_cse ) begin
      FpAdd_8U_23U_qr_9_lpi_1_dfm_5_7_4_1 <= FpAdd_8U_23U_qr_9_lpi_1_dfm_4_7_4_1;
      FpAdd_8U_23U_qr_9_lpi_1_dfm_5_3_0_1 <= FpAdd_8U_23U_qr_9_lpi_1_dfm_4_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_8_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
        & (mux_539_nl) ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_8_sva_st_3 <= MUX_s_1_2_2(alu_loop_op_8_FpAdd_8U_23U_if_3_if_acc_2_itm_7,
          FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_8_sva_st_2, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_8_sva_2 <= 6'b0;
      FpNormalize_8U_49U_if_or_7_itm_2 <= 1'b0;
    end
    else if ( IntLeadZero_49U_leading_sign_49_0_rtn_and_22_cse ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_8_sva_2 <= MUX_v_6_2_2(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_23,
          IntLeadZero_49U_leading_sign_49_0_rtn_8_sva, and_dcpl_241);
      FpNormalize_8U_49U_if_or_7_itm_2 <= MUX_s_1_2_2(FpNormalize_8U_49U_if_or_7_itm_mx0w0,
          FpNormalize_8U_49U_if_or_7_itm, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_8_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_545_nl) ) begin
      IsNaN_8U_23U_1_land_8_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_8_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_551_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_556_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_10_lpi_1_dfm_5_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_10_lpi_1_dfm_5_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_192_cse ) begin
      FpAdd_8U_23U_qr_10_lpi_1_dfm_5_7_4_1 <= FpAdd_8U_23U_qr_10_lpi_1_dfm_4_7_4_1;
      FpAdd_8U_23U_qr_10_lpi_1_dfm_5_3_0_1 <= FpAdd_8U_23U_qr_10_lpi_1_dfm_4_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_9_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
        & (mux_560_nl) ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_9_sva_st_3 <= MUX_s_1_2_2(alu_loop_op_9_FpAdd_8U_23U_if_3_if_acc_1_itm_7,
          FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_9_sva_st_2, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_9_sva_2 <= 6'b0;
      FpNormalize_8U_49U_if_or_8_itm_2 <= 1'b0;
    end
    else if ( IntLeadZero_49U_leading_sign_49_0_rtn_and_23_cse ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_9_sva_2 <= MUX_v_6_2_2(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_24,
          IntLeadZero_49U_leading_sign_49_0_rtn_9_sva, and_dcpl_241);
      FpNormalize_8U_49U_if_or_8_itm_2 <= MUX_s_1_2_2(FpNormalize_8U_49U_if_or_8_itm_mx0w0,
          FpNormalize_8U_49U_if_or_8_itm, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_9_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_566_nl) ) begin
      IsNaN_8U_23U_1_land_9_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_9_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_572_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_577_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_11_lpi_1_dfm_5_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_11_lpi_1_dfm_5_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_194_cse ) begin
      FpAdd_8U_23U_qr_11_lpi_1_dfm_5_7_4_1 <= FpAdd_8U_23U_qr_11_lpi_1_dfm_4_7_4_1;
      FpAdd_8U_23U_qr_11_lpi_1_dfm_5_3_0_1 <= FpAdd_8U_23U_qr_11_lpi_1_dfm_4_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_10_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
        & (mux_581_nl) ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_10_sva_st_3 <= MUX_s_1_2_2(alu_loop_op_10_FpAdd_8U_23U_if_3_if_acc_2_itm_7,
          FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_10_sva_st_2,
          and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_10_sva_2 <= 6'b0;
      FpNormalize_8U_49U_if_or_9_itm_2 <= 1'b0;
    end
    else if ( IntLeadZero_49U_leading_sign_49_0_rtn_and_24_cse ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_10_sva_2 <= MUX_v_6_2_2(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_25,
          IntLeadZero_49U_leading_sign_49_0_rtn_10_sva, and_dcpl_241);
      FpNormalize_8U_49U_if_or_9_itm_2 <= MUX_s_1_2_2(FpNormalize_8U_49U_if_or_9_itm_mx0w0,
          FpNormalize_8U_49U_if_or_9_itm, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_10_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_587_nl) ) begin
      IsNaN_8U_23U_1_land_10_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_10_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_593_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_598_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_12_lpi_1_dfm_5_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_12_lpi_1_dfm_5_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_196_cse ) begin
      FpAdd_8U_23U_qr_12_lpi_1_dfm_5_7_4_1 <= FpAdd_8U_23U_qr_12_lpi_1_dfm_4_7_4_1;
      FpAdd_8U_23U_qr_12_lpi_1_dfm_5_3_0_1 <= FpAdd_8U_23U_qr_12_lpi_1_dfm_4_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_11_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
        & (mux_602_nl) ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_11_sva_st_3 <= MUX_s_1_2_2(alu_loop_op_11_FpAdd_8U_23U_if_3_if_acc_1_itm_7,
          FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_11_sva_st_2,
          and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_5 <= 50'b0;
      alu_loop_op_11_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_int_mant_p1_and_26_cse ) begin
      FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_5 <= MUX_v_50_2_2(FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_mx1,
          FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm, and_dcpl_241);
      alu_loop_op_11_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 <= MUX_s_1_2_2((FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_mx2[49]),
          alu_loop_op_11_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_11_sva_2 <= 6'b0;
      FpNormalize_8U_49U_if_or_10_itm_2 <= 1'b0;
    end
    else if ( IntLeadZero_49U_leading_sign_49_0_rtn_and_25_cse ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_11_sva_2 <= MUX_v_6_2_2(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_26,
          IntLeadZero_49U_leading_sign_49_0_rtn_11_sva, and_dcpl_241);
      FpNormalize_8U_49U_if_or_10_itm_2 <= MUX_s_1_2_2(FpNormalize_8U_49U_if_or_10_itm_mx0w0,
          FpNormalize_8U_49U_if_or_10_itm, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_11_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_608_nl) ) begin
      IsNaN_8U_23U_1_land_11_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_11_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_614_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_11_lpi_1_dfm_st_5 <= 1'b0;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_11_sva_2 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_36_cse ) begin
      IsNaN_8U_23U_land_11_lpi_1_dfm_st_5 <= IsNaN_8U_23U_2_land_11_lpi_1_dfm_8;
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_11_sva_2 <= alu_loop_op_11_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_619_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_13_lpi_1_dfm_5_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_13_lpi_1_dfm_5_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_198_cse ) begin
      FpAdd_8U_23U_qr_13_lpi_1_dfm_5_7_4_1 <= FpAdd_8U_23U_qr_13_lpi_1_dfm_4_7_4_1;
      FpAdd_8U_23U_qr_13_lpi_1_dfm_5_3_0_1 <= FpAdd_8U_23U_qr_13_lpi_1_dfm_4_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_12_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
        & (mux_623_nl) ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_12_sva_st_3 <= MUX_s_1_2_2(alu_loop_op_12_FpAdd_8U_23U_if_3_if_acc_2_itm_7,
          FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_12_sva_st_2,
          and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_12_sva_2 <= 6'b0;
      FpNormalize_8U_49U_if_or_11_itm_2 <= 1'b0;
    end
    else if ( IntLeadZero_49U_leading_sign_49_0_rtn_and_26_cse ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_12_sva_2 <= MUX_v_6_2_2(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_27,
          IntLeadZero_49U_leading_sign_49_0_rtn_12_sva, and_dcpl_241);
      FpNormalize_8U_49U_if_or_11_itm_2 <= MUX_s_1_2_2(FpNormalize_8U_49U_if_or_11_itm_mx0w0,
          FpNormalize_8U_49U_if_or_11_itm, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_12_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_629_nl) ) begin
      IsNaN_8U_23U_1_land_12_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_12_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_635_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_640_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_14_lpi_1_dfm_5_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_14_lpi_1_dfm_5_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_200_cse ) begin
      FpAdd_8U_23U_qr_14_lpi_1_dfm_5_7_4_1 <= FpAdd_8U_23U_qr_14_lpi_1_dfm_4_7_4_1;
      FpAdd_8U_23U_qr_14_lpi_1_dfm_5_3_0_1 <= FpAdd_8U_23U_qr_14_lpi_1_dfm_4_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_13_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
        & (mux_644_nl) ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_13_sva_st_3 <= MUX_s_1_2_2(alu_loop_op_13_FpAdd_8U_23U_if_3_if_acc_1_itm_7,
          FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_13_sva_st_2,
          and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_13_sva_2 <= 6'b0;
      FpNormalize_8U_49U_if_or_12_itm_2 <= 1'b0;
    end
    else if ( IntLeadZero_49U_leading_sign_49_0_rtn_and_27_cse ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_13_sva_2 <= MUX_v_6_2_2(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_28,
          IntLeadZero_49U_leading_sign_49_0_rtn_13_sva, and_dcpl_241);
      FpNormalize_8U_49U_if_or_12_itm_2 <= MUX_s_1_2_2(FpNormalize_8U_49U_if_or_12_itm_mx0w0,
          FpNormalize_8U_49U_if_or_12_itm, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_13_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_650_nl) ) begin
      IsNaN_8U_23U_1_land_13_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_13_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_656_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_661_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_15_lpi_1_dfm_5_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_15_lpi_1_dfm_5_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_202_cse ) begin
      FpAdd_8U_23U_qr_15_lpi_1_dfm_5_7_4_1 <= FpAdd_8U_23U_qr_15_lpi_1_dfm_4_7_4_1;
      FpAdd_8U_23U_qr_15_lpi_1_dfm_5_3_0_1 <= FpAdd_8U_23U_qr_15_lpi_1_dfm_4_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_14_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
        & (mux_665_nl) ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_14_sva_st_3 <= MUX_s_1_2_2(alu_loop_op_14_FpAdd_8U_23U_if_3_if_acc_2_itm_7,
          FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_14_sva_st_2,
          and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_14_sva_2 <= 6'b0;
      FpNormalize_8U_49U_if_or_13_itm_2 <= 1'b0;
    end
    else if ( IntLeadZero_49U_leading_sign_49_0_rtn_and_28_cse ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_14_sva_2 <= MUX_v_6_2_2(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_29,
          IntLeadZero_49U_leading_sign_49_0_rtn_14_sva, and_dcpl_241);
      FpNormalize_8U_49U_if_or_13_itm_2 <= MUX_s_1_2_2(FpNormalize_8U_49U_if_or_13_itm_mx0w0,
          FpNormalize_8U_49U_if_or_13_itm, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_14_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_671_nl) ) begin
      IsNaN_8U_23U_1_land_14_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_14_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_677_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_681_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_16_lpi_1_dfm_5_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_16_lpi_1_dfm_5_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_204_cse ) begin
      FpAdd_8U_23U_qr_16_lpi_1_dfm_5_7_4_1 <= FpAdd_8U_23U_qr_16_lpi_1_dfm_4_7_4_1;
      FpAdd_8U_23U_qr_16_lpi_1_dfm_5_3_0_1 <= FpAdd_8U_23U_qr_16_lpi_1_dfm_4_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_15_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
        & (mux_685_nl) ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_15_sva_st_3 <= MUX_s_1_2_2(alu_loop_op_15_FpAdd_8U_23U_if_3_if_acc_1_itm_7,
          FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_15_sva_st_2,
          and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_15_sva_2 <= 6'b0;
      FpNormalize_8U_49U_if_or_14_itm_2 <= 1'b0;
    end
    else if ( IntLeadZero_49U_leading_sign_49_0_rtn_and_29_cse ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_15_sva_2 <= MUX_v_6_2_2(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_30,
          IntLeadZero_49U_leading_sign_49_0_rtn_15_sva, and_dcpl_241);
      FpNormalize_8U_49U_if_or_14_itm_2 <= MUX_s_1_2_2(FpNormalize_8U_49U_if_or_14_itm_mx0w0,
          FpNormalize_8U_49U_if_or_14_itm, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_15_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_691_nl) ) begin
      IsNaN_8U_23U_1_land_15_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_15_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_697_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_701_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_lpi_1_dfm_5_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_lpi_1_dfm_5_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_206_cse ) begin
      FpAdd_8U_23U_qr_lpi_1_dfm_5_7_4_1 <= FpAdd_8U_23U_qr_lpi_1_dfm_4_7_4_1;
      FpAdd_8U_23U_qr_lpi_1_dfm_5_3_0_1 <= FpAdd_8U_23U_qr_lpi_1_dfm_4_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_b_left_shift_FpAdd_8U_23U_b_left_shift_or_31_cse
        & (mux_705_nl) ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_st_3 <= MUX_s_1_2_2(alu_loop_op_16_FpAdd_8U_23U_if_3_if_acc_2_itm_7,
          FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_st_2, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_sva_2 <= 6'b0;
      FpNormalize_8U_49U_if_or_15_itm_2 <= 1'b0;
    end
    else if ( IntLeadZero_49U_leading_sign_49_0_rtn_and_30_cse ) begin
      IntLeadZero_49U_leading_sign_49_0_rtn_sva_2 <= MUX_v_6_2_2(libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_31,
          IntLeadZero_49U_leading_sign_49_0_rtn_sva, and_dcpl_241);
      FpNormalize_8U_49U_if_or_15_itm_2 <= MUX_s_1_2_2(FpNormalize_8U_49U_if_or_15_itm_mx0w0,
          FpNormalize_8U_49U_if_or_15_itm, and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_711_nl) ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_717_nl) ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_11 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_or_861_itm_4 <= 1'b0;
      reg_FpAlu_8U_23U_or_797_cse <= 1'b0;
      FpAlu_8U_23U_or_859_itm_4 <= 1'b0;
      reg_FpAlu_8U_23U_or_794_cse <= 1'b0;
      FpAlu_8U_23U_or_857_itm_4 <= 1'b0;
      reg_FpAlu_8U_23U_or_791_cse <= 1'b0;
      FpAlu_8U_23U_or_855_itm_4 <= 1'b0;
      reg_FpAlu_8U_23U_or_788_cse <= 1'b0;
      FpAlu_8U_23U_or_853_itm_4 <= 1'b0;
      reg_FpAlu_8U_23U_or_785_cse <= 1'b0;
      FpAlu_8U_23U_or_849_itm_4 <= 1'b0;
      reg_FpAlu_8U_23U_or_779_cse <= 1'b0;
      FpAlu_8U_23U_or_847_itm_4 <= 1'b0;
      reg_FpAlu_8U_23U_or_776_cse <= 1'b0;
      FpAlu_8U_23U_or_845_itm_4 <= 1'b0;
      reg_FpAlu_8U_23U_or_773_cse <= 1'b0;
      FpAlu_8U_23U_or_843_itm_4 <= 1'b0;
      reg_FpAlu_8U_23U_or_770_cse <= 1'b0;
      FpAlu_8U_23U_or_841_itm_4 <= 1'b0;
      reg_FpAlu_8U_23U_or_767_cse <= 1'b0;
      FpAlu_8U_23U_or_837_itm_4 <= 1'b0;
      reg_FpAlu_8U_23U_or_761_cse <= 1'b0;
      FpAlu_8U_23U_or_835_itm_4 <= 1'b0;
      reg_FpAlu_8U_23U_or_758_cse <= 1'b0;
      FpAlu_8U_23U_or_833_itm_4 <= 1'b0;
      reg_FpAlu_8U_23U_or_755_cse <= 1'b0;
      FpAlu_8U_23U_or_831_itm_4 <= 1'b0;
      reg_FpAlu_8U_23U_or_752_cse <= 1'b0;
    end
    else if ( FpAlu_8U_23U_and_849_cse ) begin
      FpAlu_8U_23U_or_861_itm_4 <= FpAlu_8U_23U_or_861_itm_3;
      reg_FpAlu_8U_23U_or_797_cse <= FpAlu_8U_23U_or_797_itm_3;
      FpAlu_8U_23U_or_859_itm_4 <= FpAlu_8U_23U_or_859_itm_3;
      reg_FpAlu_8U_23U_or_794_cse <= FpAlu_8U_23U_or_794_itm_3;
      FpAlu_8U_23U_or_857_itm_4 <= FpAlu_8U_23U_or_857_itm_3;
      reg_FpAlu_8U_23U_or_791_cse <= FpAlu_8U_23U_or_791_itm_3;
      FpAlu_8U_23U_or_855_itm_4 <= FpAlu_8U_23U_or_855_itm_3;
      reg_FpAlu_8U_23U_or_788_cse <= FpAlu_8U_23U_or_788_itm_3;
      FpAlu_8U_23U_or_853_itm_4 <= FpAlu_8U_23U_or_853_itm_3;
      reg_FpAlu_8U_23U_or_785_cse <= FpAlu_8U_23U_or_785_itm_3;
      FpAlu_8U_23U_or_849_itm_4 <= FpAlu_8U_23U_or_849_itm_3;
      reg_FpAlu_8U_23U_or_779_cse <= FpAlu_8U_23U_or_779_itm_3;
      FpAlu_8U_23U_or_847_itm_4 <= FpAlu_8U_23U_or_847_itm_3;
      reg_FpAlu_8U_23U_or_776_cse <= FpAlu_8U_23U_or_776_itm_3;
      FpAlu_8U_23U_or_845_itm_4 <= FpAlu_8U_23U_or_845_itm_3;
      reg_FpAlu_8U_23U_or_773_cse <= FpAlu_8U_23U_or_773_itm_3;
      FpAlu_8U_23U_or_843_itm_4 <= FpAlu_8U_23U_or_843_itm_3;
      reg_FpAlu_8U_23U_or_770_cse <= FpAlu_8U_23U_or_770_itm_3;
      FpAlu_8U_23U_or_841_itm_4 <= FpAlu_8U_23U_or_841_itm_3;
      reg_FpAlu_8U_23U_or_767_cse <= FpAlu_8U_23U_or_767_itm_3;
      FpAlu_8U_23U_or_837_itm_4 <= FpAlu_8U_23U_or_837_itm_3;
      reg_FpAlu_8U_23U_or_761_cse <= FpAlu_8U_23U_or_761_itm_3;
      FpAlu_8U_23U_or_835_itm_4 <= FpAlu_8U_23U_or_835_itm_3;
      reg_FpAlu_8U_23U_or_758_cse <= FpAlu_8U_23U_or_758_itm_3;
      FpAlu_8U_23U_or_833_itm_4 <= FpAlu_8U_23U_or_833_itm_3;
      reg_FpAlu_8U_23U_or_755_cse <= FpAlu_8U_23U_or_755_itm_3;
      FpAlu_8U_23U_or_831_itm_4 <= FpAlu_8U_23U_or_831_itm_3;
      reg_FpAlu_8U_23U_or_752_cse <= FpAlu_8U_23U_or_752_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_algo_1_sva_st_205 <= 2'b0;
      cfg_alu_algo_1_sva_7 <= 2'b0;
    end
    else if ( cfg_alu_algo_and_115_cse ) begin
      cfg_alu_algo_1_sva_st_205 <= cfg_alu_algo_1_sva_st_204;
      cfg_alu_algo_1_sva_7 <= cfg_alu_algo_1_sva_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_or_851_itm_4 <= 1'b0;
      reg_FpAlu_8U_23U_or_782_cse <= 1'b0;
      FpAlu_8U_23U_or_839_itm_4 <= 1'b0;
      reg_FpAlu_8U_23U_or_764_cse <= 1'b0;
    end
    else if ( FpAlu_8U_23U_and_889_cse ) begin
      FpAlu_8U_23U_or_851_itm_4 <= FpAlu_8U_23U_or_851_itm_3;
      reg_FpAlu_8U_23U_or_782_cse <= FpAlu_8U_23U_or_782_itm_3;
      FpAlu_8U_23U_or_839_itm_4 <= FpAlu_8U_23U_or_839_itm_3;
      reg_FpAlu_8U_23U_or_764_cse <= FpAlu_8U_23U_or_764_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_1 <= 1'b0;
    end
    else if ( core_wen & (or_tmp_3044 | main_stage_v_1_mx0c1) ) begin
      main_stage_v_1 <= ~ main_stage_v_1_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      AluIn_data_sva_1 <= 512'b0;
      io_read_cfg_alu_bypass_rsc_svs_st_1 <= 1'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_15_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_14_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_13_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_12_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_11_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_10_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_9_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_8_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_7_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_6_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_5_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_4_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_4 <= 1'b0;
      alu_loop_op_else_nor_tmp_16 <= 1'b0;
    end
    else if ( AluIn_data_and_cse ) begin
      AluIn_data_sva_1 <= chn_alu_in_rsci_d_mxwt;
      io_read_cfg_alu_bypass_rsc_svs_st_1 <= cfg_alu_bypass_rsci_d;
      IsNaN_8U_23U_land_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_land_15_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_15_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_land_14_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_14_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_land_13_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_13_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_land_12_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_12_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_land_11_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_11_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_land_10_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_10_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_land_9_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_9_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_land_8_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_8_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_land_7_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_7_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_land_6_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_6_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_land_5_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_5_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_land_4_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_4_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_3_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_2_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_1_lpi_1_dfm_mx1w0;
      alu_loop_op_else_nor_tmp_16 <= cfg_alu_algo_rsci_d[1];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_2_land_1_lpi_1_dfm_st_1 <= 1'b0;
      IsNaN_8U_23U_2_land_2_lpi_1_dfm_st_1 <= 1'b0;
      IsNaN_8U_23U_2_land_3_lpi_1_dfm_st_1 <= 1'b0;
      IsNaN_8U_23U_2_land_4_lpi_1_dfm_st_1 <= 1'b0;
      IsNaN_8U_23U_2_land_5_lpi_1_dfm_st_1 <= 1'b0;
      IsNaN_8U_23U_2_land_6_lpi_1_dfm_st_1 <= 1'b0;
      IsNaN_8U_23U_2_land_7_lpi_1_dfm_st_1 <= 1'b0;
      IsNaN_8U_23U_2_land_8_lpi_1_dfm_st_1 <= 1'b0;
      IsNaN_8U_23U_2_land_9_lpi_1_dfm_st_1 <= 1'b0;
      IsNaN_8U_23U_2_land_10_lpi_1_dfm_st_1 <= 1'b0;
      IsNaN_8U_23U_2_land_11_lpi_1_dfm_st_1 <= 1'b0;
      IsNaN_8U_23U_2_land_12_lpi_1_dfm_st_1 <= 1'b0;
      IsNaN_8U_23U_2_land_13_lpi_1_dfm_st_1 <= 1'b0;
      IsNaN_8U_23U_2_land_14_lpi_1_dfm_st_1 <= 1'b0;
      IsNaN_8U_23U_2_land_15_lpi_1_dfm_st_1 <= 1'b0;
      IsNaN_8U_23U_2_land_lpi_1_dfm_st_1 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_2_aelse_and_48_cse ) begin
      IsNaN_8U_23U_2_land_1_lpi_1_dfm_st_1 <= MUX_s_1_2_2(IsNaN_8U_23U_2_land_1_lpi_1_dfm_mx1w0,
          IsNaN_8U_23U_2_land_1_lpi_1_dfm_st, and_dcpl_395);
      IsNaN_8U_23U_2_land_2_lpi_1_dfm_st_1 <= MUX_s_1_2_2(IsNaN_8U_23U_2_land_2_lpi_1_dfm_mx1w0,
          IsNaN_8U_23U_2_land_2_lpi_1_dfm_st, and_dcpl_395);
      IsNaN_8U_23U_2_land_3_lpi_1_dfm_st_1 <= MUX_s_1_2_2(IsNaN_8U_23U_2_land_3_lpi_1_dfm_mx1w0,
          IsNaN_8U_23U_2_land_3_lpi_1_dfm_st, and_dcpl_395);
      IsNaN_8U_23U_2_land_4_lpi_1_dfm_st_1 <= MUX_s_1_2_2(IsNaN_8U_23U_2_land_4_lpi_1_dfm_mx1w0,
          IsNaN_8U_23U_2_land_4_lpi_1_dfm_st, and_dcpl_395);
      IsNaN_8U_23U_2_land_5_lpi_1_dfm_st_1 <= MUX_s_1_2_2(IsNaN_8U_23U_2_land_5_lpi_1_dfm_mx1w0,
          IsNaN_8U_23U_2_land_5_lpi_1_dfm_st, and_dcpl_395);
      IsNaN_8U_23U_2_land_6_lpi_1_dfm_st_1 <= MUX_s_1_2_2(IsNaN_8U_23U_2_land_6_lpi_1_dfm_mx1w0,
          IsNaN_8U_23U_2_land_6_lpi_1_dfm_st, and_dcpl_395);
      IsNaN_8U_23U_2_land_7_lpi_1_dfm_st_1 <= MUX_s_1_2_2(IsNaN_8U_23U_2_land_7_lpi_1_dfm_mx1w0,
          IsNaN_8U_23U_2_land_7_lpi_1_dfm_st, and_dcpl_395);
      IsNaN_8U_23U_2_land_8_lpi_1_dfm_st_1 <= MUX_s_1_2_2(IsNaN_8U_23U_2_land_8_lpi_1_dfm_mx1w0,
          IsNaN_8U_23U_2_land_8_lpi_1_dfm_st, and_dcpl_395);
      IsNaN_8U_23U_2_land_9_lpi_1_dfm_st_1 <= MUX_s_1_2_2(IsNaN_8U_23U_2_land_9_lpi_1_dfm_mx1w0,
          IsNaN_8U_23U_2_land_9_lpi_1_dfm_st, and_dcpl_395);
      IsNaN_8U_23U_2_land_10_lpi_1_dfm_st_1 <= MUX_s_1_2_2(IsNaN_8U_23U_2_land_10_lpi_1_dfm_mx1w0,
          IsNaN_8U_23U_2_land_10_lpi_1_dfm_st, and_dcpl_395);
      IsNaN_8U_23U_2_land_11_lpi_1_dfm_st_1 <= MUX_s_1_2_2(IsNaN_8U_23U_2_land_11_lpi_1_dfm_mx1w0,
          IsNaN_8U_23U_2_land_11_lpi_1_dfm_st, and_dcpl_395);
      IsNaN_8U_23U_2_land_12_lpi_1_dfm_st_1 <= MUX_s_1_2_2(IsNaN_8U_23U_2_land_12_lpi_1_dfm_mx1w0,
          IsNaN_8U_23U_2_land_12_lpi_1_dfm_st, and_dcpl_395);
      IsNaN_8U_23U_2_land_13_lpi_1_dfm_st_1 <= MUX_s_1_2_2(IsNaN_8U_23U_2_land_13_lpi_1_dfm_mx1w0,
          IsNaN_8U_23U_2_land_13_lpi_1_dfm_st, and_dcpl_395);
      IsNaN_8U_23U_2_land_14_lpi_1_dfm_st_1 <= MUX_s_1_2_2(IsNaN_8U_23U_2_land_14_lpi_1_dfm_mx1w0,
          IsNaN_8U_23U_2_land_14_lpi_1_dfm_st, and_dcpl_395);
      IsNaN_8U_23U_2_land_15_lpi_1_dfm_st_1 <= MUX_s_1_2_2(IsNaN_8U_23U_2_land_15_lpi_1_dfm_mx1w0,
          IsNaN_8U_23U_2_land_15_lpi_1_dfm_st, and_dcpl_395);
      IsNaN_8U_23U_2_land_lpi_1_dfm_st_1 <= MUX_s_1_2_2(IsNaN_8U_23U_2_land_lpi_1_dfm_mx1w0,
          IsNaN_8U_23U_2_land_lpi_1_dfm_st, and_dcpl_395);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_algo_1_sva_st_92 <= 2'b0;
      cfg_alu_algo_1_sva_st_96 <= 2'b0;
    end
    else if ( cfg_alu_algo_and_132_cse ) begin
      cfg_alu_algo_1_sva_st_92 <= MUX_v_2_2_2(cfg_alu_algo_rsci_d, cfg_alu_algo_1_sva_st_15,
          and_dcpl_395);
      cfg_alu_algo_1_sva_st_96 <= MUX_v_2_2_2(cfg_alu_algo_rsci_d, cfg_alu_algo_1_sva_st_31,
          and_dcpl_394);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_op_1_sva_1 <= 16'b0;
    end
    else if ( IsNaN_8U_23U_2_aelse_and_cse & and_91_tmp & (~(cfg_alu_src_rsci_d |
        cfg_alu_bypass_rsci_d)) ) begin
      cfg_alu_op_1_sva_1 <= cfg_alu_op_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_src_1_sva_st_1 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_11 & (fsm_output[1])) | cfg_alu_src_1_sva_st_1_mx0c1)
        ) begin
      cfg_alu_src_1_sva_st_1 <= MUX_s_1_2_2(cfg_alu_src_rsci_d, cfg_alu_src_1_sva_st,
          cfg_alu_src_1_sva_st_1_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_2_lpi_1_dfm_4_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_2_lpi_1_dfm_4_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_208_cse ) begin
      FpAdd_8U_23U_qr_2_lpi_1_dfm_4_7_4_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[30:27]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_9, FpAdd_8U_23U_qr_2_lpi_1_dfm_7_4,
          {and_dcpl_402 , and_dcpl_407 , and_dcpl_408});
      FpAdd_8U_23U_qr_2_lpi_1_dfm_4_3_0_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[26:23]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_9, FpAdd_8U_23U_qr_2_lpi_1_dfm_3_0,
          {and_dcpl_402 , and_dcpl_407 , and_dcpl_408});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_137) & mux_tmp_778 ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_st_2 <= alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_itm <= 1'b0;
      IntLeadZero_49U_leading_sign_49_0_rtn_1_sva <= 6'b0;
    end
    else if ( FpNormalize_8U_49U_if_and_31_cse ) begin
      FpNormalize_8U_49U_if_or_itm <= FpNormalize_8U_49U_if_or_itm_mx0w0;
      IntLeadZero_49U_leading_sign_49_0_rtn_1_sva <= libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_16;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_lpi_1_dfm <= 50'b0;
    end
    else if ( FpAdd_8U_23U_int_mant_p1_and_cse ) begin
      FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm <= FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_mx1;
      FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm <= FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_mx1;
      FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm <= FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_mx1;
      FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm <= FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_mx1;
      FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm <= FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_mx1;
      FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm <= FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_mx1;
      FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm <= FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_mx1;
      FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm <= FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_mx1;
      FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm <= FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_mx1;
      FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm <= FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_mx1;
      FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm <= FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_mx1;
      FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm <= FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_mx1;
      FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm <= FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_mx1;
      FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm <= FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_mx1;
      FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm <= FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_mx1;
      FpAdd_8U_23U_int_mant_p1_lpi_1_dfm <= FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_mx1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm <= 1'b0;
      alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm <= 1'b0;
      alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm <= 1'b0;
      alu_loop_op_5_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm <= 1'b0;
      alu_loop_op_6_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm <= 1'b0;
      alu_loop_op_7_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm <= 1'b0;
      alu_loop_op_8_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm <= 1'b0;
      alu_loop_op_9_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm <= 1'b0;
      alu_loop_op_10_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm <= 1'b0;
      alu_loop_op_11_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm <= 1'b0;
      alu_loop_op_12_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm <= 1'b0;
      alu_loop_op_13_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm <= 1'b0;
      alu_loop_op_14_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm <= 1'b0;
      alu_loop_op_15_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm <= 1'b0;
      alu_loop_op_16_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm <= 1'b0;
    end
    else if ( FpAdd_8U_23U_if_3_and_cse ) begin
      alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm <= FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_mx2[49];
      alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm <= FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_mx2[49];
      alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm <= FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_mx2[49];
      alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm <= FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_mx2[49];
      alu_loop_op_5_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm <= FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_mx2[49];
      alu_loop_op_6_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm <= FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_mx2[49];
      alu_loop_op_7_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm <= FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_mx2[49];
      alu_loop_op_8_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm <= FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_mx2[49];
      alu_loop_op_9_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm <= FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_mx2[49];
      alu_loop_op_10_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm <= FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_mx2[49];
      alu_loop_op_11_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm <= FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_mx2[49];
      alu_loop_op_12_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm <= FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_mx2[49];
      alu_loop_op_13_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm <= FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_mx2[49];
      alu_loop_op_14_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm <= FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_mx2[49];
      alu_loop_op_15_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm <= FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_mx2[49];
      alu_loop_op_16_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm <= FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_mx2[49];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_3_lpi_1_dfm_4_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_3_lpi_1_dfm_4_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_210_cse ) begin
      FpAdd_8U_23U_qr_3_lpi_1_dfm_4_7_4_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[62:59]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_9, FpAdd_8U_23U_qr_3_lpi_1_dfm_7_4,
          {and_dcpl_417 , and_dcpl_422 , and_dcpl_408});
      FpAdd_8U_23U_qr_3_lpi_1_dfm_4_3_0_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[58:55]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_9, FpAdd_8U_23U_qr_3_lpi_1_dfm_3_0,
          {and_dcpl_417 , and_dcpl_422 , and_dcpl_408});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_137) & mux_tmp_779 ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_st_2 <= alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_1_itm <= 1'b0;
      IntLeadZero_49U_leading_sign_49_0_rtn_2_sva <= 6'b0;
    end
    else if ( FpNormalize_8U_49U_if_and_32_cse ) begin
      FpNormalize_8U_49U_if_or_1_itm <= FpNormalize_8U_49U_if_or_1_itm_mx0w0;
      IntLeadZero_49U_leading_sign_49_0_rtn_2_sva <= libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_17;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_4_lpi_1_dfm_4_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_4_lpi_1_dfm_4_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_212_cse ) begin
      FpAdd_8U_23U_qr_4_lpi_1_dfm_4_7_4_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[94:91]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_9, FpAdd_8U_23U_qr_4_lpi_1_dfm_7_4,
          {and_dcpl_432 , and_dcpl_437 , and_dcpl_408});
      FpAdd_8U_23U_qr_4_lpi_1_dfm_4_3_0_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[90:87]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_9, FpAdd_8U_23U_qr_4_lpi_1_dfm_3_0,
          {and_dcpl_432 , and_dcpl_437 , and_dcpl_408});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_137) & mux_tmp_781 ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_st_2 <= alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_2_itm <= 1'b0;
      IntLeadZero_49U_leading_sign_49_0_rtn_3_sva <= 6'b0;
    end
    else if ( FpNormalize_8U_49U_if_and_33_cse ) begin
      FpNormalize_8U_49U_if_or_2_itm <= FpNormalize_8U_49U_if_or_2_itm_mx0w0;
      IntLeadZero_49U_leading_sign_49_0_rtn_3_sva <= libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_18;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_5_lpi_1_dfm_4_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_5_lpi_1_dfm_4_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_214_cse ) begin
      FpAdd_8U_23U_qr_5_lpi_1_dfm_4_7_4_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[126:123]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_9, FpAdd_8U_23U_qr_5_lpi_1_dfm_7_4,
          {and_dcpl_447 , and_dcpl_452 , and_dcpl_408});
      FpAdd_8U_23U_qr_5_lpi_1_dfm_4_3_0_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[122:119]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_9, FpAdd_8U_23U_qr_5_lpi_1_dfm_3_0,
          {and_dcpl_447 , and_dcpl_452 , and_dcpl_408});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_4_sva_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_137) & mux_tmp_782 ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_4_sva_st_2 <= alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_3_itm <= 1'b0;
      IntLeadZero_49U_leading_sign_49_0_rtn_4_sva <= 6'b0;
    end
    else if ( FpNormalize_8U_49U_if_and_34_cse ) begin
      FpNormalize_8U_49U_if_or_3_itm <= FpNormalize_8U_49U_if_or_3_itm_mx0w0;
      IntLeadZero_49U_leading_sign_49_0_rtn_4_sva <= libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_19;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_5_sva_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_137) & mux_tmp_783 ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_5_sva_st_2 <= alu_loop_op_5_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_4_itm <= 1'b0;
      IntLeadZero_49U_leading_sign_49_0_rtn_5_sva <= 6'b0;
    end
    else if ( FpNormalize_8U_49U_if_and_35_cse ) begin
      FpNormalize_8U_49U_if_or_4_itm <= FpNormalize_8U_49U_if_or_4_itm_mx0w0;
      IntLeadZero_49U_leading_sign_49_0_rtn_5_sva <= libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_20;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_6_sva_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_137) & mux_tmp_785 ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_6_sva_st_2 <= alu_loop_op_6_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_5_itm <= 1'b0;
      IntLeadZero_49U_leading_sign_49_0_rtn_6_sva <= 6'b0;
    end
    else if ( FpNormalize_8U_49U_if_and_36_cse ) begin
      FpNormalize_8U_49U_if_or_5_itm <= FpNormalize_8U_49U_if_or_5_itm_mx0w0;
      IntLeadZero_49U_leading_sign_49_0_rtn_6_sva <= libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_21;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_7_sva_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_137) & mux_tmp_786 ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_7_sva_st_2 <= alu_loop_op_7_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_6_itm <= 1'b0;
      IntLeadZero_49U_leading_sign_49_0_rtn_7_sva <= 6'b0;
    end
    else if ( FpNormalize_8U_49U_if_and_37_cse ) begin
      FpNormalize_8U_49U_if_or_6_itm <= FpNormalize_8U_49U_if_or_6_itm_mx0w0;
      IntLeadZero_49U_leading_sign_49_0_rtn_7_sva <= libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_22;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_9_lpi_1_dfm_4_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_9_lpi_1_dfm_4_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_216_cse ) begin
      FpAdd_8U_23U_qr_9_lpi_1_dfm_4_7_4_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[254:251]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_9, FpAdd_8U_23U_qr_9_lpi_1_dfm_7_4,
          {and_dcpl_474 , and_dcpl_479 , and_dcpl_408});
      FpAdd_8U_23U_qr_9_lpi_1_dfm_4_3_0_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[250:247]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_9, FpAdd_8U_23U_qr_9_lpi_1_dfm_3_0,
          {and_dcpl_474 , and_dcpl_479 , and_dcpl_408});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_8_sva_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_137) & mux_tmp_787 ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_8_sva_st_2 <= alu_loop_op_8_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_7_itm <= 1'b0;
      IntLeadZero_49U_leading_sign_49_0_rtn_8_sva <= 6'b0;
    end
    else if ( FpNormalize_8U_49U_if_and_38_cse ) begin
      FpNormalize_8U_49U_if_or_7_itm <= FpNormalize_8U_49U_if_or_7_itm_mx0w0;
      IntLeadZero_49U_leading_sign_49_0_rtn_8_sva <= libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_23;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_9_sva_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_137) & mux_tmp_788 ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_9_sva_st_2 <= alu_loop_op_9_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_8_itm <= 1'b0;
      IntLeadZero_49U_leading_sign_49_0_rtn_9_sva <= 6'b0;
    end
    else if ( FpNormalize_8U_49U_if_and_39_cse ) begin
      FpNormalize_8U_49U_if_or_8_itm <= FpNormalize_8U_49U_if_or_8_itm_mx0w0;
      IntLeadZero_49U_leading_sign_49_0_rtn_9_sva <= libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_24;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_10_sva_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_137) & mux_tmp_789 ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_10_sva_st_2 <= alu_loop_op_10_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_9_itm <= 1'b0;
      IntLeadZero_49U_leading_sign_49_0_rtn_10_sva <= 6'b0;
    end
    else if ( FpNormalize_8U_49U_if_and_40_cse ) begin
      FpNormalize_8U_49U_if_or_9_itm <= FpNormalize_8U_49U_if_or_9_itm_mx0w0;
      IntLeadZero_49U_leading_sign_49_0_rtn_10_sva <= libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_25;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_11_sva_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_137) & mux_tmp_790 ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_11_sva_st_2 <= alu_loop_op_11_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_10_itm <= 1'b0;
      IntLeadZero_49U_leading_sign_49_0_rtn_11_sva <= 6'b0;
    end
    else if ( FpNormalize_8U_49U_if_and_41_cse ) begin
      FpNormalize_8U_49U_if_or_10_itm <= FpNormalize_8U_49U_if_or_10_itm_mx0w0;
      IntLeadZero_49U_leading_sign_49_0_rtn_11_sva <= libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_26;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_12_sva_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_137) & mux_tmp_791 ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_12_sva_st_2 <= alu_loop_op_12_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_11_itm <= 1'b0;
      IntLeadZero_49U_leading_sign_49_0_rtn_12_sva <= 6'b0;
    end
    else if ( FpNormalize_8U_49U_if_and_42_cse ) begin
      FpNormalize_8U_49U_if_or_11_itm <= FpNormalize_8U_49U_if_or_11_itm_mx0w0;
      IntLeadZero_49U_leading_sign_49_0_rtn_12_sva <= libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_27;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_14_lpi_1_dfm_4_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_14_lpi_1_dfm_4_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_218_cse ) begin
      FpAdd_8U_23U_qr_14_lpi_1_dfm_4_7_4_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[414:411]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_9, FpAdd_8U_23U_qr_14_lpi_1_dfm_7_4,
          {and_dcpl_505 , and_dcpl_510 , and_dcpl_408});
      FpAdd_8U_23U_qr_14_lpi_1_dfm_4_3_0_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[410:407]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_9, FpAdd_8U_23U_qr_14_lpi_1_dfm_3_0,
          {and_dcpl_505 , and_dcpl_510 , and_dcpl_408});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_13_sva_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_137) & mux_tmp_792 ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_13_sva_st_2 <= alu_loop_op_13_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_12_itm <= 1'b0;
      IntLeadZero_49U_leading_sign_49_0_rtn_13_sva <= 6'b0;
    end
    else if ( FpNormalize_8U_49U_if_and_43_cse ) begin
      FpNormalize_8U_49U_if_or_12_itm <= FpNormalize_8U_49U_if_or_12_itm_mx0w0;
      IntLeadZero_49U_leading_sign_49_0_rtn_13_sva <= libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_28;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_15_lpi_1_dfm_4_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_15_lpi_1_dfm_4_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_220_cse ) begin
      FpAdd_8U_23U_qr_15_lpi_1_dfm_4_7_4_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[446:443]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_9, FpAdd_8U_23U_qr_15_lpi_1_dfm_7_4,
          {and_dcpl_520 , and_dcpl_525 , and_dcpl_408});
      FpAdd_8U_23U_qr_15_lpi_1_dfm_4_3_0_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[442:439]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_9, FpAdd_8U_23U_qr_15_lpi_1_dfm_3_0,
          {and_dcpl_520 , and_dcpl_525 , and_dcpl_408});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_14_sva_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_137) & mux_tmp_793 ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_14_sva_st_2 <= alu_loop_op_14_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_13_itm <= 1'b0;
      IntLeadZero_49U_leading_sign_49_0_rtn_14_sva <= 6'b0;
    end
    else if ( FpNormalize_8U_49U_if_and_44_cse ) begin
      FpNormalize_8U_49U_if_or_13_itm <= FpNormalize_8U_49U_if_or_13_itm_mx0w0;
      IntLeadZero_49U_leading_sign_49_0_rtn_14_sva <= libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_29;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_16_lpi_1_dfm_4_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_16_lpi_1_dfm_4_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_222_cse ) begin
      FpAdd_8U_23U_qr_16_lpi_1_dfm_4_7_4_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[478:475]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_9, FpAdd_8U_23U_qr_16_lpi_1_dfm_7_4,
          {and_dcpl_535 , and_dcpl_540 , and_dcpl_408});
      FpAdd_8U_23U_qr_16_lpi_1_dfm_4_3_0_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[474:471]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_9, FpAdd_8U_23U_qr_16_lpi_1_dfm_3_0,
          {and_dcpl_535 , and_dcpl_540 , and_dcpl_408});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_15_sva_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_137) & mux_tmp_795 ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_15_sva_st_2 <= alu_loop_op_15_FpAdd_8U_23U_if_3_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_14_itm <= 1'b0;
      IntLeadZero_49U_leading_sign_49_0_rtn_15_sva <= 6'b0;
    end
    else if ( FpNormalize_8U_49U_if_and_45_cse ) begin
      FpNormalize_8U_49U_if_or_14_itm <= FpNormalize_8U_49U_if_or_14_itm_mx0w0;
      IntLeadZero_49U_leading_sign_49_0_rtn_15_sva <= libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_30;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_lpi_1_dfm_4_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_lpi_1_dfm_4_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_224_cse ) begin
      FpAdd_8U_23U_qr_lpi_1_dfm_4_7_4_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[510:507]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_9, FpAdd_8U_23U_qr_lpi_1_dfm_7_4,
          {and_dcpl_550 , and_dcpl_555 , and_dcpl_408});
      FpAdd_8U_23U_qr_lpi_1_dfm_4_3_0_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[506:503]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_9, FpAdd_8U_23U_qr_lpi_1_dfm_3_0,
          {and_dcpl_550 , and_dcpl_555 , and_dcpl_408});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_137) & mux_tmp_796 ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_st_2 <= alu_loop_op_16_FpAdd_8U_23U_if_3_if_acc_2_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_15_itm <= 1'b0;
      IntLeadZero_49U_leading_sign_49_0_rtn_sva <= 6'b0;
    end
    else if ( FpNormalize_8U_49U_if_and_46_cse ) begin
      FpNormalize_8U_49U_if_or_15_itm <= FpNormalize_8U_49U_if_or_15_itm_mx0w0;
      IntLeadZero_49U_leading_sign_49_0_rtn_sva <= libraries_leading_sign_49_0_b604f59be2905c01c81f2d0a2ea3fe5a83a3_31;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_else_if_conc_itm_31 <= 1'b0;
      alu_loop_op_1_else_if_conc_itm_0 <= 1'b0;
      alu_loop_op_1_else_if_conc_itm_30_1 <= 30'b0;
      alu_loop_op_2_else_if_conc_1_itm_31 <= 1'b0;
      alu_loop_op_2_else_if_conc_1_itm_0 <= 1'b0;
      alu_loop_op_2_else_if_conc_1_itm_30_1 <= 30'b0;
      alu_loop_op_4_else_if_conc_1_itm_31 <= 1'b0;
      alu_loop_op_4_else_if_conc_1_itm_0 <= 1'b0;
      alu_loop_op_4_else_if_conc_1_itm_30_1 <= 30'b0;
    end
    else if ( alu_loop_op_else_if_and_cse ) begin
      alu_loop_op_1_else_if_conc_itm_31 <= alu_loop_op_else_else_if_mux_itm_2;
      alu_loop_op_1_else_if_conc_itm_0 <= alu_loop_op_else_else_if_mux_2_itm_2;
      alu_loop_op_1_else_if_conc_itm_30_1 <= alu_loop_op_else_else_if_mux_1_itm_2;
      alu_loop_op_2_else_if_conc_1_itm_31 <= alu_loop_op_else_else_if_mux_3_itm_2;
      alu_loop_op_2_else_if_conc_1_itm_0 <= alu_loop_op_else_else_if_mux_5_itm_2;
      alu_loop_op_2_else_if_conc_1_itm_30_1 <= alu_loop_op_else_else_if_mux_4_itm_2;
      alu_loop_op_4_else_if_conc_1_itm_31 <= alu_loop_op_else_else_if_mux_9_itm_2;
      alu_loop_op_4_else_if_conc_1_itm_0 <= alu_loop_op_else_else_if_mux_11_itm_2;
      alu_loop_op_4_else_if_conc_1_itm_30_1 <= alu_loop_op_else_else_if_mux_10_itm_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_else_else_if_conc_itm_31 <= 1'b0;
      alu_loop_op_1_else_else_if_conc_itm_0 <= 1'b0;
      alu_loop_op_1_else_else_if_conc_itm_30_1 <= 30'b0;
      alu_loop_op_2_else_else_if_conc_1_itm_31 <= 1'b0;
      alu_loop_op_2_else_else_if_conc_1_itm_0 <= 1'b0;
      alu_loop_op_2_else_else_if_conc_1_itm_30_1 <= 30'b0;
      alu_loop_op_4_else_else_if_conc_1_itm_31 <= 1'b0;
      alu_loop_op_4_else_else_if_conc_1_itm_0 <= 1'b0;
      alu_loop_op_4_else_else_if_conc_1_itm_30_1 <= 30'b0;
    end
    else if ( alu_loop_op_else_else_if_and_cse ) begin
      alu_loop_op_1_else_else_if_conc_itm_31 <= alu_loop_op_else_else_if_mux_itm_2;
      alu_loop_op_1_else_else_if_conc_itm_0 <= alu_loop_op_else_else_if_mux_2_itm_2;
      alu_loop_op_1_else_else_if_conc_itm_30_1 <= alu_loop_op_else_else_if_mux_1_itm_2;
      alu_loop_op_2_else_else_if_conc_1_itm_31 <= alu_loop_op_else_else_if_mux_3_itm_2;
      alu_loop_op_2_else_else_if_conc_1_itm_0 <= alu_loop_op_else_else_if_mux_5_itm_2;
      alu_loop_op_2_else_else_if_conc_1_itm_30_1 <= alu_loop_op_else_else_if_mux_4_itm_2;
      alu_loop_op_4_else_else_if_conc_1_itm_31 <= alu_loop_op_else_else_if_mux_9_itm_2;
      alu_loop_op_4_else_else_if_conc_1_itm_0 <= alu_loop_op_else_else_if_mux_11_itm_2;
      alu_loop_op_4_else_else_if_conc_1_itm_30_1 <= alu_loop_op_else_else_if_mux_10_itm_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_6_lpi_1_dfm_4_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_6_lpi_1_dfm_4_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_226_cse ) begin
      FpAdd_8U_23U_qr_6_lpi_1_dfm_4_7_4_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[158:155]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_9, FpAdd_8U_23U_qr_6_lpi_1_dfm_7_4,
          {and_dcpl_565 , and_dcpl_570 , and_dcpl_408});
      FpAdd_8U_23U_qr_6_lpi_1_dfm_4_3_0_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[154:151]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_9, FpAdd_8U_23U_qr_6_lpi_1_dfm_3_0,
          {and_dcpl_565 , and_dcpl_570 , and_dcpl_408});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_7_lpi_1_dfm_4_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_7_lpi_1_dfm_4_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_228_cse ) begin
      FpAdd_8U_23U_qr_7_lpi_1_dfm_4_7_4_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[190:187]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_9, FpAdd_8U_23U_qr_7_lpi_1_dfm_7_4,
          {and_dcpl_576 , and_dcpl_581 , and_dcpl_408});
      FpAdd_8U_23U_qr_7_lpi_1_dfm_4_3_0_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[186:183]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_9, FpAdd_8U_23U_qr_7_lpi_1_dfm_3_0,
          {and_dcpl_576 , and_dcpl_581 , and_dcpl_408});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_8_lpi_1_dfm_4_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_8_lpi_1_dfm_4_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_230_cse ) begin
      FpAdd_8U_23U_qr_8_lpi_1_dfm_4_7_4_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[222:219]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_9, FpAdd_8U_23U_qr_8_lpi_1_dfm_7_4,
          {and_dcpl_587 , and_dcpl_592 , and_dcpl_408});
      FpAdd_8U_23U_qr_8_lpi_1_dfm_4_3_0_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[218:215]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_9, FpAdd_8U_23U_qr_8_lpi_1_dfm_3_0,
          {and_dcpl_587 , and_dcpl_592 , and_dcpl_408});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_10_lpi_1_dfm_4_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_10_lpi_1_dfm_4_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_232_cse ) begin
      FpAdd_8U_23U_qr_10_lpi_1_dfm_4_7_4_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[286:283]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_9, FpAdd_8U_23U_qr_10_lpi_1_dfm_7_4,
          {and_dcpl_598 , and_dcpl_603 , and_dcpl_408});
      FpAdd_8U_23U_qr_10_lpi_1_dfm_4_3_0_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[282:279]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_9, FpAdd_8U_23U_qr_10_lpi_1_dfm_3_0,
          {and_dcpl_598 , and_dcpl_603 , and_dcpl_408});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_11_lpi_1_dfm_4_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_11_lpi_1_dfm_4_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_234_cse ) begin
      FpAdd_8U_23U_qr_11_lpi_1_dfm_4_7_4_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[318:315]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_9, FpAdd_8U_23U_qr_11_lpi_1_dfm_7_4,
          {and_dcpl_609 , and_dcpl_614 , and_dcpl_408});
      FpAdd_8U_23U_qr_11_lpi_1_dfm_4_3_0_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[314:311]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_9, FpAdd_8U_23U_qr_11_lpi_1_dfm_3_0,
          {and_dcpl_609 , and_dcpl_614 , and_dcpl_408});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_12_lpi_1_dfm_4_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_12_lpi_1_dfm_4_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_236_cse ) begin
      FpAdd_8U_23U_qr_12_lpi_1_dfm_4_7_4_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[350:347]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_9, FpAdd_8U_23U_qr_12_lpi_1_dfm_7_4,
          {and_dcpl_620 , and_dcpl_625 , and_dcpl_408});
      FpAdd_8U_23U_qr_12_lpi_1_dfm_4_3_0_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[346:343]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_9, FpAdd_8U_23U_qr_12_lpi_1_dfm_3_0,
          {and_dcpl_620 , and_dcpl_625 , and_dcpl_408});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_13_lpi_1_dfm_4_7_4_1 <= 4'b0;
      FpAdd_8U_23U_qr_13_lpi_1_dfm_4_3_0_1 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_238_cse ) begin
      FpAdd_8U_23U_qr_13_lpi_1_dfm_4_7_4_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[382:379]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_9, FpAdd_8U_23U_qr_13_lpi_1_dfm_7_4,
          {and_dcpl_631 , and_dcpl_636 , and_dcpl_408});
      FpAdd_8U_23U_qr_13_lpi_1_dfm_4_3_0_1 <= MUX1HOT_v_4_3_2((AluIn_data_sva_501[378:375]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_9, FpAdd_8U_23U_qr_13_lpi_1_dfm_3_0,
          {and_dcpl_631 , and_dcpl_636 , and_dcpl_408});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm
          <= 1'b0;
      alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_itm <= 8'b0;
      alu_loop_op_1_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm
          <= 1'b0;
      alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_itm <= 8'b0;
      alu_loop_op_2_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm
          <= 1'b0;
      alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_1_itm <= 8'b0;
      alu_loop_op_2_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm
          <= 1'b0;
      alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_1_itm <= 8'b0;
      alu_loop_op_3_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm
          <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_itm <= 8'b0;
      alu_loop_op_3_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm
          <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_itm <= 8'b0;
      alu_loop_op_4_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm
          <= 1'b0;
      alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_1_itm <= 8'b0;
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= 1'b0;
      alu_loop_op_4_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm
          <= 1'b0;
      alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_1_itm <= 8'b0;
      alu_loop_op_5_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm
          <= 1'b0;
      alu_loop_op_5_FpAdd_8U_23U_b_left_shift_acc_itm <= 8'b0;
      alu_loop_op_5_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm
          <= 1'b0;
      alu_loop_op_5_FpAdd_8U_23U_a_left_shift_acc_itm <= 8'b0;
      alu_loop_op_6_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm
          <= 1'b0;
      alu_loop_op_6_FpAdd_8U_23U_b_left_shift_acc_1_itm <= 8'b0;
      alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= 1'b0;
      alu_loop_op_6_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm
          <= 1'b0;
      alu_loop_op_6_FpAdd_8U_23U_a_left_shift_acc_1_itm <= 8'b0;
      alu_loop_op_7_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm
          <= 1'b0;
      alu_loop_op_7_FpAdd_8U_23U_b_left_shift_acc_itm <= 8'b0;
      alu_loop_op_7_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm
          <= 1'b0;
      alu_loop_op_7_FpAdd_8U_23U_a_left_shift_acc_itm <= 8'b0;
      alu_loop_op_8_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm
          <= 1'b0;
      alu_loop_op_8_FpAdd_8U_23U_b_left_shift_acc_1_itm <= 8'b0;
      alu_loop_op_8_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm
          <= 1'b0;
      alu_loop_op_8_FpAdd_8U_23U_a_left_shift_acc_1_itm <= 8'b0;
      alu_loop_op_9_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm
          <= 1'b0;
      alu_loop_op_9_FpAdd_8U_23U_b_left_shift_acc_itm <= 8'b0;
      alu_loop_op_9_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm
          <= 1'b0;
      alu_loop_op_9_FpAdd_8U_23U_a_left_shift_acc_itm <= 8'b0;
      alu_loop_op_10_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm
          <= 1'b0;
      alu_loop_op_10_FpAdd_8U_23U_b_left_shift_acc_1_itm <= 8'b0;
      alu_loop_op_10_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm
          <= 1'b0;
      alu_loop_op_10_FpAdd_8U_23U_a_left_shift_acc_1_itm <= 8'b0;
      alu_loop_op_11_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm
          <= 1'b0;
      alu_loop_op_11_FpAdd_8U_23U_b_left_shift_acc_itm <= 8'b0;
      alu_loop_op_11_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm
          <= 1'b0;
      alu_loop_op_11_FpAdd_8U_23U_a_left_shift_acc_itm <= 8'b0;
      alu_loop_op_12_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm
          <= 1'b0;
      alu_loop_op_12_FpAdd_8U_23U_b_left_shift_acc_1_itm <= 8'b0;
      alu_loop_op_12_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm
          <= 1'b0;
      alu_loop_op_12_FpAdd_8U_23U_a_left_shift_acc_1_itm <= 8'b0;
      alu_loop_op_13_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm
          <= 1'b0;
      alu_loop_op_13_FpAdd_8U_23U_b_left_shift_acc_itm <= 8'b0;
      alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= 1'b0;
      alu_loop_op_13_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm
          <= 1'b0;
      alu_loop_op_13_FpAdd_8U_23U_a_left_shift_acc_itm <= 8'b0;
      alu_loop_op_14_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm
          <= 1'b0;
      alu_loop_op_14_FpAdd_8U_23U_b_left_shift_acc_1_itm <= 8'b0;
      alu_loop_op_14_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm
          <= 1'b0;
      alu_loop_op_14_FpAdd_8U_23U_a_left_shift_acc_1_itm <= 8'b0;
      alu_loop_op_15_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm
          <= 1'b0;
      alu_loop_op_15_FpAdd_8U_23U_b_left_shift_acc_itm <= 8'b0;
      alu_loop_op_15_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm
          <= 1'b0;
      alu_loop_op_15_FpAdd_8U_23U_a_left_shift_acc_itm <= 8'b0;
      alu_loop_op_16_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm
          <= 1'b0;
      alu_loop_op_16_FpAdd_8U_23U_b_left_shift_acc_1_itm <= 8'b0;
      alu_loop_op_16_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm
          <= 1'b0;
      alu_loop_op_16_FpAdd_8U_23U_a_left_shift_acc_1_itm <= 8'b0;
    end
    else if ( FpAdd_8U_23U_b_left_shift_and_cse ) begin
      alu_loop_op_1_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm
          <= FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm[0];
      alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_itm <= alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
      alu_loop_op_1_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm
          <= FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm[0];
      alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_itm <= alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
      alu_loop_op_2_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm
          <= FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm[0];
      alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_1_itm <= alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
      alu_loop_op_2_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm
          <= FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm[0];
      alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_1_itm <= alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
      alu_loop_op_3_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm
          <= FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm[0];
      alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_itm <= alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
      alu_loop_op_3_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm
          <= FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm[0];
      alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_itm <= alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
      alu_loop_op_4_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm
          <= FpAdd_8U_23U_b_right_shift_qr_4_lpi_1_dfm[0];
      alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_1_itm <= alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
      alu_loop_op_4_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm
          <= FpAdd_8U_23U_a_right_shift_qr_4_lpi_1_dfm[0];
      alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_1_itm <= alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
      alu_loop_op_5_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm
          <= FpAdd_8U_23U_b_right_shift_qr_5_lpi_1_dfm[0];
      alu_loop_op_5_FpAdd_8U_23U_b_left_shift_acc_itm <= alu_loop_op_5_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
      alu_loop_op_5_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm
          <= FpAdd_8U_23U_a_right_shift_qr_5_lpi_1_dfm[0];
      alu_loop_op_5_FpAdd_8U_23U_a_left_shift_acc_itm <= alu_loop_op_5_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
      alu_loop_op_6_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm
          <= FpAdd_8U_23U_b_right_shift_qr_6_lpi_1_dfm[0];
      alu_loop_op_6_FpAdd_8U_23U_b_left_shift_acc_1_itm <= alu_loop_op_6_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
      alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
      alu_loop_op_6_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm
          <= FpAdd_8U_23U_a_right_shift_qr_6_lpi_1_dfm[0];
      alu_loop_op_6_FpAdd_8U_23U_a_left_shift_acc_1_itm <= alu_loop_op_6_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
      alu_loop_op_7_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm
          <= FpAdd_8U_23U_b_right_shift_qr_7_lpi_1_dfm[0];
      alu_loop_op_7_FpAdd_8U_23U_b_left_shift_acc_itm <= alu_loop_op_7_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
      alu_loop_op_7_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm
          <= FpAdd_8U_23U_a_right_shift_qr_7_lpi_1_dfm[0];
      alu_loop_op_7_FpAdd_8U_23U_a_left_shift_acc_itm <= alu_loop_op_7_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
      alu_loop_op_8_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm
          <= FpAdd_8U_23U_b_right_shift_qr_8_lpi_1_dfm[0];
      alu_loop_op_8_FpAdd_8U_23U_b_left_shift_acc_1_itm <= alu_loop_op_8_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
      alu_loop_op_8_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm
          <= FpAdd_8U_23U_a_right_shift_qr_8_lpi_1_dfm[0];
      alu_loop_op_8_FpAdd_8U_23U_a_left_shift_acc_1_itm <= alu_loop_op_8_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
      alu_loop_op_9_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm
          <= FpAdd_8U_23U_b_right_shift_qr_9_lpi_1_dfm[0];
      alu_loop_op_9_FpAdd_8U_23U_b_left_shift_acc_itm <= alu_loop_op_9_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
      alu_loop_op_9_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm
          <= FpAdd_8U_23U_a_right_shift_qr_9_lpi_1_dfm[0];
      alu_loop_op_9_FpAdd_8U_23U_a_left_shift_acc_itm <= alu_loop_op_9_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
      alu_loop_op_10_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm
          <= FpAdd_8U_23U_b_right_shift_qr_10_lpi_1_dfm[0];
      alu_loop_op_10_FpAdd_8U_23U_b_left_shift_acc_1_itm <= alu_loop_op_10_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
      alu_loop_op_10_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm
          <= FpAdd_8U_23U_a_right_shift_qr_10_lpi_1_dfm[0];
      alu_loop_op_10_FpAdd_8U_23U_a_left_shift_acc_1_itm <= alu_loop_op_10_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
      alu_loop_op_11_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm
          <= FpAdd_8U_23U_b_right_shift_qr_11_lpi_1_dfm[0];
      alu_loop_op_11_FpAdd_8U_23U_b_left_shift_acc_itm <= alu_loop_op_11_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
      alu_loop_op_11_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm
          <= FpAdd_8U_23U_a_right_shift_qr_11_lpi_1_dfm[0];
      alu_loop_op_11_FpAdd_8U_23U_a_left_shift_acc_itm <= alu_loop_op_11_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
      alu_loop_op_12_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm
          <= FpAdd_8U_23U_b_right_shift_qr_12_lpi_1_dfm[0];
      alu_loop_op_12_FpAdd_8U_23U_b_left_shift_acc_1_itm <= alu_loop_op_12_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
      alu_loop_op_12_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm
          <= FpAdd_8U_23U_a_right_shift_qr_12_lpi_1_dfm[0];
      alu_loop_op_12_FpAdd_8U_23U_a_left_shift_acc_1_itm <= alu_loop_op_12_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
      alu_loop_op_13_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm
          <= FpAdd_8U_23U_b_right_shift_qr_13_lpi_1_dfm[0];
      alu_loop_op_13_FpAdd_8U_23U_b_left_shift_acc_itm <= alu_loop_op_13_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
      alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
      alu_loop_op_13_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm
          <= FpAdd_8U_23U_a_right_shift_qr_13_lpi_1_dfm[0];
      alu_loop_op_13_FpAdd_8U_23U_a_left_shift_acc_itm <= alu_loop_op_13_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
      alu_loop_op_14_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm
          <= FpAdd_8U_23U_b_right_shift_qr_14_lpi_1_dfm[0];
      alu_loop_op_14_FpAdd_8U_23U_b_left_shift_acc_1_itm <= alu_loop_op_14_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
      alu_loop_op_14_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm
          <= FpAdd_8U_23U_a_right_shift_qr_14_lpi_1_dfm[0];
      alu_loop_op_14_FpAdd_8U_23U_a_left_shift_acc_1_itm <= alu_loop_op_14_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
      alu_loop_op_15_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_itm
          <= FpAdd_8U_23U_b_right_shift_qr_15_lpi_1_dfm[0];
      alu_loop_op_15_FpAdd_8U_23U_b_left_shift_acc_itm <= alu_loop_op_15_FpAdd_8U_23U_b_left_shift_acc_itm_mx0w0;
      alu_loop_op_15_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_itm
          <= FpAdd_8U_23U_a_right_shift_qr_15_lpi_1_dfm[0];
      alu_loop_op_15_FpAdd_8U_23U_a_left_shift_acc_itm <= alu_loop_op_15_FpAdd_8U_23U_a_left_shift_acc_itm_mx0w0;
      alu_loop_op_16_FpAdd_8U_23U_b_left_shift_slc_FpAdd_8U_23U_b_right_shift_0_1_itm
          <= FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm[0];
      alu_loop_op_16_FpAdd_8U_23U_b_left_shift_acc_1_itm <= alu_loop_op_16_FpAdd_8U_23U_b_left_shift_acc_1_itm_mx0w0;
      alu_loop_op_16_FpAdd_8U_23U_a_left_shift_slc_FpAdd_8U_23U_a_right_shift_0_1_itm
          <= FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm[0];
      alu_loop_op_16_FpAdd_8U_23U_a_left_shift_acc_1_itm <= alu_loop_op_16_FpAdd_8U_23U_a_left_shift_acc_1_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3 <= 1'b0;
      alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2 <= 1'b0;
    end
    else if ( IsZero_8U_23U_1_and_24_cse ) begin
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3 <= MUX_s_1_2_2(alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0,
          alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm, and_1106_rgt);
      alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2 <= MUX_s_1_2_2(alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0,
          alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm, and_1106_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2 <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3 <= 1'b0;
      alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2 <= 1'b0;
      alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3 <= 1'b0;
      alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3 <= 1'b0;
      alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2 <= 1'b0;
      alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2 <= 1'b0;
      alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2 <= 1'b0;
      alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2 <= 1'b0;
      alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3 <= 1'b0;
      alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3 <= 1'b0;
    end
    else if ( IsZero_8U_23U_1_and_25_cse ) begin
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2 <= MUX_s_1_2_2(alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0,
          alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm, and_1108_rgt);
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3 <= MUX_s_1_2_2(alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0,
          alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm, and_1108_rgt);
      alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2 <= MUX_s_1_2_2(alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0,
          alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm, and_1108_rgt);
      alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3 <= MUX_s_1_2_2(alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0,
          alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm, and_1108_rgt);
      alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3 <= MUX_s_1_2_2(alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0,
          alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm, and_1108_rgt);
      alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2 <= MUX_s_1_2_2(alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0,
          alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm, and_1108_rgt);
      alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2 <= MUX_s_1_2_2(alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0,
          alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm, and_1108_rgt);
      alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2 <= MUX_s_1_2_2(alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0,
          alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm, and_1108_rgt);
      alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2 <= MUX_s_1_2_2(alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0,
          alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm, and_1108_rgt);
      alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3 <= MUX_s_1_2_2(alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0,
          alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm, and_1108_rgt);
      alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_3 <= MUX_s_1_2_2(alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0,
          alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm, and_1108_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_1_aelse_or_5_cse & (~
        (mux_813_nl)) ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_1_land_lpi_1_dfm_7,
          IsNaN_8U_23U_4_land_lpi_1_dfm_6, IsNaN_8U_23U_1_aelse_or_5_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_15_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_14_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_13_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_12_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_11_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_10_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_9_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_8_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_7_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_6_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_5_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_4_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_47_cse ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_9 <= IsNaN_8U_23U_land_lpi_1_dfm_8;
      IsNaN_8U_23U_land_15_lpi_1_dfm_9 <= IsNaN_8U_23U_land_15_lpi_1_dfm_8;
      IsNaN_8U_23U_land_14_lpi_1_dfm_9 <= IsNaN_8U_23U_land_14_lpi_1_dfm_8;
      IsNaN_8U_23U_land_13_lpi_1_dfm_9 <= IsNaN_8U_23U_land_13_lpi_1_dfm_8;
      IsNaN_8U_23U_land_12_lpi_1_dfm_9 <= IsNaN_8U_23U_land_12_lpi_1_dfm_8;
      IsNaN_8U_23U_land_11_lpi_1_dfm_9 <= IsNaN_8U_23U_land_11_lpi_1_dfm_8;
      IsNaN_8U_23U_land_10_lpi_1_dfm_9 <= IsNaN_8U_23U_land_10_lpi_1_dfm_8;
      IsNaN_8U_23U_land_9_lpi_1_dfm_9 <= IsNaN_8U_23U_land_9_lpi_1_dfm_8;
      IsNaN_8U_23U_land_8_lpi_1_dfm_9 <= IsNaN_8U_23U_land_8_lpi_1_dfm_8;
      IsNaN_8U_23U_land_7_lpi_1_dfm_9 <= IsNaN_8U_23U_land_7_lpi_1_dfm_8;
      IsNaN_8U_23U_land_6_lpi_1_dfm_9 <= IsNaN_8U_23U_land_6_lpi_1_dfm_8;
      IsNaN_8U_23U_land_5_lpi_1_dfm_9 <= IsNaN_8U_23U_land_5_lpi_1_dfm_8;
      IsNaN_8U_23U_land_4_lpi_1_dfm_9 <= IsNaN_8U_23U_land_4_lpi_1_dfm_8;
      IsNaN_8U_23U_land_3_lpi_1_dfm_9 <= IsNaN_8U_23U_land_3_lpi_1_dfm_8;
      IsNaN_8U_23U_land_2_lpi_1_dfm_9 <= IsNaN_8U_23U_land_2_lpi_1_dfm_8;
      IsNaN_8U_23U_land_1_lpi_1_dfm_9 <= IsNaN_8U_23U_land_1_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_15_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_1_aelse_or_5_cse & (mux_825_nl)
        ) begin
      IsNaN_8U_23U_1_land_15_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_1_land_15_lpi_1_dfm_7,
          IsNaN_8U_23U_4_land_15_lpi_1_dfm_6, IsNaN_8U_23U_1_aelse_or_5_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_14_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_1_land_13_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_1_land_12_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_1_land_11_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_1_land_5_lpi_1_dfm_8 <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_10 <= 4'b0;
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_10 <= 4'b0;
      IsNaN_8U_23U_1_land_4_lpi_1_dfm_8 <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_10 <= 4'b0;
      IsNaN_8U_23U_1_land_6_lpi_1_dfm_8 <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_10 <= 4'b0;
      IsNaN_8U_23U_1_land_9_lpi_1_dfm_8 <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_10 <= 4'b0;
      IsNaN_8U_23U_1_land_10_lpi_1_dfm_8 <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_10 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( IsNaN_8U_23U_1_aelse_and_34_cse ) begin
      IsNaN_8U_23U_1_land_14_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_14_lpi_1_dfm_7;
      IsNaN_8U_23U_1_land_13_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_13_lpi_1_dfm_7;
      IsNaN_8U_23U_1_land_12_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_12_lpi_1_dfm_7;
      IsNaN_8U_23U_1_land_11_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_11_lpi_1_dfm_7;
      IsNaN_8U_23U_1_land_5_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_5_lpi_1_dfm_7;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_9;
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_9;
      IsNaN_8U_23U_1_land_4_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_4_lpi_1_dfm_7;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_9;
      IsNaN_8U_23U_1_land_6_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_6_lpi_1_dfm_7;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_9;
      IsNaN_8U_23U_1_land_9_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_9_lpi_1_dfm_7;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_9;
      IsNaN_8U_23U_1_land_10_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_10_lpi_1_dfm_7;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_9;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_8_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_1_aelse_or_3_cse & (mux_857_nl)
        ) begin
      IsNaN_8U_23U_1_land_8_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_1_land_8_lpi_1_dfm_7,
          IsNaN_8U_23U_4_land_8_lpi_1_dfm_6, IsNaN_8U_23U_1_aelse_or_3_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_7_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_1_aelse_or_5_cse & (~
        (mux_870_nl)) ) begin
      IsNaN_8U_23U_1_land_7_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_1_land_7_lpi_1_dfm_7,
          IsNaN_8U_23U_4_land_7_lpi_1_dfm_6, IsNaN_8U_23U_1_aelse_or_5_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_1_aelse_or_3_cse & (mux_892_nl)
        ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_1_land_3_lpi_1_dfm_7,
          IsNaN_8U_23U_4_land_3_lpi_1_dfm_6, IsNaN_8U_23U_1_aelse_or_3_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_1_aelse_or_5_cse & (~
        (mux_908_nl)) ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_1_land_1_lpi_1_dfm_7,
          IsNaN_8U_23U_4_land_1_lpi_1_dfm_6, IsNaN_8U_23U_1_aelse_or_5_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      AluOut_data_15_sva_7 <= 33'b0;
      AluOut_data_14_sva_7 <= 33'b0;
      AluOut_data_13_sva_7 <= 33'b0;
      AluOut_data_12_sva_7 <= 33'b0;
      AluOut_data_11_sva_7 <= 33'b0;
      AluOut_data_10_sva_7 <= 33'b0;
      AluOut_data_9_sva_7 <= 33'b0;
      AluOut_data_8_sva_7 <= 33'b0;
      AluOut_data_7_sva_7 <= 33'b0;
      AluOut_data_6_sva_7 <= 33'b0;
      AluOut_data_5_sva_7 <= 33'b0;
      AluOut_data_4_sva_7 <= 33'b0;
      AluOut_data_3_sva_7 <= 33'b0;
      AluOut_data_2_sva_7 <= 33'b0;
      AluOut_data_1_sva_7 <= 33'b0;
      AluOut_data_0_sva_7 <= 33'b0;
    end
    else if ( AluOut_data_and_16_cse ) begin
      AluOut_data_15_sva_7 <= nl_AluOut_data_15_sva_7[32:0];
      AluOut_data_14_sva_7 <= nl_AluOut_data_14_sva_7[32:0];
      AluOut_data_13_sva_7 <= nl_AluOut_data_13_sva_7[32:0];
      AluOut_data_12_sva_7 <= nl_AluOut_data_12_sva_7[32:0];
      AluOut_data_11_sva_7 <= nl_AluOut_data_11_sva_7[32:0];
      AluOut_data_10_sva_7 <= nl_AluOut_data_10_sva_7[32:0];
      AluOut_data_9_sva_7 <= nl_AluOut_data_9_sva_7[32:0];
      AluOut_data_8_sva_7 <= nl_AluOut_data_8_sva_7[32:0];
      AluOut_data_7_sva_7 <= nl_AluOut_data_7_sva_7[32:0];
      AluOut_data_6_sva_7 <= nl_AluOut_data_6_sva_7[32:0];
      AluOut_data_5_sva_7 <= nl_AluOut_data_5_sva_7[32:0];
      AluOut_data_4_sva_7 <= nl_AluOut_data_4_sva_7[32:0];
      AluOut_data_3_sva_7 <= nl_AluOut_data_3_sva_7[32:0];
      AluOut_data_2_sva_7 <= nl_AluOut_data_2_sva_7[32:0];
      AluOut_data_1_sva_7 <= nl_AluOut_data_1_sva_7[32:0];
      AluOut_data_0_sva_7 <= nl_AluOut_data_0_sva_7[32:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_o_0_sva_6 <= 1'b0;
      FpAlu_8U_23U_o_0_15_sva_6 <= 1'b0;
      FpAlu_8U_23U_o_0_14_sva_6 <= 1'b0;
      FpAlu_8U_23U_o_0_13_sva_6 <= 1'b0;
      FpAlu_8U_23U_o_0_12_sva_6 <= 1'b0;
      FpAlu_8U_23U_o_0_11_sva_6 <= 1'b0;
      FpAlu_8U_23U_o_0_10_sva_6 <= 1'b0;
      FpAlu_8U_23U_o_0_9_sva_6 <= 1'b0;
      FpAlu_8U_23U_o_0_8_sva_6 <= 1'b0;
      FpAlu_8U_23U_o_0_7_sva_6 <= 1'b0;
      FpAlu_8U_23U_o_0_6_sva_6 <= 1'b0;
      FpAlu_8U_23U_o_0_5_sva_6 <= 1'b0;
      FpAlu_8U_23U_o_0_4_sva_6 <= 1'b0;
      FpAlu_8U_23U_o_0_3_sva_6 <= 1'b0;
      FpAlu_8U_23U_o_0_2_sva_6 <= 1'b0;
      FpAlu_8U_23U_o_0_1_sva_6 <= 1'b0;
    end
    else if ( FpAlu_8U_23U_o_and_16_cse ) begin
      FpAlu_8U_23U_o_0_sva_6 <= (AluIn_data_sva_501[511:480]) != ({alu_nan_to_zero_op_sign_lpi_1_dfm_3
          , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_9
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp_2});
      FpAlu_8U_23U_o_0_15_sva_6 <= (AluIn_data_sva_501[479:448]) != ({alu_nan_to_zero_op_sign_15_lpi_1_dfm_3
          , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_9
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_6_tmp_2});
      FpAlu_8U_23U_o_0_14_sva_6 <= (AluIn_data_sva_501[447:416]) != ({alu_nan_to_zero_op_sign_14_lpi_1_dfm_3
          , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_9
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_6_tmp_2});
      FpAlu_8U_23U_o_0_13_sva_6 <= (AluIn_data_sva_501[415:384]) != ({alu_nan_to_zero_op_sign_13_lpi_1_dfm_3
          , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_9
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp_2});
      FpAlu_8U_23U_o_0_12_sva_6 <= (AluIn_data_sva_501[383:352]) != ({alu_nan_to_zero_op_sign_12_lpi_1_dfm_3
          , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_9
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp_2});
      FpAlu_8U_23U_o_0_11_sva_6 <= (AluIn_data_sva_501[351:320]) != ({alu_nan_to_zero_op_sign_11_lpi_1_dfm_3
          , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_9
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp_2});
      FpAlu_8U_23U_o_0_10_sva_6 <= (AluIn_data_sva_501[319:288]) != ({alu_nan_to_zero_op_sign_10_lpi_1_dfm_3
          , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_9
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp_2});
      FpAlu_8U_23U_o_0_9_sva_6 <= (AluIn_data_sva_501[287:256]) != ({alu_nan_to_zero_op_sign_9_lpi_1_dfm_3
          , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_9
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp_2});
      FpAlu_8U_23U_o_0_8_sva_6 <= (AluIn_data_sva_501[255:224]) != ({alu_nan_to_zero_op_sign_8_lpi_1_dfm_3
          , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_9
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp_2});
      FpAlu_8U_23U_o_0_7_sva_6 <= (AluIn_data_sva_501[223:192]) != ({alu_nan_to_zero_op_sign_7_lpi_1_dfm_4
          , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_9
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp_2});
      FpAlu_8U_23U_o_0_6_sva_6 <= (AluIn_data_sva_501[191:160]) != ({alu_nan_to_zero_op_sign_6_lpi_1_dfm_4
          , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_9
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp_2});
      FpAlu_8U_23U_o_0_5_sva_6 <= (AluIn_data_sva_501[159:128]) != ({alu_nan_to_zero_op_sign_5_lpi_1_dfm_4
          , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_9
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp_2});
      FpAlu_8U_23U_o_0_4_sva_6 <= (AluIn_data_sva_501[127:96]) != ({alu_nan_to_zero_op_sign_4_lpi_1_dfm_4
          , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_9
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp_2});
      FpAlu_8U_23U_o_0_3_sva_6 <= (AluIn_data_sva_501[95:64]) != ({alu_nan_to_zero_op_sign_3_lpi_1_dfm_4
          , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_9
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp_2});
      FpAlu_8U_23U_o_0_2_sva_6 <= (AluIn_data_sva_501[63:32]) != ({alu_nan_to_zero_op_sign_2_lpi_1_dfm_4
          , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_9
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp_2});
      FpAlu_8U_23U_o_0_1_sva_6 <= (AluIn_data_sva_501[31:0]) != ({alu_nan_to_zero_op_sign_1_lpi_1_dfm_4
          , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_9
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp_1
          , reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp_2});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_6_itm_3 <= 1'b0;
      alu_loop_op_else_else_if_mux_7_itm_3 <= 30'b0;
      alu_loop_op_else_else_if_mux_8_itm_3 <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_105_cse ) begin
      alu_loop_op_else_else_if_mux_6_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[95]),
          IntShiftLeft_16U_6U_32U_return_31_3_sva_2, alu_loop_op_else_else_if_mux_6_itm,
          alu_loop_op_else_if_mux_6_itm, {and_dcpl_698 , and_dcpl_701 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_7_itm_3 <= MUX1HOT_v_30_4_2((AluIn_data_sva_501[94:65]),
          IntShiftLeft_16U_6U_32U_return_30_1_3_sva_2, alu_loop_op_else_else_if_mux_7_itm,
          alu_loop_op_else_if_mux_7_itm, {and_dcpl_698 , and_dcpl_701 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_8_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[64]),
          IntShiftLeft_16U_6U_32U_return_0_3_sva_2, alu_loop_op_else_else_if_mux_8_itm,
          alu_loop_op_else_if_mux_8_itm, {and_dcpl_698 , and_dcpl_701 , and_dcpl_704
          , and_dcpl_707});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_12_itm_3 <= 1'b0;
      alu_loop_op_else_else_if_mux_13_itm_3 <= 30'b0;
      alu_loop_op_else_else_if_mux_14_itm_3 <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_108_cse ) begin
      alu_loop_op_else_else_if_mux_12_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[159]),
          IntShiftLeft_16U_6U_32U_return_31_5_sva_2, alu_loop_op_else_else_if_mux_12_itm,
          alu_loop_op_else_if_mux_12_itm, {and_dcpl_711 , and_dcpl_714 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_13_itm_3 <= MUX1HOT_v_30_4_2((AluIn_data_sva_501[158:129]),
          IntShiftLeft_16U_6U_32U_return_30_1_5_sva_2, alu_loop_op_else_else_if_mux_13_itm,
          alu_loop_op_else_if_mux_13_itm, {and_dcpl_711 , and_dcpl_714 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_14_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[128]),
          IntShiftLeft_16U_6U_32U_return_0_5_sva_2, alu_loop_op_else_else_if_mux_14_itm,
          alu_loop_op_else_if_mux_14_itm, {and_dcpl_711 , and_dcpl_714 , and_dcpl_704
          , and_dcpl_707});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_15_itm_3 <= 1'b0;
      alu_loop_op_else_else_if_mux_16_itm_3 <= 30'b0;
      alu_loop_op_else_else_if_mux_17_itm_3 <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_111_cse ) begin
      alu_loop_op_else_else_if_mux_15_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[191]),
          IntShiftLeft_16U_6U_32U_return_31_6_sva_2, alu_loop_op_else_else_if_mux_15_itm,
          alu_loop_op_else_if_mux_15_itm, {and_dcpl_722 , and_dcpl_725 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_16_itm_3 <= MUX1HOT_v_30_4_2((AluIn_data_sva_501[190:161]),
          IntShiftLeft_16U_6U_32U_return_30_1_6_sva_2, alu_loop_op_else_else_if_mux_16_itm,
          alu_loop_op_else_if_mux_16_itm, {and_dcpl_722 , and_dcpl_725 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_17_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[160]),
          IntShiftLeft_16U_6U_32U_return_0_6_sva_2, alu_loop_op_else_else_if_mux_17_itm,
          alu_loop_op_else_if_mux_17_itm, {and_dcpl_722 , and_dcpl_725 , and_dcpl_704
          , and_dcpl_707});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_18_itm_3 <= 1'b0;
      alu_loop_op_else_else_if_mux_19_itm_3 <= 30'b0;
      alu_loop_op_else_else_if_mux_20_itm_3 <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_114_cse ) begin
      alu_loop_op_else_else_if_mux_18_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[223]),
          IntShiftLeft_16U_6U_32U_return_31_7_sva_2, alu_loop_op_else_else_if_mux_18_itm,
          alu_loop_op_else_if_mux_18_itm, {and_dcpl_733 , and_dcpl_736 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_19_itm_3 <= MUX1HOT_v_30_4_2((AluIn_data_sva_501[222:193]),
          IntShiftLeft_16U_6U_32U_return_30_1_7_sva_2, alu_loop_op_else_else_if_mux_19_itm,
          alu_loop_op_else_if_mux_19_itm, {and_dcpl_733 , and_dcpl_736 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_20_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[192]),
          IntShiftLeft_16U_6U_32U_return_0_7_sva_2, alu_loop_op_else_else_if_mux_20_itm,
          alu_loop_op_else_if_mux_20_itm, {and_dcpl_733 , and_dcpl_736 , and_dcpl_704
          , and_dcpl_707});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_21_itm_3 <= 1'b0;
      alu_loop_op_else_else_if_mux_22_itm_3 <= 30'b0;
      alu_loop_op_else_else_if_mux_23_itm_3 <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_117_cse ) begin
      alu_loop_op_else_else_if_mux_21_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[255]),
          IntShiftLeft_16U_6U_32U_return_31_8_sva_2, alu_loop_op_else_else_if_mux_21_itm,
          alu_loop_op_else_if_mux_21_itm, {and_dcpl_744 , and_dcpl_747 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_22_itm_3 <= MUX1HOT_v_30_4_2((AluIn_data_sva_501[254:225]),
          IntShiftLeft_16U_6U_32U_return_30_1_8_sva_2, alu_loop_op_else_else_if_mux_22_itm,
          alu_loop_op_else_if_mux_22_itm, {and_dcpl_744 , and_dcpl_747 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_23_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[224]),
          IntShiftLeft_16U_6U_32U_return_0_8_sva_2, alu_loop_op_else_else_if_mux_23_itm,
          alu_loop_op_else_if_mux_23_itm, {and_dcpl_744 , and_dcpl_747 , and_dcpl_704
          , and_dcpl_707});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_24_itm_3 <= 1'b0;
      alu_loop_op_else_else_if_mux_25_itm_3 <= 30'b0;
      alu_loop_op_else_else_if_mux_26_itm_3 <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_120_cse ) begin
      alu_loop_op_else_else_if_mux_24_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[287]),
          IntShiftLeft_16U_6U_32U_return_31_9_sva_2, alu_loop_op_else_else_if_mux_24_itm,
          alu_loop_op_else_if_mux_24_itm, {and_dcpl_755 , and_dcpl_758 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_25_itm_3 <= MUX1HOT_v_30_4_2((AluIn_data_sva_501[286:257]),
          IntShiftLeft_16U_6U_32U_return_30_1_9_sva_2, alu_loop_op_else_else_if_mux_25_itm,
          alu_loop_op_else_if_mux_25_itm, {and_dcpl_755 , and_dcpl_758 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_26_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[256]),
          IntShiftLeft_16U_6U_32U_return_0_9_sva_2, alu_loop_op_else_else_if_mux_26_itm,
          alu_loop_op_else_if_mux_26_itm, {and_dcpl_755 , and_dcpl_758 , and_dcpl_704
          , and_dcpl_707});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_27_itm_3 <= 1'b0;
      alu_loop_op_else_else_if_mux_28_itm_3 <= 30'b0;
      alu_loop_op_else_else_if_mux_29_itm_3 <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_123_cse ) begin
      alu_loop_op_else_else_if_mux_27_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[319]),
          IntShiftLeft_16U_6U_32U_return_31_10_sva_2, alu_loop_op_else_else_if_mux_27_itm,
          alu_loop_op_else_if_mux_27_itm, {and_dcpl_766 , and_dcpl_769 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_28_itm_3 <= MUX1HOT_v_30_4_2((AluIn_data_sva_501[318:289]),
          IntShiftLeft_16U_6U_32U_return_30_1_10_sva_2, alu_loop_op_else_else_if_mux_28_itm,
          alu_loop_op_else_if_mux_28_itm, {and_dcpl_766 , and_dcpl_769 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_29_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[288]),
          IntShiftLeft_16U_6U_32U_return_0_10_sva_2, alu_loop_op_else_else_if_mux_29_itm,
          alu_loop_op_else_if_mux_29_itm, {and_dcpl_766 , and_dcpl_769 , and_dcpl_704
          , and_dcpl_707});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_30_itm_3 <= 1'b0;
      alu_loop_op_else_else_if_mux_31_itm_3 <= 30'b0;
      alu_loop_op_else_else_if_mux_32_itm_3 <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_126_cse ) begin
      alu_loop_op_else_else_if_mux_30_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[351]),
          IntShiftLeft_16U_6U_32U_return_31_11_sva_2, alu_loop_op_else_else_if_mux_30_itm,
          alu_loop_op_else_if_mux_30_itm, {and_dcpl_777 , and_dcpl_780 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_31_itm_3 <= MUX1HOT_v_30_4_2((AluIn_data_sva_501[350:321]),
          IntShiftLeft_16U_6U_32U_return_30_1_11_sva_2, alu_loop_op_else_else_if_mux_31_itm,
          alu_loop_op_else_if_mux_31_itm, {and_dcpl_777 , and_dcpl_780 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_32_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[320]),
          IntShiftLeft_16U_6U_32U_return_0_11_sva_2, alu_loop_op_else_else_if_mux_32_itm,
          alu_loop_op_else_if_mux_32_itm, {and_dcpl_777 , and_dcpl_780 , and_dcpl_704
          , and_dcpl_707});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_33_itm_3 <= 1'b0;
      alu_loop_op_else_else_if_mux_34_itm_3 <= 30'b0;
      alu_loop_op_else_else_if_mux_35_itm_3 <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_129_cse ) begin
      alu_loop_op_else_else_if_mux_33_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[383]),
          IntShiftLeft_16U_6U_32U_return_31_12_sva_2, alu_loop_op_else_else_if_mux_33_itm,
          alu_loop_op_else_if_mux_33_itm, {and_dcpl_788 , and_dcpl_791 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_34_itm_3 <= MUX1HOT_v_30_4_2((AluIn_data_sva_501[382:353]),
          IntShiftLeft_16U_6U_32U_return_30_1_12_sva_2, alu_loop_op_else_else_if_mux_34_itm,
          alu_loop_op_else_if_mux_34_itm, {and_dcpl_788 , and_dcpl_791 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_35_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[352]),
          IntShiftLeft_16U_6U_32U_return_0_12_sva_2, alu_loop_op_else_else_if_mux_35_itm,
          alu_loop_op_else_if_mux_35_itm, {and_dcpl_788 , and_dcpl_791 , and_dcpl_704
          , and_dcpl_707});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_36_itm_3 <= 1'b0;
      alu_loop_op_else_else_if_mux_37_itm_3 <= 30'b0;
      alu_loop_op_else_else_if_mux_38_itm_3 <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_132_cse ) begin
      alu_loop_op_else_else_if_mux_36_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[415]),
          IntShiftLeft_16U_6U_32U_return_31_13_sva_2, alu_loop_op_else_else_if_mux_36_itm,
          alu_loop_op_else_if_mux_36_itm, {and_dcpl_799 , and_dcpl_802 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_37_itm_3 <= MUX1HOT_v_30_4_2((AluIn_data_sva_501[414:385]),
          IntShiftLeft_16U_6U_32U_return_30_1_13_sva_2, alu_loop_op_else_else_if_mux_37_itm,
          alu_loop_op_else_if_mux_37_itm, {and_dcpl_799 , and_dcpl_802 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_38_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[384]),
          IntShiftLeft_16U_6U_32U_return_0_13_sva_2, alu_loop_op_else_else_if_mux_38_itm,
          alu_loop_op_else_if_mux_38_itm, {and_dcpl_799 , and_dcpl_802 , and_dcpl_704
          , and_dcpl_707});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_39_itm_3 <= 1'b0;
      alu_loop_op_else_else_if_mux_40_itm_3 <= 30'b0;
      alu_loop_op_else_else_if_mux_41_itm_3 <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_135_cse ) begin
      alu_loop_op_else_else_if_mux_39_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[447]),
          IntShiftLeft_16U_6U_32U_return_31_14_sva_2, alu_loop_op_else_else_if_mux_39_itm,
          alu_loop_op_else_if_mux_39_itm, {and_dcpl_810 , and_dcpl_813 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_40_itm_3 <= MUX1HOT_v_30_4_2((AluIn_data_sva_501[446:417]),
          IntShiftLeft_16U_6U_32U_return_30_1_14_sva_2, alu_loop_op_else_else_if_mux_40_itm,
          alu_loop_op_else_if_mux_40_itm, {and_dcpl_810 , and_dcpl_813 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_41_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[416]),
          IntShiftLeft_16U_6U_32U_return_0_14_sva_2, alu_loop_op_else_else_if_mux_41_itm,
          alu_loop_op_else_if_mux_41_itm, {and_dcpl_810 , and_dcpl_813 , and_dcpl_704
          , and_dcpl_707});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_42_itm_3 <= 1'b0;
      alu_loop_op_else_else_if_mux_43_itm_3 <= 30'b0;
      alu_loop_op_else_else_if_mux_44_itm_3 <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_138_cse ) begin
      alu_loop_op_else_else_if_mux_42_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[479]),
          IntShiftLeft_16U_6U_32U_return_31_15_sva_2, alu_loop_op_else_else_if_mux_42_itm,
          alu_loop_op_else_if_mux_42_itm, {and_dcpl_821 , and_dcpl_824 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_43_itm_3 <= MUX1HOT_v_30_4_2((AluIn_data_sva_501[478:449]),
          IntShiftLeft_16U_6U_32U_return_30_1_15_sva_2, alu_loop_op_else_else_if_mux_43_itm,
          alu_loop_op_else_if_mux_43_itm, {and_dcpl_821 , and_dcpl_824 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_44_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[448]),
          IntShiftLeft_16U_6U_32U_return_0_15_sva_2, alu_loop_op_else_else_if_mux_44_itm,
          alu_loop_op_else_if_mux_44_itm, {and_dcpl_821 , and_dcpl_824 , and_dcpl_704
          , and_dcpl_707});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_45_itm_3 <= 1'b0;
      alu_loop_op_else_else_if_mux_46_itm_3 <= 30'b0;
      alu_loop_op_else_else_if_mux_47_itm_3 <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_141_cse ) begin
      alu_loop_op_else_else_if_mux_45_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[511]),
          IntShiftLeft_16U_6U_32U_return_31_sva_2, alu_loop_op_else_else_if_mux_45_itm,
          alu_loop_op_else_if_mux_45_itm, {and_dcpl_832 , and_dcpl_834 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_46_itm_3 <= MUX1HOT_v_30_4_2((AluIn_data_sva_501[510:481]),
          IntShiftLeft_16U_6U_32U_return_30_1_sva_2, alu_loop_op_else_else_if_mux_46_itm,
          alu_loop_op_else_if_mux_46_itm, {and_dcpl_832 , and_dcpl_834 , and_dcpl_704
          , and_dcpl_707});
      alu_loop_op_else_else_if_mux_47_itm_3 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[480]),
          IntShiftLeft_16U_6U_32U_return_0_sva_2, alu_loop_op_else_else_if_mux_47_itm,
          alu_loop_op_else_if_mux_47_itm, {and_dcpl_832 , and_dcpl_834 , and_dcpl_704
          , and_dcpl_707});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_or_831_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_752_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_833_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_755_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_835_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_758_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_837_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_761_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_839_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_764_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_841_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_767_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_843_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_770_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_845_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_773_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_847_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_776_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_849_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_779_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_851_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_782_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_853_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_785_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_855_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_788_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_857_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_791_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_859_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_794_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_861_itm_3 <= 1'b0;
      FpAlu_8U_23U_or_797_itm_3 <= 1'b0;
    end
    else if ( FpAlu_8U_23U_and_976_cse ) begin
      FpAlu_8U_23U_or_831_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_831_itm_mx0w0, FpAlu_8U_23U_or_832_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_752_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_752_itm_mx0w0, FpAlu_8U_23U_or_753_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_833_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_833_itm_mx0w0, FpAlu_8U_23U_or_834_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_755_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_755_itm_mx0w0, FpAlu_8U_23U_or_756_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_835_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_835_itm_mx0w0, FpAlu_8U_23U_or_836_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_758_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_758_itm_mx0w0, FpAlu_8U_23U_or_759_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_837_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_837_itm_mx0w0, FpAlu_8U_23U_or_838_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_761_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_761_itm_mx0w0, FpAlu_8U_23U_or_762_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_839_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_839_itm_mx0w0, FpAlu_8U_23U_or_840_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_764_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_764_itm_mx0w0, FpAlu_8U_23U_or_765_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_841_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_841_itm_mx0w0, FpAlu_8U_23U_or_842_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_767_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_767_itm_mx0w0, FpAlu_8U_23U_or_768_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_843_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_843_itm_mx0w0, FpAlu_8U_23U_or_844_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_770_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_770_itm_mx0w0, FpAlu_8U_23U_or_771_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_845_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_845_itm_mx0w0, FpAlu_8U_23U_or_846_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_773_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_773_itm_mx0w0, FpAlu_8U_23U_or_774_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_847_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_847_itm_mx0w0, FpAlu_8U_23U_or_848_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_776_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_776_itm_mx0w0, FpAlu_8U_23U_or_777_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_849_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_849_itm_mx0w0, FpAlu_8U_23U_or_850_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_779_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_779_itm_mx0w0, FpAlu_8U_23U_or_780_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_851_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_851_itm_mx0w0, FpAlu_8U_23U_or_852_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_782_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_782_itm_mx0w0, FpAlu_8U_23U_or_783_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_853_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_853_itm_mx0w0, FpAlu_8U_23U_or_854_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_785_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_785_itm_mx0w0, FpAlu_8U_23U_or_786_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_855_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_855_itm_mx0w0, FpAlu_8U_23U_or_856_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_788_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_788_itm_mx0w0, FpAlu_8U_23U_or_789_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_857_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_857_itm_mx0w0, FpAlu_8U_23U_or_858_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_791_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_791_itm_mx0w0, FpAlu_8U_23U_or_792_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_859_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_859_itm_mx0w0, FpAlu_8U_23U_or_860_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_794_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_794_itm_mx0w0, FpAlu_8U_23U_or_795_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_861_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_861_itm_mx0w0, FpAlu_8U_23U_or_862_itm,
          and_dcpl_241);
      FpAlu_8U_23U_or_797_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_or_797_itm_mx0w0, FpAlu_8U_23U_or_798_itm,
          and_dcpl_241);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_and_itm_3 <= 1'b0;
      FpAlu_8U_23U_and_4_itm_3 <= 1'b0;
      FpAlu_8U_23U_and_8_itm_3 <= 1'b0;
      FpAlu_8U_23U_and_12_itm_3 <= 1'b0;
      FpAlu_8U_23U_and_16_itm_3 <= 1'b0;
      FpAlu_8U_23U_and_20_itm_3 <= 1'b0;
      FpAlu_8U_23U_and_24_itm_3 <= 1'b0;
      FpAlu_8U_23U_and_28_itm_3 <= 1'b0;
      FpAlu_8U_23U_and_32_itm_3 <= 1'b0;
      FpAlu_8U_23U_and_36_itm_3 <= 1'b0;
      FpAlu_8U_23U_and_40_itm_3 <= 1'b0;
      FpAlu_8U_23U_and_44_itm_3 <= 1'b0;
      FpAlu_8U_23U_and_48_itm_3 <= 1'b0;
      FpAlu_8U_23U_and_52_itm_3 <= 1'b0;
      FpAlu_8U_23U_and_56_itm_3 <= 1'b0;
      FpAlu_8U_23U_and_60_itm_3 <= 1'b0;
    end
    else if ( FpAlu_8U_23U_and_1040_cse ) begin
      FpAlu_8U_23U_and_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_and_itm_mx0w0, FpAlu_8U_23U_and_itm,
          and_dcpl_840);
      FpAlu_8U_23U_and_4_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_and_4_itm_mx0w0, FpAlu_8U_23U_and_4_itm,
          and_dcpl_840);
      FpAlu_8U_23U_and_8_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_and_8_itm_mx0w0, FpAlu_8U_23U_and_8_itm,
          and_dcpl_840);
      FpAlu_8U_23U_and_12_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_and_12_itm_mx0w0, FpAlu_8U_23U_and_12_itm,
          and_dcpl_840);
      FpAlu_8U_23U_and_16_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_and_16_itm_mx0w0, FpAlu_8U_23U_and_16_itm,
          and_dcpl_840);
      FpAlu_8U_23U_and_20_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_and_20_itm_mx0w0, FpAlu_8U_23U_and_20_itm,
          and_dcpl_840);
      FpAlu_8U_23U_and_24_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_and_24_itm_mx0w0, FpAlu_8U_23U_and_24_itm,
          and_dcpl_840);
      FpAlu_8U_23U_and_28_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_and_28_itm_mx0w0, FpAlu_8U_23U_and_28_itm,
          and_dcpl_840);
      FpAlu_8U_23U_and_32_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_and_32_itm_mx0w0, FpAlu_8U_23U_and_32_itm,
          and_dcpl_840);
      FpAlu_8U_23U_and_36_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_and_36_itm_mx0w0, FpAlu_8U_23U_and_36_itm,
          and_dcpl_840);
      FpAlu_8U_23U_and_40_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_and_40_itm_mx0w0, FpAlu_8U_23U_and_40_itm,
          and_dcpl_840);
      FpAlu_8U_23U_and_44_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_and_44_itm_mx0w0, FpAlu_8U_23U_and_44_itm,
          and_dcpl_840);
      FpAlu_8U_23U_and_48_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_and_48_itm_mx0w0, FpAlu_8U_23U_and_48_itm,
          and_dcpl_840);
      FpAlu_8U_23U_and_52_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_and_52_itm_mx0w0, FpAlu_8U_23U_and_52_itm,
          and_dcpl_840);
      FpAlu_8U_23U_and_56_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_and_56_itm_mx0w0, FpAlu_8U_23U_and_56_itm,
          and_dcpl_840);
      FpAlu_8U_23U_and_60_itm_3 <= MUX_s_1_2_2(FpAlu_8U_23U_and_60_itm_mx0w0, FpAlu_8U_23U_and_60_itm,
          and_dcpl_840);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_equal_tmp_144 <= 1'b0;
      FpAlu_8U_23U_equal_tmp_146 <= 1'b0;
      FpAlu_8U_23U_equal_tmp_148 <= 1'b0;
      FpAlu_8U_23U_nor_dfs_48 <= 1'b0;
    end
    else if ( FpAlu_8U_23U_and_1056_cse ) begin
      FpAlu_8U_23U_equal_tmp_144 <= MUX_s_1_2_2(FpAlu_8U_23U_equal_tmp_mx0w0, FpAlu_8U_23U_equal_tmp,
          and_dcpl_840);
      FpAlu_8U_23U_equal_tmp_146 <= MUX_s_1_2_2(and_3689_cse, FpAlu_8U_23U_equal_tmp_1,
          and_dcpl_840);
      FpAlu_8U_23U_equal_tmp_148 <= MUX_s_1_2_2(FpAlu_8U_23U_equal_tmp_2_mx0w0, FpAlu_8U_23U_equal_tmp_2,
          and_dcpl_840);
      FpAlu_8U_23U_nor_dfs_48 <= MUX_s_1_2_2(FpAlu_8U_23U_nor_dfs_mx0w0, FpAlu_8U_23U_nor_dfs,
          and_dcpl_840);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_3_land_1_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_2_land_2_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_2_land_4_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_2_land_5_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_3_land_7_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_2_land_9_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_2_land_11_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_2_land_12_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_3_land_15_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_3_land_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_3_aelse_and_cse ) begin
      IsNaN_8U_23U_3_land_1_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_1_lpi_1_dfm_6,
          alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_st_2, and_1308_rgt);
      IsNaN_8U_23U_2_land_2_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_4_land_2_lpi_1_dfm_6,
          alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_st_2, and_1308_rgt);
      IsNaN_8U_23U_2_land_4_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_4_land_4_lpi_1_dfm_6,
          alu_loop_op_4_FpCmp_8U_23U_false_slc_8_1_svs_st_2, and_1308_rgt);
      IsNaN_8U_23U_2_land_5_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_4_land_5_lpi_1_dfm_6,
          alu_loop_op_5_FpCmp_8U_23U_false_slc_8_svs_st_2, and_1308_rgt);
      IsNaN_8U_23U_3_land_7_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_7_lpi_1_dfm_6,
          alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_st_2, and_1308_rgt);
      IsNaN_8U_23U_2_land_9_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_4_land_9_lpi_1_dfm_6,
          alu_loop_op_9_FpCmp_8U_23U_false_slc_8_svs_st_2, and_1308_rgt);
      IsNaN_8U_23U_2_land_11_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_4_land_11_lpi_1_dfm_6,
          alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_st_2, and_1308_rgt);
      IsNaN_8U_23U_2_land_12_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_4_land_12_lpi_1_dfm_6,
          alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_st_2, and_1308_rgt);
      IsNaN_8U_23U_3_land_15_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_15_lpi_1_dfm_6,
          alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_st_2, and_1308_rgt);
      IsNaN_8U_23U_3_land_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_lpi_1_dfm_6,
          alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_st_2, and_1308_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_is_a_greater_1_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_1311_rgt | and_1313_rgt | and_1315_rgt | and_1316_rgt
        | and_1141_cse) & mux_1092_cse ) begin
      FpCmp_8U_23U_false_is_a_greater_1_lpi_1_dfm_7 <= MUX1HOT_s_1_5_2(FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_mx0w0,
          FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_mx0w1, FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_mx0w2,
          FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_mx0w3, FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w4,
          {and_1311_rgt , and_1313_rgt , and_1315_rgt , and_1316_rgt , and_1141_cse});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_3_land_2_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_3_land_5_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_3_land_9_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_3_land_11_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_3_land_12_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_3_aelse_and_1_cse ) begin
      IsNaN_8U_23U_3_land_2_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_2_lpi_1_dfm_6,
          alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2, and_1308_rgt);
      IsNaN_8U_23U_3_land_5_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_5_lpi_1_dfm_6,
          alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2, and_1308_rgt);
      IsNaN_8U_23U_3_land_9_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_9_lpi_1_dfm_6,
          alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2, and_1308_rgt);
      IsNaN_8U_23U_3_land_11_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_11_lpi_1_dfm_6,
          alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2, and_1308_rgt);
      IsNaN_8U_23U_3_land_12_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_12_lpi_1_dfm_6,
          alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2, and_1308_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_is_a_greater_2_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_1323_rgt | and_1325_rgt | and_1327_rgt | and_1328_rgt
        | and_1141_cse) & mux_1092_cse ) begin
      FpCmp_8U_23U_false_is_a_greater_2_lpi_1_dfm_7 <= MUX1HOT_s_1_5_2(FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_1_mx0w0,
          FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_1_mx0w1, FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_1_mx0w2,
          FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_1_mx0w3, FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w4,
          {and_1323_rgt , and_1325_rgt , and_1327_rgt , and_1328_rgt , and_1141_cse});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_3_land_3_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_2_land_6_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_3_land_8_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_2_land_10_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_2_land_13_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_2_land_14_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_3_aelse_and_2_cse ) begin
      IsNaN_8U_23U_3_land_3_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_3_lpi_1_dfm_6,
          alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_st_2, and_1308_rgt);
      IsNaN_8U_23U_2_land_6_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_4_land_6_lpi_1_dfm_6,
          alu_loop_op_6_FpCmp_8U_23U_false_slc_8_1_svs_st_2, and_1308_rgt);
      IsNaN_8U_23U_3_land_8_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_8_lpi_1_dfm_6,
          alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_st_2, and_1308_rgt);
      IsNaN_8U_23U_2_land_10_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_4_land_10_lpi_1_dfm_6,
          alu_loop_op_10_FpCmp_8U_23U_false_slc_8_1_svs_st_2, and_1308_rgt);
      IsNaN_8U_23U_2_land_13_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_4_land_13_lpi_1_dfm_6,
          alu_loop_op_13_FpCmp_8U_23U_false_slc_8_svs_st_2, and_1308_rgt);
      IsNaN_8U_23U_2_land_14_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_4_land_14_lpi_1_dfm_6,
          alu_loop_op_14_FpCmp_8U_23U_false_slc_8_1_svs_st_2, and_1308_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_is_a_greater_3_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_1333_rgt | and_1335_rgt | and_1337_rgt | and_1339_rgt
        | and_1308_rgt) & mux_1092_cse ) begin
      FpCmp_8U_23U_false_is_a_greater_3_lpi_1_dfm_7 <= MUX1HOT_s_1_5_2(FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_2_mx0w0,
          FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_2_mx0w1, FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_2_mx0w2,
          FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_2_mx0w3, FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w4,
          {and_1333_rgt , and_1335_rgt , and_1337_rgt , and_1339_rgt , and_1308_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_3_land_4_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_1318_cse | and_1307_cse | and_1346_rgt | and_1347_rgt)
        & mux_1092_cse ) begin
      IsNaN_8U_23U_3_land_4_lpi_1_dfm_7 <= MUX1HOT_s_1_3_2(IsNaN_8U_23U_3_land_4_lpi_1_dfm_6,
          alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0, alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm,
          {(IsNaN_8U_23U_3_aelse_or_nl) , and_1346_rgt , and_1347_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_is_a_greater_4_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_1351_rgt | and_1353_rgt | and_1355_rgt | and_1356_rgt
        | and_1141_cse) & mux_1092_cse ) begin
      FpCmp_8U_23U_false_is_a_greater_4_lpi_1_dfm_7 <= MUX1HOT_s_1_5_2(FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_3_mx0w0,
          FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_3_mx0w1, FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_3_mx0w2,
          FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_3_mx0w3, FpAdd_8U_23U_is_a_greater_lor_4_lpi_1_dfm_1_mx0w4,
          {and_1351_rgt , and_1353_rgt , and_1355_rgt , and_1356_rgt , and_1141_cse});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_is_a_greater_5_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_1364_rgt | and_1366_rgt | and_1368_rgt | and_1369_rgt
        | and_1141_cse) & mux_1092_cse ) begin
      FpCmp_8U_23U_false_is_a_greater_5_lpi_1_dfm_7 <= MUX1HOT_s_1_5_2(FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_4_mx0w0,
          FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_4_mx0w1, FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_4_mx0w2,
          FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_4_mx0w3, FpAdd_8U_23U_is_a_greater_lor_5_lpi_1_dfm_1_mx0w4,
          {and_1364_rgt , and_1366_rgt , and_1368_rgt , and_1369_rgt , and_1141_cse});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_3_land_6_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_3_land_13_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_3_aelse_and_5_cse ) begin
      IsNaN_8U_23U_3_land_6_lpi_1_dfm_7 <= MUX1HOT_s_1_3_2(IsNaN_8U_23U_3_land_6_lpi_1_dfm_6,
          alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0, alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm,
          {IsNaN_8U_23U_3_aelse_or_1_cse , and_1346_rgt , and_1347_rgt});
      IsNaN_8U_23U_3_land_13_lpi_1_dfm_7 <= MUX1HOT_s_1_3_2(IsNaN_8U_23U_3_land_13_lpi_1_dfm_6,
          alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0, alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm,
          {IsNaN_8U_23U_3_aelse_or_1_cse , and_1346_rgt , and_1347_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_is_a_greater_6_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_1380_rgt | and_1382_rgt | and_1384_rgt | and_1386_rgt
        | and_1308_rgt) & mux_1092_cse ) begin
      FpCmp_8U_23U_false_is_a_greater_6_lpi_1_dfm_7 <= MUX1HOT_s_1_5_2(FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_5_mx0w0,
          FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_5_mx0w1, FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_5_mx0w2,
          FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_5_mx0w3, FpAdd_8U_23U_is_a_greater_lor_6_lpi_1_dfm_1_mx0w4,
          {and_1380_rgt , and_1382_rgt , and_1384_rgt , and_1386_rgt , and_1308_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_is_a_greater_7_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_1391_rgt | and_1393_rgt | and_1395_rgt | and_1396_rgt
        | and_1141_cse) & mux_1092_cse ) begin
      FpCmp_8U_23U_false_is_a_greater_7_lpi_1_dfm_7 <= MUX1HOT_s_1_5_2(FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_6_mx0w0,
          FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_6_mx0w1, FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_6_mx0w2,
          FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_6_mx0w3, FpAdd_8U_23U_is_a_greater_lor_7_lpi_1_dfm_1_mx0w4,
          {and_1391_rgt , and_1393_rgt , and_1395_rgt , and_1396_rgt , and_1141_cse});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_is_a_greater_8_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_1400_rgt | and_1402_rgt | and_1404_rgt | and_1406_rgt
        | and_1308_rgt) & mux_1092_cse ) begin
      FpCmp_8U_23U_false_is_a_greater_8_lpi_1_dfm_7 <= MUX1HOT_s_1_5_2(FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_7_mx0w0,
          FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_7_mx0w1, FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_7_mx0w2,
          FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_7_mx0w3, FpAdd_8U_23U_is_a_greater_lor_8_lpi_1_dfm_1_mx0w4,
          {and_1400_rgt , and_1402_rgt , and_1404_rgt , and_1406_rgt , and_1308_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_is_a_greater_9_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_1413_rgt | and_1415_rgt | and_1417_rgt | and_1418_rgt
        | and_1141_cse) & mux_1092_cse ) begin
      FpCmp_8U_23U_false_is_a_greater_9_lpi_1_dfm_7 <= MUX1HOT_s_1_5_2(FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_8_mx0w0,
          FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_8_mx0w1, FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_8_mx0w2,
          FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_8_mx0w3, FpAdd_8U_23U_is_a_greater_lor_9_lpi_1_dfm_1_mx0w4,
          {and_1413_rgt , and_1415_rgt , and_1417_rgt , and_1418_rgt , and_1141_cse});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_3_land_10_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_3_land_14_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_3_aelse_and_9_cse ) begin
      IsNaN_8U_23U_3_land_10_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_10_lpi_1_dfm_6,
          alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2, and_1308_rgt);
      IsNaN_8U_23U_3_land_14_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_14_lpi_1_dfm_6,
          alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_2, and_1308_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_is_a_greater_10_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_1425_rgt | and_1427_rgt | and_1429_rgt | and_1431_rgt
        | and_1308_rgt) & mux_1092_cse ) begin
      FpCmp_8U_23U_false_is_a_greater_10_lpi_1_dfm_7 <= MUX1HOT_s_1_5_2(FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_9_mx0w0,
          FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_9_mx0w1, FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_9_mx0w2,
          FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_9_mx0w3, FpAdd_8U_23U_is_a_greater_lor_10_lpi_1_dfm_1_mx0w4,
          {and_1425_rgt , and_1427_rgt , and_1429_rgt , and_1431_rgt , and_1308_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_is_a_greater_11_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_1438_rgt | and_1440_rgt | and_1442_rgt | and_1444_rgt
        | and_1141_cse) & mux_1092_cse ) begin
      FpCmp_8U_23U_false_is_a_greater_11_lpi_1_dfm_7 <= MUX1HOT_s_1_5_2(FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_10_mx0w0,
          FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_10_mx0w1, FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_10_mx0w2,
          FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_10_mx0w3, FpAdd_8U_23U_is_a_greater_lor_11_lpi_1_dfm_1_mx0w4,
          {and_1438_rgt , and_1440_rgt , and_1442_rgt , and_1444_rgt , and_1141_cse});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_is_a_greater_12_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_1452_rgt | and_1454_rgt | and_1456_rgt | and_1458_rgt
        | and_1141_cse) & mux_1092_cse ) begin
      FpCmp_8U_23U_false_is_a_greater_12_lpi_1_dfm_7 <= MUX1HOT_s_1_5_2(FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_11_mx0w0,
          FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_11_mx0w1, FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_11_mx0w2,
          FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_11_mx0w3, FpAdd_8U_23U_is_a_greater_lor_12_lpi_1_dfm_1_mx0w4,
          {and_1452_rgt , and_1454_rgt , and_1456_rgt , and_1458_rgt , and_1141_cse});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_is_a_greater_13_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_1469_rgt | and_1471_rgt | and_1473_rgt | and_1475_rgt
        | and_1308_rgt) & mux_1092_cse ) begin
      FpCmp_8U_23U_false_is_a_greater_13_lpi_1_dfm_7 <= MUX1HOT_s_1_5_2(FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_12_mx0w0,
          FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_12_mx0w1, FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_12_mx0w2,
          FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_12_mx0w3, FpAdd_8U_23U_is_a_greater_lor_13_lpi_1_dfm_1_mx0w4,
          {and_1469_rgt , and_1471_rgt , and_1473_rgt , and_1475_rgt , and_1308_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_is_a_greater_14_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_1481_rgt | and_1483_rgt | and_1485_rgt | and_1487_rgt
        | and_1308_rgt) & mux_1092_cse ) begin
      FpCmp_8U_23U_false_is_a_greater_14_lpi_1_dfm_7 <= MUX1HOT_s_1_5_2(FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_13_mx0w0,
          FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_13_mx0w1, FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_13_mx0w2,
          FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_13_mx0w3, FpAdd_8U_23U_is_a_greater_lor_14_lpi_1_dfm_1_mx0w4,
          {and_1481_rgt , and_1483_rgt , and_1485_rgt , and_1487_rgt , and_1308_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_is_a_greater_15_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_1492_rgt | and_1494_rgt | and_1496_rgt | and_1498_rgt
        | and_1141_cse) & mux_1092_cse ) begin
      FpCmp_8U_23U_false_is_a_greater_15_lpi_1_dfm_7 <= MUX1HOT_s_1_5_2(FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_14_mx0w0,
          FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_14_mx0w1, FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_14_mx0w2,
          FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_14_mx0w3, FpAdd_8U_23U_is_a_greater_lor_15_lpi_1_dfm_1_mx0w4,
          {and_1492_rgt , and_1494_rgt , and_1496_rgt , and_1498_rgt , and_1141_cse});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_is_a_greater_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_1503_rgt | and_1505_rgt | and_1507_rgt | and_1508_rgt
        | and_1141_cse) & mux_1092_cse ) begin
      FpCmp_8U_23U_false_is_a_greater_lpi_1_dfm_7 <= MUX1HOT_s_1_5_2(FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_15_mx0w0,
          FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_15_mx0w1, FpCmp_8U_23U_true_else_1_FpCmp_8U_23U_true_else_1_and_15_mx0w2,
          FpCmp_8U_23U_true_if_1_FpCmp_8U_23U_true_if_1_or_15_mx0w3, FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w4,
          {and_1503_rgt , and_1505_rgt , and_1507_rgt , and_1508_rgt , and_1141_cse});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_itm_2 <= 1'b0;
      alu_loop_op_else_else_if_mux_2_itm_2 <= 1'b0;
      alu_loop_op_else_else_if_mux_1_itm_2 <= 30'b0;
    end
    else if ( alu_loop_op_else_else_if_and_144_cse ) begin
      alu_loop_op_else_else_if_mux_itm_2 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[31]),
          IntShiftLeft_16U_6U_32U_return_31_1_sva_2, alu_loop_op_else_else_if_mux_itm,
          alu_loop_op_else_if_mux_itm, {and_dcpl_1044 , and_dcpl_1046 , and_dcpl_1048
          , and_dcpl_1050});
      alu_loop_op_else_else_if_mux_2_itm_2 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[0]),
          IntShiftLeft_16U_6U_32U_return_0_1_sva_2, alu_loop_op_else_else_if_mux_2_itm,
          alu_loop_op_else_if_mux_2_itm, {and_dcpl_1044 , and_dcpl_1046 , and_dcpl_1048
          , and_dcpl_1050});
      alu_loop_op_else_else_if_mux_1_itm_2 <= MUX1HOT_v_30_4_2((AluIn_data_sva_501[30:1]),
          IntShiftLeft_16U_6U_32U_return_30_1_1_sva_2, alu_loop_op_else_else_if_mux_1_itm,
          alu_loop_op_else_if_mux_1_itm, {and_dcpl_1044 , and_dcpl_1046 , and_dcpl_1048
          , and_dcpl_1050});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_3_itm_2 <= 1'b0;
      alu_loop_op_else_else_if_mux_5_itm_2 <= 1'b0;
      alu_loop_op_else_else_if_mux_4_itm_2 <= 30'b0;
    end
    else if ( alu_loop_op_else_else_if_and_147_cse ) begin
      alu_loop_op_else_else_if_mux_3_itm_2 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[63]),
          IntShiftLeft_16U_6U_32U_return_31_2_sva_2, alu_loop_op_else_else_if_mux_3_itm,
          alu_loop_op_else_if_mux_3_itm, {and_dcpl_1052 , and_dcpl_1054 , and_dcpl_1048
          , and_dcpl_1050});
      alu_loop_op_else_else_if_mux_5_itm_2 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[32]),
          IntShiftLeft_16U_6U_32U_return_0_2_sva_2, alu_loop_op_else_else_if_mux_5_itm,
          alu_loop_op_else_if_mux_5_itm, {and_dcpl_1052 , and_dcpl_1054 , and_dcpl_1048
          , and_dcpl_1050});
      alu_loop_op_else_else_if_mux_4_itm_2 <= MUX1HOT_v_30_4_2((AluIn_data_sva_501[62:33]),
          IntShiftLeft_16U_6U_32U_return_30_1_2_sva_2, alu_loop_op_else_else_if_mux_4_itm,
          alu_loop_op_else_if_mux_4_itm, {and_dcpl_1052 , and_dcpl_1054 , and_dcpl_1048
          , and_dcpl_1050});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_9_itm_2 <= 1'b0;
      alu_loop_op_else_else_if_mux_11_itm_2 <= 1'b0;
      alu_loop_op_else_else_if_mux_10_itm_2 <= 30'b0;
    end
    else if ( alu_loop_op_else_else_if_and_150_cse ) begin
      alu_loop_op_else_else_if_mux_9_itm_2 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[127]),
          IntShiftLeft_16U_6U_32U_return_31_4_sva_2, alu_loop_op_else_else_if_mux_9_itm,
          alu_loop_op_else_if_mux_9_itm, {and_dcpl_1060 , and_dcpl_1062 , and_dcpl_1048
          , and_dcpl_1050});
      alu_loop_op_else_else_if_mux_11_itm_2 <= MUX1HOT_s_1_4_2((AluIn_data_sva_501[96]),
          IntShiftLeft_16U_6U_32U_return_0_4_sva_2, alu_loop_op_else_else_if_mux_11_itm,
          alu_loop_op_else_if_mux_11_itm, {and_dcpl_1060 , and_dcpl_1062 , and_dcpl_1048
          , and_dcpl_1050});
      alu_loop_op_else_else_if_mux_10_itm_2 <= MUX1HOT_v_30_4_2((AluIn_data_sva_501[126:97]),
          IntShiftLeft_16U_6U_32U_return_30_1_4_sva_2, alu_loop_op_else_else_if_mux_10_itm,
          alu_loop_op_else_if_mux_10_itm, {and_dcpl_1060 , and_dcpl_1062 , and_dcpl_1048
          , and_dcpl_1050});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_14_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_1_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_65_mx0w1,
          or_tmp_3190);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_1_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_64_mx0w1,
          or_tmp_3190);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_12_10 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_12_10 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_12_10 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_12_10 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_12_10 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_12_10 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_12_10 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_12_10 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_12_10 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_12_10 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_12_10 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_12_10 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_12_10 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_12_10 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_12_10 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_12_10 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3 <= 4'b0;
      alu_nan_to_zero_op_sign_1_lpi_1_dfm <= 1'b0;
      alu_nan_to_zero_op_sign_2_lpi_1_dfm <= 1'b0;
      alu_nan_to_zero_op_sign_3_lpi_1_dfm <= 1'b0;
      alu_nan_to_zero_op_sign_4_lpi_1_dfm <= 1'b0;
      alu_nan_to_zero_op_sign_5_lpi_1_dfm <= 1'b0;
      alu_nan_to_zero_op_sign_6_lpi_1_dfm <= 1'b0;
      alu_nan_to_zero_op_sign_7_lpi_1_dfm <= 1'b0;
      alu_nan_to_zero_op_sign_8_lpi_1_dfm <= 1'b0;
      alu_nan_to_zero_op_sign_9_lpi_1_dfm <= 1'b0;
      alu_nan_to_zero_op_sign_10_lpi_1_dfm <= 1'b0;
      alu_nan_to_zero_op_sign_11_lpi_1_dfm <= 1'b0;
      alu_nan_to_zero_op_sign_12_lpi_1_dfm <= 1'b0;
      alu_nan_to_zero_op_sign_13_lpi_1_dfm <= 1'b0;
      alu_nan_to_zero_op_sign_14_lpi_1_dfm <= 1'b0;
      alu_nan_to_zero_op_sign_15_lpi_1_dfm <= 1'b0;
      alu_nan_to_zero_op_sign_lpi_1_dfm <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_15_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_12_10_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_12_10_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_12_10_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_12_10_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_12_10_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_12_10_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_12_10_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_12_10_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_12_10_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_12_10_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_12_10_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_12_10_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_12_10_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_12_10_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_12_10_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_12_10_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w0;
      alu_nan_to_zero_op_sign_1_lpi_1_dfm <= alu_nan_to_zero_op_sign_1_lpi_1_dfm_mx0w0;
      alu_nan_to_zero_op_sign_2_lpi_1_dfm <= alu_nan_to_zero_op_sign_2_lpi_1_dfm_mx0w0;
      alu_nan_to_zero_op_sign_3_lpi_1_dfm <= alu_nan_to_zero_op_sign_3_lpi_1_dfm_mx0w0;
      alu_nan_to_zero_op_sign_4_lpi_1_dfm <= alu_nan_to_zero_op_sign_4_lpi_1_dfm_mx0w0;
      alu_nan_to_zero_op_sign_5_lpi_1_dfm <= alu_nan_to_zero_op_sign_5_lpi_1_dfm_mx0w0;
      alu_nan_to_zero_op_sign_6_lpi_1_dfm <= alu_nan_to_zero_op_sign_6_lpi_1_dfm_mx0w0;
      alu_nan_to_zero_op_sign_7_lpi_1_dfm <= alu_nan_to_zero_op_sign_7_lpi_1_dfm_mx0w0;
      alu_nan_to_zero_op_sign_8_lpi_1_dfm <= alu_nan_to_zero_op_sign_8_lpi_1_dfm_mx0w0;
      alu_nan_to_zero_op_sign_9_lpi_1_dfm <= alu_nan_to_zero_op_sign_9_lpi_1_dfm_mx0w0;
      alu_nan_to_zero_op_sign_10_lpi_1_dfm <= alu_nan_to_zero_op_sign_10_lpi_1_dfm_mx0w0;
      alu_nan_to_zero_op_sign_11_lpi_1_dfm <= alu_nan_to_zero_op_sign_11_lpi_1_dfm_mx0w0;
      alu_nan_to_zero_op_sign_12_lpi_1_dfm <= alu_nan_to_zero_op_sign_12_lpi_1_dfm_mx0w0;
      alu_nan_to_zero_op_sign_13_lpi_1_dfm <= alu_nan_to_zero_op_sign_13_lpi_1_dfm_mx0w0;
      alu_nan_to_zero_op_sign_14_lpi_1_dfm <= alu_nan_to_zero_op_sign_14_lpi_1_dfm_mx0w0;
      alu_nan_to_zero_op_sign_15_lpi_1_dfm <= alu_nan_to_zero_op_sign_15_lpi_1_dfm_mx0w0;
      alu_nan_to_zero_op_sign_lpi_1_dfm <= alu_nan_to_zero_op_sign_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_393 | (cfg_alu_algo_1_sva_st_92[0]) | FpCmp_8U_23U_true_if_acc_16_itm_8_1
        | (~ (cfg_alu_algo_1_sva_st_92[1])))) ) begin
      alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_svs <= alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_FpAdd_8U_23U_is_a_greater_slc_8_svs <= 1'b0;
      alu_loop_op_10_FpAdd_8U_23U_is_a_greater_slc_8_1_svs <= 1'b0;
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= 1'b0;
      alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st
          <= 1'b0;
      alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= 1'b0;
      alu_loop_op_10_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st
          <= 1'b0;
    end
    else if ( FpAdd_8U_23U_is_a_greater_and_cse ) begin
      alu_loop_op_1_FpAdd_8U_23U_is_a_greater_slc_8_svs <= FpCmp_8U_23U_true_if_acc_16_itm_8_1;
      alu_loop_op_10_FpAdd_8U_23U_is_a_greater_slc_8_1_svs <= FpCmp_8U_23U_true_if_acc_34_itm_8_1;
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
      alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st
          <= alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0;
      alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
      alu_loop_op_10_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st
          <= alu_loop_op_10_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_FpCmp_8U_23U_true_slc_8_svs_st <= 1'b0;
      alu_loop_op_2_FpCmp_8U_23U_true_slc_8_1_svs_st <= 1'b0;
      alu_loop_op_3_FpCmp_8U_23U_true_slc_8_svs_st <= 1'b0;
      alu_loop_op_4_FpCmp_8U_23U_true_slc_8_1_svs_st <= 1'b0;
      alu_loop_op_5_FpCmp_8U_23U_true_slc_8_svs_st <= 1'b0;
      alu_loop_op_6_FpCmp_8U_23U_true_slc_8_1_svs_st <= 1'b0;
      alu_loop_op_7_FpCmp_8U_23U_true_slc_8_svs_st <= 1'b0;
      alu_loop_op_9_FpCmp_8U_23U_true_slc_8_svs_st <= 1'b0;
      alu_loop_op_10_FpCmp_8U_23U_true_slc_8_1_svs_st <= 1'b0;
      alu_loop_op_11_FpCmp_8U_23U_true_slc_8_svs_st <= 1'b0;
      alu_loop_op_13_FpCmp_8U_23U_true_slc_8_svs_st <= 1'b0;
      alu_loop_op_14_FpCmp_8U_23U_true_slc_8_1_svs_st <= 1'b0;
      alu_loop_op_15_FpCmp_8U_23U_true_slc_8_svs_st <= 1'b0;
      alu_loop_op_16_FpCmp_8U_23U_true_slc_8_1_svs_st <= 1'b0;
    end
    else if ( FpCmp_8U_23U_true_if_and_cse ) begin
      alu_loop_op_1_FpCmp_8U_23U_true_slc_8_svs_st <= FpCmp_8U_23U_true_if_acc_16_itm_8_1;
      alu_loop_op_2_FpCmp_8U_23U_true_slc_8_1_svs_st <= FpCmp_8U_23U_true_if_acc_18_itm_8_1;
      alu_loop_op_3_FpCmp_8U_23U_true_slc_8_svs_st <= FpCmp_8U_23U_true_if_acc_20_itm_8_1;
      alu_loop_op_4_FpCmp_8U_23U_true_slc_8_1_svs_st <= FpCmp_8U_23U_true_if_acc_22_itm_8_1;
      alu_loop_op_5_FpCmp_8U_23U_true_slc_8_svs_st <= FpCmp_8U_23U_true_if_acc_24_itm_8_1;
      alu_loop_op_6_FpCmp_8U_23U_true_slc_8_1_svs_st <= FpCmp_8U_23U_true_if_acc_26_itm_8_1;
      alu_loop_op_7_FpCmp_8U_23U_true_slc_8_svs_st <= FpCmp_8U_23U_true_if_acc_28_itm_8_1;
      alu_loop_op_9_FpCmp_8U_23U_true_slc_8_svs_st <= FpCmp_8U_23U_true_if_acc_32_itm_8_1;
      alu_loop_op_10_FpCmp_8U_23U_true_slc_8_1_svs_st <= FpCmp_8U_23U_true_if_acc_34_itm_8_1;
      alu_loop_op_11_FpCmp_8U_23U_true_slc_8_svs_st <= FpCmp_8U_23U_true_if_acc_36_itm_8_1;
      alu_loop_op_13_FpCmp_8U_23U_true_slc_8_svs_st <= FpCmp_8U_23U_true_if_acc_40_itm_8_1;
      alu_loop_op_14_FpCmp_8U_23U_true_slc_8_1_svs_st <= FpCmp_8U_23U_true_if_acc_42_itm_8_1;
      alu_loop_op_15_FpCmp_8U_23U_true_slc_8_svs_st <= FpCmp_8U_23U_true_if_acc_44_itm_8_1;
      alu_loop_op_16_FpCmp_8U_23U_true_slc_8_1_svs_st <= FpCmp_8U_23U_true_if_acc_46_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_st <= 1'b0;
      alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_st <= 1'b0;
      alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_st <= 1'b0;
      alu_loop_op_4_FpCmp_8U_23U_false_slc_8_1_svs_st <= 1'b0;
      alu_loop_op_5_FpCmp_8U_23U_false_slc_8_svs_st <= 1'b0;
      alu_loop_op_6_FpCmp_8U_23U_false_slc_8_1_svs_st <= 1'b0;
      alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_st <= 1'b0;
      alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_st <= 1'b0;
      alu_loop_op_9_FpCmp_8U_23U_false_slc_8_svs_st <= 1'b0;
      alu_loop_op_10_FpCmp_8U_23U_false_slc_8_1_svs_st <= 1'b0;
      alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_st <= 1'b0;
      alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_st <= 1'b0;
      alu_loop_op_13_FpCmp_8U_23U_false_slc_8_svs_st <= 1'b0;
      alu_loop_op_14_FpCmp_8U_23U_false_slc_8_1_svs_st <= 1'b0;
      alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_st <= 1'b0;
      alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_st <= 1'b0;
    end
    else if ( FpCmp_8U_23U_false_if_and_cse ) begin
      alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_st <= FpCmp_8U_23U_true_if_acc_16_itm_8_1;
      alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_st <= FpCmp_8U_23U_true_if_acc_18_itm_8_1;
      alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_st <= FpCmp_8U_23U_true_if_acc_20_itm_8_1;
      alu_loop_op_4_FpCmp_8U_23U_false_slc_8_1_svs_st <= FpCmp_8U_23U_true_if_acc_22_itm_8_1;
      alu_loop_op_5_FpCmp_8U_23U_false_slc_8_svs_st <= FpCmp_8U_23U_true_if_acc_24_itm_8_1;
      alu_loop_op_6_FpCmp_8U_23U_false_slc_8_1_svs_st <= FpCmp_8U_23U_true_if_acc_26_itm_8_1;
      alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_st <= FpCmp_8U_23U_true_if_acc_28_itm_8_1;
      alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_st <= FpCmp_8U_23U_true_if_acc_30_itm_8_1;
      alu_loop_op_9_FpCmp_8U_23U_false_slc_8_svs_st <= FpCmp_8U_23U_true_if_acc_32_itm_8_1;
      alu_loop_op_10_FpCmp_8U_23U_false_slc_8_1_svs_st <= FpCmp_8U_23U_true_if_acc_34_itm_8_1;
      alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_st <= FpCmp_8U_23U_true_if_acc_36_itm_8_1;
      alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_st <= FpCmp_8U_23U_true_if_acc_38_itm_8_1;
      alu_loop_op_13_FpCmp_8U_23U_false_slc_8_svs_st <= FpCmp_8U_23U_true_if_acc_40_itm_8_1;
      alu_loop_op_14_FpCmp_8U_23U_false_slc_8_1_svs_st <= FpCmp_8U_23U_true_if_acc_42_itm_8_1;
      alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_st <= FpCmp_8U_23U_true_if_acc_44_itm_8_1;
      alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_st <= FpCmp_8U_23U_true_if_acc_46_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_17_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_2_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_67_mx0w1,
          or_tmp_3201);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_2_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_66_mx0w1,
          or_tmp_3201);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_st <= 1'b0;
    end
    else if ( IsNaN_8U_23U_2_aelse_and_cse & (~ or_dcpl_414) & (~ (mux_1359_nl))
        ) begin
      alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_st <= alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_13 | (cfg_precision[0]) | FpCmp_8U_23U_true_if_acc_18_itm_8_1
        | or_dcpl_413)) ) begin
      alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs <= alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_alu_loop_op_2_FpAdd_8U_23U_is_a_greater_slc_8_1_svs_cse <= 1'b0;
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= 1'b0;
      alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st
          <= 1'b0;
    end
    else if ( FpAdd_8U_23U_is_a_greater_and_1_cse ) begin
      reg_alu_loop_op_2_FpAdd_8U_23U_is_a_greater_slc_8_1_svs_cse <= FpCmp_8U_23U_true_if_acc_18_itm_8_1;
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
      alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st
          <= alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_20_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_3_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_69_mx0w1,
          or_tmp_3212);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_3_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_68_mx0w1,
          or_tmp_3212);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_13 | (cfg_precision[0]) | FpCmp_8U_23U_true_if_acc_20_itm_8_1
        | or_dcpl_413)) ) begin
      alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_svs <= alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_3_FpAdd_8U_23U_is_a_greater_slc_8_svs <= 1'b0;
      alu_loop_op_4_FpAdd_8U_23U_is_a_greater_slc_8_1_svs <= 1'b0;
      alu_loop_op_5_FpAdd_8U_23U_is_a_greater_slc_8_svs <= 1'b0;
      alu_loop_op_6_FpAdd_8U_23U_is_a_greater_slc_8_1_svs <= 1'b0;
      alu_loop_op_7_FpAdd_8U_23U_is_a_greater_slc_8_svs <= 1'b0;
      alu_loop_op_9_FpAdd_8U_23U_is_a_greater_slc_8_svs <= 1'b0;
      alu_loop_op_11_FpAdd_8U_23U_is_a_greater_slc_8_svs <= 1'b0;
      alu_loop_op_13_FpAdd_8U_23U_is_a_greater_slc_8_svs <= 1'b0;
      alu_loop_op_14_FpAdd_8U_23U_is_a_greater_slc_8_1_svs <= 1'b0;
      alu_loop_op_15_FpAdd_8U_23U_is_a_greater_slc_8_svs <= 1'b0;
      alu_loop_op_16_FpAdd_8U_23U_is_a_greater_slc_8_1_svs <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st
          <= 1'b0;
      alu_loop_op_4_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm <= 1'b0;
      alu_loop_op_4_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm <= 1'b0;
      alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st
          <= 1'b0;
      alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= 1'b0;
      alu_loop_op_5_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st
          <= 1'b0;
      alu_loop_op_6_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm <= 1'b0;
      alu_loop_op_6_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm <= 1'b0;
      alu_loop_op_6_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st
          <= 1'b0;
      alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= 1'b0;
      alu_loop_op_7_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st
          <= 1'b0;
      alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= 1'b0;
      alu_loop_op_9_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st
          <= 1'b0;
      alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= 1'b0;
      alu_loop_op_11_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st
          <= 1'b0;
      alu_loop_op_13_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_itm <= 1'b0;
      alu_loop_op_13_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_itm <= 1'b0;
      alu_loop_op_13_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st
          <= 1'b0;
      alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= 1'b0;
      alu_loop_op_14_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st
          <= 1'b0;
      alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= 1'b0;
      alu_loop_op_15_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st
          <= 1'b0;
      alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= 1'b0;
      alu_loop_op_16_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st
          <= 1'b0;
    end
    else if ( FpAdd_8U_23U_is_a_greater_and_3_cse ) begin
      alu_loop_op_3_FpAdd_8U_23U_is_a_greater_slc_8_svs <= FpCmp_8U_23U_true_if_acc_20_itm_8_1;
      alu_loop_op_4_FpAdd_8U_23U_is_a_greater_slc_8_1_svs <= FpCmp_8U_23U_true_if_acc_22_itm_8_1;
      alu_loop_op_5_FpAdd_8U_23U_is_a_greater_slc_8_svs <= FpCmp_8U_23U_true_if_acc_24_itm_8_1;
      alu_loop_op_6_FpAdd_8U_23U_is_a_greater_slc_8_1_svs <= FpCmp_8U_23U_true_if_acc_26_itm_8_1;
      alu_loop_op_7_FpAdd_8U_23U_is_a_greater_slc_8_svs <= FpCmp_8U_23U_true_if_acc_28_itm_8_1;
      alu_loop_op_9_FpAdd_8U_23U_is_a_greater_slc_8_svs <= FpCmp_8U_23U_true_if_acc_32_itm_8_1;
      alu_loop_op_11_FpAdd_8U_23U_is_a_greater_slc_8_svs <= FpCmp_8U_23U_true_if_acc_36_itm_8_1;
      alu_loop_op_13_FpAdd_8U_23U_is_a_greater_slc_8_svs <= FpCmp_8U_23U_true_if_acc_40_itm_8_1;
      alu_loop_op_14_FpAdd_8U_23U_is_a_greater_slc_8_1_svs <= FpCmp_8U_23U_true_if_acc_42_itm_8_1;
      alu_loop_op_15_FpAdd_8U_23U_is_a_greater_slc_8_svs <= FpCmp_8U_23U_true_if_acc_44_itm_8_1;
      alu_loop_op_16_FpAdd_8U_23U_is_a_greater_slc_8_1_svs <= FpCmp_8U_23U_true_if_acc_46_itm_8_1;
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
      alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st
          <= alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0;
      alu_loop_op_4_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm <= alu_loop_op_4_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm_mx0w0;
      alu_loop_op_4_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm <= alu_loop_op_4_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm_mx0w0;
      alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st
          <= alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0;
      alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
      alu_loop_op_5_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st
          <= alu_loop_op_5_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0;
      alu_loop_op_6_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm <= alu_loop_op_6_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_itm_mx0w0;
      alu_loop_op_6_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm <= alu_loop_op_6_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_1_itm_mx0w0;
      alu_loop_op_6_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st
          <= alu_loop_op_6_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0;
      alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
      alu_loop_op_7_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st
          <= alu_loop_op_7_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0;
      alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
      alu_loop_op_9_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st
          <= alu_loop_op_9_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0;
      alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
      alu_loop_op_11_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st
          <= alu_loop_op_11_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0;
      alu_loop_op_13_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_itm <= alu_loop_op_13_IsZero_8U_23U_1_IsZero_8U_23U_1_nor_itm_mx0w0;
      alu_loop_op_13_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_itm <= alu_loop_op_13_IsZero_8U_23U_1_aif_IsZero_8U_23U_1_aelse_nor_itm_mx0w0;
      alu_loop_op_13_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st
          <= alu_loop_op_13_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0;
      alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
      alu_loop_op_14_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st
          <= alu_loop_op_14_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0;
      alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
      alu_loop_op_15_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st
          <= alu_loop_op_15_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0;
      alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
      alu_loop_op_16_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st
          <= alu_loop_op_16_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_23_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_4_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_71_mx0w1,
          or_tmp_3223);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_4_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_70_mx0w1,
          or_tmp_3223);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_13 | (cfg_precision[0]) | FpCmp_8U_23U_true_if_acc_22_itm_8_1
        | or_dcpl_413)) ) begin
      alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs <= alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_26_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_5_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_73_mx0w1,
          or_tmp_3234);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_5_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_72_mx0w1,
          or_tmp_3234);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_5_FpAdd_8U_23U_is_a_greater_oif_equal_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_13 | (cfg_precision[0]) | FpCmp_8U_23U_true_if_acc_24_itm_8_1
        | or_dcpl_413)) ) begin
      alu_loop_op_5_FpAdd_8U_23U_is_a_greater_oif_equal_svs <= alu_loop_op_5_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_29_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_6_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_75_mx0w1,
          or_tmp_3245);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_6_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_74_mx0w1,
          or_tmp_3245);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_6_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_13 | (cfg_precision[0]) | FpCmp_8U_23U_true_if_acc_26_itm_8_1
        | or_dcpl_413)) ) begin
      alu_loop_op_6_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs <= alu_loop_op_6_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_32_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_7_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_77_mx0w1,
          or_tmp_3256);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_7_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_76_mx0w1,
          or_tmp_3256);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_7_FpAdd_8U_23U_is_a_greater_oif_equal_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_13 | (cfg_precision[0]) | FpCmp_8U_23U_true_if_acc_28_itm_8_1
        | or_dcpl_413)) ) begin
      alu_loop_op_7_FpAdd_8U_23U_is_a_greater_oif_equal_svs <= alu_loop_op_7_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_35_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_8_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_79_mx0w1,
          or_tmp_3267);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_8_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_78_mx0w1,
          or_tmp_3267);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_8_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_13 | (cfg_precision[0]) | FpCmp_8U_23U_true_if_acc_30_itm_8_1
        | or_dcpl_520)) ) begin
      alu_loop_op_8_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs <= alu_loop_op_8_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_8_FpAdd_8U_23U_is_a_greater_slc_8_1_svs <= 1'b0;
      alu_loop_op_12_FpAdd_8U_23U_is_a_greater_slc_8_1_svs <= 1'b0;
      alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= 1'b0;
      alu_loop_op_8_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st
          <= 1'b0;
      alu_loop_op_12_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st
          <= 1'b0;
      alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= 1'b0;
    end
    else if ( FpAdd_8U_23U_is_a_greater_and_8_cse ) begin
      alu_loop_op_8_FpAdd_8U_23U_is_a_greater_slc_8_1_svs <= FpCmp_8U_23U_true_if_acc_30_itm_8_1;
      alu_loop_op_12_FpAdd_8U_23U_is_a_greater_slc_8_1_svs <= FpCmp_8U_23U_true_if_acc_38_itm_8_1;
      alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
      alu_loop_op_8_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st
          <= alu_loop_op_8_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0;
      alu_loop_op_12_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st
          <= alu_loop_op_12_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0;
      alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm <= alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_1_nand_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_8_FpCmp_8U_23U_true_slc_8_1_svs_st <= 1'b0;
      alu_loop_op_12_FpCmp_8U_23U_true_slc_8_1_svs_st <= 1'b0;
    end
    else if ( FpCmp_8U_23U_true_if_and_7_cse ) begin
      alu_loop_op_8_FpCmp_8U_23U_true_slc_8_1_svs_st <= FpCmp_8U_23U_true_if_acc_30_itm_8_1;
      alu_loop_op_12_FpCmp_8U_23U_true_slc_8_1_svs_st <= FpCmp_8U_23U_true_if_acc_38_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_38_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_9_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_81_mx0w1,
          or_tmp_3278);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_9_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_80_mx0w1,
          or_tmp_3278);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_9_FpAdd_8U_23U_is_a_greater_oif_equal_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_13 | (cfg_precision[0]) | FpCmp_8U_23U_true_if_acc_32_itm_8_1
        | or_dcpl_413)) ) begin
      alu_loop_op_9_FpAdd_8U_23U_is_a_greater_oif_equal_svs <= alu_loop_op_9_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_41_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_10_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_83_mx0w1,
          or_tmp_3289);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_10_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_82_mx0w1,
          or_tmp_3289);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_10_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_393 | (cfg_alu_algo_1_sva_st_92[0]) | FpCmp_8U_23U_true_if_acc_34_itm_8_1
        | (~ (cfg_alu_algo_1_sva_st_92[1])))) ) begin
      alu_loop_op_10_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs <= alu_loop_op_10_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_44_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_11_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_85_mx0w1,
          or_tmp_3300);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_11_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_84_mx0w1,
          or_tmp_3300);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_11_FpAdd_8U_23U_is_a_greater_oif_equal_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_13 | (cfg_precision[0]) | FpCmp_8U_23U_true_if_acc_36_itm_8_1
        | or_dcpl_413)) ) begin
      alu_loop_op_11_FpAdd_8U_23U_is_a_greater_oif_equal_svs <= alu_loop_op_11_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_47_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_12_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_87_mx0w1,
          or_tmp_3311);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_12_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_86_mx0w1,
          or_tmp_3311);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_12_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_13 | (cfg_precision[0]) | FpCmp_8U_23U_true_if_acc_38_itm_8_1
        | or_dcpl_520)) ) begin
      alu_loop_op_12_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs <= alu_loop_op_12_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_50_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_13_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_89_mx0w1,
          or_tmp_3322);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_13_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_88_mx0w1,
          or_tmp_3322);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_13_FpAdd_8U_23U_is_a_greater_oif_equal_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_13 | (cfg_precision[0]) | FpCmp_8U_23U_true_if_acc_40_itm_8_1
        | or_dcpl_413)) ) begin
      alu_loop_op_13_FpAdd_8U_23U_is_a_greater_oif_equal_svs <= alu_loop_op_13_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_53_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_14_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_91_mx0w1,
          or_tmp_3333);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_14_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_90_mx0w1,
          or_tmp_3333);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_14_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_13 | (cfg_precision[0]) | FpCmp_8U_23U_true_if_acc_42_itm_8_1
        | or_dcpl_413)) ) begin
      alu_loop_op_14_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs <= alu_loop_op_14_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_56_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_15_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_93_mx0w1,
          or_tmp_3344);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_15_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_92_mx0w1,
          or_tmp_3344);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_15_FpAdd_8U_23U_is_a_greater_oif_equal_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_13 | (cfg_precision[0]) | FpCmp_8U_23U_true_if_acc_44_itm_8_1
        | or_dcpl_413)) ) begin
      alu_loop_op_15_FpAdd_8U_23U_is_a_greater_oif_equal_svs <= alu_loop_op_15_FpAdd_8U_23U_is_a_greater_oif_equal_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_59_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_95_mx0w1,
          or_tmp_3355);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_94_mx0w1,
          or_tmp_3355);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_16_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_13 | (cfg_precision[0]) | FpCmp_8U_23U_true_if_acc_46_itm_8_1
        | or_dcpl_413)) ) begin
      alu_loop_op_16_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs <= alu_loop_op_16_FpAdd_8U_23U_is_a_greater_oif_equal_1_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_2_land_1_lpi_1_dfm_st <= 1'b0;
      IsNaN_8U_23U_2_land_2_lpi_1_dfm_st <= 1'b0;
      IsNaN_8U_23U_2_land_3_lpi_1_dfm_st <= 1'b0;
      IsNaN_8U_23U_2_land_4_lpi_1_dfm_st <= 1'b0;
      IsNaN_8U_23U_2_land_5_lpi_1_dfm_st <= 1'b0;
      IsNaN_8U_23U_2_land_6_lpi_1_dfm_st <= 1'b0;
      IsNaN_8U_23U_2_land_7_lpi_1_dfm_st <= 1'b0;
      IsNaN_8U_23U_2_land_8_lpi_1_dfm_st <= 1'b0;
      IsNaN_8U_23U_2_land_9_lpi_1_dfm_st <= 1'b0;
      IsNaN_8U_23U_2_land_10_lpi_1_dfm_st <= 1'b0;
      IsNaN_8U_23U_2_land_11_lpi_1_dfm_st <= 1'b0;
      IsNaN_8U_23U_2_land_12_lpi_1_dfm_st <= 1'b0;
      IsNaN_8U_23U_2_land_13_lpi_1_dfm_st <= 1'b0;
      IsNaN_8U_23U_2_land_14_lpi_1_dfm_st <= 1'b0;
      IsNaN_8U_23U_2_land_15_lpi_1_dfm_st <= 1'b0;
      IsNaN_8U_23U_2_land_lpi_1_dfm_st <= 1'b0;
    end
    else if ( IsNaN_8U_23U_2_aelse_and_74_cse ) begin
      IsNaN_8U_23U_2_land_1_lpi_1_dfm_st <= IsNaN_8U_23U_2_land_1_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_2_land_2_lpi_1_dfm_st <= IsNaN_8U_23U_2_land_2_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_2_land_3_lpi_1_dfm_st <= IsNaN_8U_23U_2_land_3_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_2_land_4_lpi_1_dfm_st <= IsNaN_8U_23U_2_land_4_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_2_land_5_lpi_1_dfm_st <= IsNaN_8U_23U_2_land_5_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_2_land_6_lpi_1_dfm_st <= IsNaN_8U_23U_2_land_6_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_2_land_7_lpi_1_dfm_st <= IsNaN_8U_23U_2_land_7_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_2_land_8_lpi_1_dfm_st <= IsNaN_8U_23U_2_land_8_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_2_land_9_lpi_1_dfm_st <= IsNaN_8U_23U_2_land_9_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_2_land_10_lpi_1_dfm_st <= IsNaN_8U_23U_2_land_10_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_2_land_11_lpi_1_dfm_st <= IsNaN_8U_23U_2_land_11_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_2_land_12_lpi_1_dfm_st <= IsNaN_8U_23U_2_land_12_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_2_land_13_lpi_1_dfm_st <= IsNaN_8U_23U_2_land_13_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_2_land_14_lpi_1_dfm_st <= IsNaN_8U_23U_2_land_14_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_2_land_15_lpi_1_dfm_st <= IsNaN_8U_23U_2_land_15_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_2_land_lpi_1_dfm_st <= IsNaN_8U_23U_2_land_lpi_1_dfm_mx1w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_algo_1_sva_st_15 <= 2'b0;
    end
    else if ( core_wen & (~(or_dcpl_675 | (fsm_output[0]))) ) begin
      cfg_alu_algo_1_sva_st_15 <= cfg_alu_algo_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_src_1_sva_st <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_3 | (fsm_output[0]))) ) begin
      cfg_alu_src_1_sva_st <= cfg_alu_src_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_2_lpi_1_dfm_7_4 <= 4'b0;
      FpAdd_8U_23U_qr_2_lpi_1_dfm_3_0 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_144_cse ) begin
      FpAdd_8U_23U_qr_2_lpi_1_dfm_7_4 <= MUX_v_4_2_2((AluIn_data_sva_501[30:27]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_9, and_dcpl_1335);
      FpAdd_8U_23U_qr_2_lpi_1_dfm_3_0 <= MUX_v_4_2_2((AluIn_data_sva_501[26:23]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_9, and_dcpl_1335);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_3_lpi_1_dfm_7_4 <= 4'b0;
      FpAdd_8U_23U_qr_3_lpi_1_dfm_3_0 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_146_cse ) begin
      FpAdd_8U_23U_qr_3_lpi_1_dfm_7_4 <= MUX_v_4_2_2((AluIn_data_sva_501[62:59]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_9, and_dcpl_1341);
      FpAdd_8U_23U_qr_3_lpi_1_dfm_3_0 <= MUX_v_4_2_2((AluIn_data_sva_501[58:55]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_9, and_dcpl_1341);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_4_lpi_1_dfm_7_4 <= 4'b0;
      FpAdd_8U_23U_qr_4_lpi_1_dfm_3_0 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_148_cse ) begin
      FpAdd_8U_23U_qr_4_lpi_1_dfm_7_4 <= MUX_v_4_2_2((AluIn_data_sva_501[94:91]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_9, and_dcpl_1347);
      FpAdd_8U_23U_qr_4_lpi_1_dfm_3_0 <= MUX_v_4_2_2((AluIn_data_sva_501[90:87]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_9, and_dcpl_1347);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_5_lpi_1_dfm_7_4 <= 4'b0;
      FpAdd_8U_23U_qr_5_lpi_1_dfm_3_0 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_150_cse ) begin
      FpAdd_8U_23U_qr_5_lpi_1_dfm_7_4 <= MUX_v_4_2_2((AluIn_data_sva_501[126:123]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_9, and_dcpl_1353);
      FpAdd_8U_23U_qr_5_lpi_1_dfm_3_0 <= MUX_v_4_2_2((AluIn_data_sva_501[122:119]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_9, and_dcpl_1353);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_6_lpi_1_dfm_7_4 <= 4'b0;
      FpAdd_8U_23U_qr_6_lpi_1_dfm_3_0 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_152_cse ) begin
      FpAdd_8U_23U_qr_6_lpi_1_dfm_7_4 <= MUX_v_4_2_2((AluIn_data_sva_501[158:155]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_9, and_dcpl_1359);
      FpAdd_8U_23U_qr_6_lpi_1_dfm_3_0 <= MUX_v_4_2_2((AluIn_data_sva_501[154:151]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_9, and_dcpl_1359);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_7_lpi_1_dfm_7_4 <= 4'b0;
      FpAdd_8U_23U_qr_7_lpi_1_dfm_3_0 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_154_cse ) begin
      FpAdd_8U_23U_qr_7_lpi_1_dfm_7_4 <= MUX_v_4_2_2((AluIn_data_sva_501[190:187]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_9, and_dcpl_1365);
      FpAdd_8U_23U_qr_7_lpi_1_dfm_3_0 <= MUX_v_4_2_2((AluIn_data_sva_501[186:183]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_9, and_dcpl_1365);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_8_lpi_1_dfm_7_4 <= 4'b0;
      FpAdd_8U_23U_qr_8_lpi_1_dfm_3_0 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_156_cse ) begin
      FpAdd_8U_23U_qr_8_lpi_1_dfm_7_4 <= MUX_v_4_2_2((AluIn_data_sva_501[222:219]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_9, and_dcpl_1371);
      FpAdd_8U_23U_qr_8_lpi_1_dfm_3_0 <= MUX_v_4_2_2((AluIn_data_sva_501[218:215]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_9, and_dcpl_1371);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_9_lpi_1_dfm_7_4 <= 4'b0;
      FpAdd_8U_23U_qr_9_lpi_1_dfm_3_0 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_158_cse ) begin
      FpAdd_8U_23U_qr_9_lpi_1_dfm_7_4 <= MUX_v_4_2_2((AluIn_data_sva_501[254:251]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_9, and_dcpl_1377);
      FpAdd_8U_23U_qr_9_lpi_1_dfm_3_0 <= MUX_v_4_2_2((AluIn_data_sva_501[250:247]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_9, and_dcpl_1377);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_10_lpi_1_dfm_7_4 <= 4'b0;
      FpAdd_8U_23U_qr_10_lpi_1_dfm_3_0 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_160_cse ) begin
      FpAdd_8U_23U_qr_10_lpi_1_dfm_7_4 <= MUX_v_4_2_2((AluIn_data_sva_501[286:283]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_9, and_dcpl_1383);
      FpAdd_8U_23U_qr_10_lpi_1_dfm_3_0 <= MUX_v_4_2_2((AluIn_data_sva_501[282:279]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_9, and_dcpl_1383);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_11_lpi_1_dfm_7_4 <= 4'b0;
      FpAdd_8U_23U_qr_11_lpi_1_dfm_3_0 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_162_cse ) begin
      FpAdd_8U_23U_qr_11_lpi_1_dfm_7_4 <= MUX_v_4_2_2((AluIn_data_sva_501[318:315]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_9, and_dcpl_1389);
      FpAdd_8U_23U_qr_11_lpi_1_dfm_3_0 <= MUX_v_4_2_2((AluIn_data_sva_501[314:311]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_9, and_dcpl_1389);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_12_lpi_1_dfm_7_4 <= 4'b0;
      FpAdd_8U_23U_qr_12_lpi_1_dfm_3_0 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_164_cse ) begin
      FpAdd_8U_23U_qr_12_lpi_1_dfm_7_4 <= MUX_v_4_2_2((AluIn_data_sva_501[350:347]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_9, and_dcpl_1395);
      FpAdd_8U_23U_qr_12_lpi_1_dfm_3_0 <= MUX_v_4_2_2((AluIn_data_sva_501[346:343]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_9, and_dcpl_1395);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_13_lpi_1_dfm_7_4 <= 4'b0;
      FpAdd_8U_23U_qr_13_lpi_1_dfm_3_0 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_166_cse ) begin
      FpAdd_8U_23U_qr_13_lpi_1_dfm_7_4 <= MUX_v_4_2_2((AluIn_data_sva_501[382:379]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_9, and_dcpl_1401);
      FpAdd_8U_23U_qr_13_lpi_1_dfm_3_0 <= MUX_v_4_2_2((AluIn_data_sva_501[378:375]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_9, and_dcpl_1401);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_14_lpi_1_dfm_7_4 <= 4'b0;
      FpAdd_8U_23U_qr_14_lpi_1_dfm_3_0 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_168_cse ) begin
      FpAdd_8U_23U_qr_14_lpi_1_dfm_7_4 <= MUX_v_4_2_2((AluIn_data_sva_501[414:411]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_9, and_dcpl_1407);
      FpAdd_8U_23U_qr_14_lpi_1_dfm_3_0 <= MUX_v_4_2_2((AluIn_data_sva_501[410:407]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_9, and_dcpl_1407);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_15_lpi_1_dfm_7_4 <= 4'b0;
      FpAdd_8U_23U_qr_15_lpi_1_dfm_3_0 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_170_cse ) begin
      FpAdd_8U_23U_qr_15_lpi_1_dfm_7_4 <= MUX_v_4_2_2((AluIn_data_sva_501[446:443]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_9, and_dcpl_1413);
      FpAdd_8U_23U_qr_15_lpi_1_dfm_3_0 <= MUX_v_4_2_2((AluIn_data_sva_501[442:439]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_9, and_dcpl_1413);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_16_lpi_1_dfm_7_4 <= 4'b0;
      FpAdd_8U_23U_qr_16_lpi_1_dfm_3_0 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_172_cse ) begin
      FpAdd_8U_23U_qr_16_lpi_1_dfm_7_4 <= MUX_v_4_2_2((AluIn_data_sva_501[478:475]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_9, and_dcpl_1419);
      FpAdd_8U_23U_qr_16_lpi_1_dfm_3_0 <= MUX_v_4_2_2((AluIn_data_sva_501[474:471]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_9, and_dcpl_1419);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_lpi_1_dfm_7_4 <= 4'b0;
      FpAdd_8U_23U_qr_lpi_1_dfm_3_0 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_and_174_cse ) begin
      FpAdd_8U_23U_qr_lpi_1_dfm_7_4 <= MUX_v_4_2_2((AluIn_data_sva_501[510:507]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_9, and_dcpl_1425);
      FpAdd_8U_23U_qr_lpi_1_dfm_3_0 <= MUX_v_4_2_2((AluIn_data_sva_501[506:503]),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_9, and_dcpl_1425);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_or_798_itm <= 1'b0;
      FpAlu_8U_23U_or_862_itm <= 1'b0;
      FpAlu_8U_23U_or_795_itm <= 1'b0;
      FpAlu_8U_23U_or_860_itm <= 1'b0;
      FpAlu_8U_23U_or_792_itm <= 1'b0;
      FpAlu_8U_23U_or_858_itm <= 1'b0;
      FpAlu_8U_23U_or_789_itm <= 1'b0;
      FpAlu_8U_23U_or_856_itm <= 1'b0;
      FpAlu_8U_23U_or_786_itm <= 1'b0;
      FpAlu_8U_23U_or_854_itm <= 1'b0;
      FpAlu_8U_23U_or_783_itm <= 1'b0;
      FpAlu_8U_23U_or_852_itm <= 1'b0;
      FpAlu_8U_23U_or_780_itm <= 1'b0;
      FpAlu_8U_23U_or_850_itm <= 1'b0;
      FpAlu_8U_23U_or_777_itm <= 1'b0;
      FpAlu_8U_23U_or_848_itm <= 1'b0;
      FpAlu_8U_23U_or_774_itm <= 1'b0;
      FpAlu_8U_23U_or_846_itm <= 1'b0;
      FpAlu_8U_23U_or_771_itm <= 1'b0;
      FpAlu_8U_23U_or_844_itm <= 1'b0;
      FpAlu_8U_23U_or_768_itm <= 1'b0;
      FpAlu_8U_23U_or_842_itm <= 1'b0;
      FpAlu_8U_23U_or_765_itm <= 1'b0;
      FpAlu_8U_23U_or_840_itm <= 1'b0;
      FpAlu_8U_23U_or_762_itm <= 1'b0;
      FpAlu_8U_23U_or_838_itm <= 1'b0;
      FpAlu_8U_23U_or_759_itm <= 1'b0;
      FpAlu_8U_23U_or_836_itm <= 1'b0;
      FpAlu_8U_23U_or_756_itm <= 1'b0;
      FpAlu_8U_23U_or_834_itm <= 1'b0;
      FpAlu_8U_23U_or_753_itm <= 1'b0;
      FpAlu_8U_23U_or_832_itm <= 1'b0;
    end
    else if ( FpAlu_8U_23U_and_1120_cse ) begin
      FpAlu_8U_23U_or_798_itm <= FpAlu_8U_23U_or_797_itm_mx0w0;
      FpAlu_8U_23U_or_862_itm <= FpAlu_8U_23U_or_861_itm_mx0w0;
      FpAlu_8U_23U_or_795_itm <= FpAlu_8U_23U_or_794_itm_mx0w0;
      FpAlu_8U_23U_or_860_itm <= FpAlu_8U_23U_or_859_itm_mx0w0;
      FpAlu_8U_23U_or_792_itm <= FpAlu_8U_23U_or_791_itm_mx0w0;
      FpAlu_8U_23U_or_858_itm <= FpAlu_8U_23U_or_857_itm_mx0w0;
      FpAlu_8U_23U_or_789_itm <= FpAlu_8U_23U_or_788_itm_mx0w0;
      FpAlu_8U_23U_or_856_itm <= FpAlu_8U_23U_or_855_itm_mx0w0;
      FpAlu_8U_23U_or_786_itm <= FpAlu_8U_23U_or_785_itm_mx0w0;
      FpAlu_8U_23U_or_854_itm <= FpAlu_8U_23U_or_853_itm_mx0w0;
      FpAlu_8U_23U_or_783_itm <= FpAlu_8U_23U_or_782_itm_mx0w0;
      FpAlu_8U_23U_or_852_itm <= FpAlu_8U_23U_or_851_itm_mx0w0;
      FpAlu_8U_23U_or_780_itm <= FpAlu_8U_23U_or_779_itm_mx0w0;
      FpAlu_8U_23U_or_850_itm <= FpAlu_8U_23U_or_849_itm_mx0w0;
      FpAlu_8U_23U_or_777_itm <= FpAlu_8U_23U_or_776_itm_mx0w0;
      FpAlu_8U_23U_or_848_itm <= FpAlu_8U_23U_or_847_itm_mx0w0;
      FpAlu_8U_23U_or_774_itm <= FpAlu_8U_23U_or_773_itm_mx0w0;
      FpAlu_8U_23U_or_846_itm <= FpAlu_8U_23U_or_845_itm_mx0w0;
      FpAlu_8U_23U_or_771_itm <= FpAlu_8U_23U_or_770_itm_mx0w0;
      FpAlu_8U_23U_or_844_itm <= FpAlu_8U_23U_or_843_itm_mx0w0;
      FpAlu_8U_23U_or_768_itm <= FpAlu_8U_23U_or_767_itm_mx0w0;
      FpAlu_8U_23U_or_842_itm <= FpAlu_8U_23U_or_841_itm_mx0w0;
      FpAlu_8U_23U_or_765_itm <= FpAlu_8U_23U_or_764_itm_mx0w0;
      FpAlu_8U_23U_or_840_itm <= FpAlu_8U_23U_or_839_itm_mx0w0;
      FpAlu_8U_23U_or_762_itm <= FpAlu_8U_23U_or_761_itm_mx0w0;
      FpAlu_8U_23U_or_838_itm <= FpAlu_8U_23U_or_837_itm_mx0w0;
      FpAlu_8U_23U_or_759_itm <= FpAlu_8U_23U_or_758_itm_mx0w0;
      FpAlu_8U_23U_or_836_itm <= FpAlu_8U_23U_or_835_itm_mx0w0;
      FpAlu_8U_23U_or_756_itm <= FpAlu_8U_23U_or_755_itm_mx0w0;
      FpAlu_8U_23U_or_834_itm <= FpAlu_8U_23U_or_833_itm_mx0w0;
      FpAlu_8U_23U_or_753_itm <= FpAlu_8U_23U_or_752_itm_mx0w0;
      FpAlu_8U_23U_or_832_itm <= FpAlu_8U_23U_or_831_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_and_60_itm <= 1'b0;
      FpAlu_8U_23U_nor_dfs <= 1'b0;
      FpAlu_8U_23U_equal_tmp_1 <= 1'b0;
      FpAlu_8U_23U_equal_tmp_2 <= 1'b0;
      FpAlu_8U_23U_equal_tmp <= 1'b0;
      FpAlu_8U_23U_and_56_itm <= 1'b0;
      FpAlu_8U_23U_and_52_itm <= 1'b0;
      FpAlu_8U_23U_and_48_itm <= 1'b0;
      FpAlu_8U_23U_and_44_itm <= 1'b0;
      FpAlu_8U_23U_and_40_itm <= 1'b0;
      FpAlu_8U_23U_and_36_itm <= 1'b0;
      FpAlu_8U_23U_and_32_itm <= 1'b0;
      FpAlu_8U_23U_and_28_itm <= 1'b0;
      FpAlu_8U_23U_and_24_itm <= 1'b0;
      FpAlu_8U_23U_and_20_itm <= 1'b0;
      FpAlu_8U_23U_and_16_itm <= 1'b0;
      FpAlu_8U_23U_and_12_itm <= 1'b0;
      FpAlu_8U_23U_and_8_itm <= 1'b0;
      FpAlu_8U_23U_and_4_itm <= 1'b0;
      FpAlu_8U_23U_and_itm <= 1'b0;
    end
    else if ( FpAlu_8U_23U_and_692_cse ) begin
      FpAlu_8U_23U_and_60_itm <= FpAlu_8U_23U_and_60_itm_mx0w0;
      FpAlu_8U_23U_nor_dfs <= FpAlu_8U_23U_nor_dfs_mx0w0;
      FpAlu_8U_23U_equal_tmp_1 <= and_3689_cse;
      FpAlu_8U_23U_equal_tmp_2 <= FpAlu_8U_23U_equal_tmp_2_mx0w0;
      FpAlu_8U_23U_equal_tmp <= FpAlu_8U_23U_equal_tmp_mx0w0;
      FpAlu_8U_23U_and_56_itm <= FpAlu_8U_23U_and_56_itm_mx0w0;
      FpAlu_8U_23U_and_52_itm <= FpAlu_8U_23U_and_52_itm_mx0w0;
      FpAlu_8U_23U_and_48_itm <= FpAlu_8U_23U_and_48_itm_mx0w0;
      FpAlu_8U_23U_and_44_itm <= FpAlu_8U_23U_and_44_itm_mx0w0;
      FpAlu_8U_23U_and_40_itm <= FpAlu_8U_23U_and_40_itm_mx0w0;
      FpAlu_8U_23U_and_36_itm <= FpAlu_8U_23U_and_36_itm_mx0w0;
      FpAlu_8U_23U_and_32_itm <= FpAlu_8U_23U_and_32_itm_mx0w0;
      FpAlu_8U_23U_and_28_itm <= FpAlu_8U_23U_and_28_itm_mx0w0;
      FpAlu_8U_23U_and_24_itm <= FpAlu_8U_23U_and_24_itm_mx0w0;
      FpAlu_8U_23U_and_20_itm <= FpAlu_8U_23U_and_20_itm_mx0w0;
      FpAlu_8U_23U_and_16_itm <= FpAlu_8U_23U_and_16_itm_mx0w0;
      FpAlu_8U_23U_and_12_itm <= FpAlu_8U_23U_and_12_itm_mx0w0;
      FpAlu_8U_23U_and_8_itm <= FpAlu_8U_23U_and_8_itm_mx0w0;
      FpAlu_8U_23U_and_4_itm <= FpAlu_8U_23U_and_4_itm_mx0w0;
      FpAlu_8U_23U_and_itm <= FpAlu_8U_23U_and_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_29 & and_dcpl_1426 & (~ IsNaN_8U_23U_2_land_lpi_1_dfm_st_1))
        | and_1895_rgt) & (~ mux_1425_itm) ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_1_land_lpi_1_dfm, and_1895_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_15_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_29 & and_dcpl_1426 & (~ IsNaN_8U_23U_2_land_15_lpi_1_dfm_st_1))
        | and_1899_rgt) & (~ mux_1425_itm) ) begin
      IsNaN_8U_23U_1_land_15_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_15_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_1_land_15_lpi_1_dfm, and_1899_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_14_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_29 & and_dcpl_1426 & (~ IsNaN_8U_23U_2_land_14_lpi_1_dfm_st_1))
        | and_1903_rgt) & (~ mux_1425_itm) ) begin
      IsNaN_8U_23U_1_land_14_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_14_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_1_land_14_lpi_1_dfm, and_1903_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_13_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_29 & and_dcpl_1426 & (~ IsNaN_8U_23U_2_land_13_lpi_1_dfm_st_1))
        | and_1907_rgt) & (~ mux_1425_itm) ) begin
      IsNaN_8U_23U_1_land_13_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_13_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_1_land_13_lpi_1_dfm, and_1907_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_11_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_29 & and_dcpl_1426 & (~ IsNaN_8U_23U_2_land_11_lpi_1_dfm_st_1))
        | and_1911_rgt) & (~ mux_1425_itm) ) begin
      IsNaN_8U_23U_1_land_11_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_11_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_1_land_11_lpi_1_dfm, and_1911_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_8_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & and_89_tmp & (~ mux_1425_itm) ) begin
      IsNaN_8U_23U_1_land_8_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_8_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_1_land_8_lpi_1_dfm, and_1917_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_7_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_29 & and_dcpl_1426 & (~ IsNaN_8U_23U_2_land_7_lpi_1_dfm_st_1))
        | and_1921_rgt) & (~ mux_1425_itm) ) begin
      IsNaN_8U_23U_1_land_7_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_7_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_1_land_7_lpi_1_dfm, and_1921_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_5_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_29 & and_dcpl_1426 & (~ IsNaN_8U_23U_2_land_5_lpi_1_dfm_st_1))
        | and_1925_rgt) & (~ mux_1425_itm) ) begin
      IsNaN_8U_23U_1_land_5_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_5_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_1_land_5_lpi_1_dfm, and_1925_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_29 & and_dcpl_1426 & (~ IsNaN_8U_23U_2_land_3_lpi_1_dfm_st_1))
        | and_1929_rgt) & (~ mux_1425_itm) ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_3_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_1_land_3_lpi_1_dfm, and_1929_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_29 & (~ (cfg_alu_algo_1_sva_st_92[0])) & (~ IsNaN_8U_23U_2_land_1_lpi_1_dfm_st_1)
        & (cfg_alu_algo_1_sva_st_92[1])) | and_1933_rgt) & (~ mux_1425_itm) ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_1_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_1_land_1_lpi_1_dfm, and_1933_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_if_mux_2_itm <= 1'b0;
      alu_loop_op_else_if_mux_1_itm <= 30'b0;
      alu_loop_op_else_if_mux_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_if_and_9_cse ) begin
      alu_loop_op_else_if_mux_2_itm <= MUX_s_1_2_2((AluIn_data_sva_501[0]), IntShiftLeft_16U_6U_32U_return_0_1_sva_2,
          and_dcpl_1476);
      alu_loop_op_else_if_mux_1_itm <= MUX_v_30_2_2((AluIn_data_sva_501[30:1]), IntShiftLeft_16U_6U_32U_return_30_1_1_sva_2,
          and_dcpl_1476);
      alu_loop_op_else_if_mux_itm <= MUX_s_1_2_2((AluIn_data_sva_501[31]), IntShiftLeft_16U_6U_32U_return_31_1_sva_2,
          and_dcpl_1476);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_2_itm <= 1'b0;
      alu_loop_op_else_else_if_mux_1_itm <= 30'b0;
      alu_loop_op_else_else_if_mux_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_9_cse ) begin
      alu_loop_op_else_else_if_mux_2_itm <= MUX_s_1_2_2((AluIn_data_sva_501[0]),
          IntShiftLeft_16U_6U_32U_return_0_1_sva_2, and_dcpl_1483);
      alu_loop_op_else_else_if_mux_1_itm <= MUX_v_30_2_2((AluIn_data_sva_501[30:1]),
          IntShiftLeft_16U_6U_32U_return_30_1_1_sva_2, and_dcpl_1483);
      alu_loop_op_else_else_if_mux_itm <= MUX_s_1_2_2((AluIn_data_sva_501[31]), IntShiftLeft_16U_6U_32U_return_31_1_sva_2,
          and_dcpl_1483);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_if_mux_5_itm <= 1'b0;
      alu_loop_op_else_if_mux_4_itm <= 30'b0;
      alu_loop_op_else_if_mux_3_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_if_and_12_cse ) begin
      alu_loop_op_else_if_mux_5_itm <= MUX_s_1_2_2((AluIn_data_sva_501[32]), IntShiftLeft_16U_6U_32U_return_0_2_sva_2,
          and_dcpl_1490);
      alu_loop_op_else_if_mux_4_itm <= MUX_v_30_2_2((AluIn_data_sva_501[62:33]),
          IntShiftLeft_16U_6U_32U_return_30_1_2_sva_2, and_dcpl_1490);
      alu_loop_op_else_if_mux_3_itm <= MUX_s_1_2_2((AluIn_data_sva_501[63]), IntShiftLeft_16U_6U_32U_return_31_2_sva_2,
          and_dcpl_1490);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_5_itm <= 1'b0;
      alu_loop_op_else_else_if_mux_4_itm <= 30'b0;
      alu_loop_op_else_else_if_mux_3_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_12_cse ) begin
      alu_loop_op_else_else_if_mux_5_itm <= MUX_s_1_2_2((AluIn_data_sva_501[32]),
          IntShiftLeft_16U_6U_32U_return_0_2_sva_2, and_dcpl_1497);
      alu_loop_op_else_else_if_mux_4_itm <= MUX_v_30_2_2((AluIn_data_sva_501[62:33]),
          IntShiftLeft_16U_6U_32U_return_30_1_2_sva_2, and_dcpl_1497);
      alu_loop_op_else_else_if_mux_3_itm <= MUX_s_1_2_2((AluIn_data_sva_501[63]),
          IntShiftLeft_16U_6U_32U_return_31_2_sva_2, and_dcpl_1497);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_if_mux_8_itm <= 1'b0;
      alu_loop_op_else_if_mux_7_itm <= 30'b0;
      alu_loop_op_else_if_mux_6_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_if_and_15_cse ) begin
      alu_loop_op_else_if_mux_8_itm <= MUX_s_1_2_2((AluIn_data_sva_501[64]), IntShiftLeft_16U_6U_32U_return_0_3_sva_2,
          and_dcpl_1504);
      alu_loop_op_else_if_mux_7_itm <= MUX_v_30_2_2((AluIn_data_sva_501[94:65]),
          IntShiftLeft_16U_6U_32U_return_30_1_3_sva_2, and_dcpl_1504);
      alu_loop_op_else_if_mux_6_itm <= MUX_s_1_2_2((AluIn_data_sva_501[95]), IntShiftLeft_16U_6U_32U_return_31_3_sva_2,
          and_dcpl_1504);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_8_itm <= 1'b0;
      alu_loop_op_else_else_if_mux_7_itm <= 30'b0;
      alu_loop_op_else_else_if_mux_6_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_15_cse ) begin
      alu_loop_op_else_else_if_mux_8_itm <= MUX_s_1_2_2((AluIn_data_sva_501[64]),
          IntShiftLeft_16U_6U_32U_return_0_3_sva_2, and_dcpl_1511);
      alu_loop_op_else_else_if_mux_7_itm <= MUX_v_30_2_2((AluIn_data_sva_501[94:65]),
          IntShiftLeft_16U_6U_32U_return_30_1_3_sva_2, and_dcpl_1511);
      alu_loop_op_else_else_if_mux_6_itm <= MUX_s_1_2_2((AluIn_data_sva_501[95]),
          IntShiftLeft_16U_6U_32U_return_31_3_sva_2, and_dcpl_1511);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_if_mux_11_itm <= 1'b0;
      alu_loop_op_else_if_mux_10_itm <= 30'b0;
      alu_loop_op_else_if_mux_9_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_if_and_18_cse ) begin
      alu_loop_op_else_if_mux_11_itm <= MUX_s_1_2_2((AluIn_data_sva_501[96]), IntShiftLeft_16U_6U_32U_return_0_4_sva_2,
          and_dcpl_1518);
      alu_loop_op_else_if_mux_10_itm <= MUX_v_30_2_2((AluIn_data_sva_501[126:97]),
          IntShiftLeft_16U_6U_32U_return_30_1_4_sva_2, and_dcpl_1518);
      alu_loop_op_else_if_mux_9_itm <= MUX_s_1_2_2((AluIn_data_sva_501[127]), IntShiftLeft_16U_6U_32U_return_31_4_sva_2,
          and_dcpl_1518);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_11_itm <= 1'b0;
      alu_loop_op_else_else_if_mux_10_itm <= 30'b0;
      alu_loop_op_else_else_if_mux_9_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_18_cse ) begin
      alu_loop_op_else_else_if_mux_11_itm <= MUX_s_1_2_2((AluIn_data_sva_501[96]),
          IntShiftLeft_16U_6U_32U_return_0_4_sva_2, and_dcpl_1525);
      alu_loop_op_else_else_if_mux_10_itm <= MUX_v_30_2_2((AluIn_data_sva_501[126:97]),
          IntShiftLeft_16U_6U_32U_return_30_1_4_sva_2, and_dcpl_1525);
      alu_loop_op_else_else_if_mux_9_itm <= MUX_s_1_2_2((AluIn_data_sva_501[127]),
          IntShiftLeft_16U_6U_32U_return_31_4_sva_2, and_dcpl_1525);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_if_mux_14_itm <= 1'b0;
      alu_loop_op_else_if_mux_13_itm <= 30'b0;
      alu_loop_op_else_if_mux_12_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_if_and_21_cse ) begin
      alu_loop_op_else_if_mux_14_itm <= MUX_s_1_2_2((AluIn_data_sva_501[128]), IntShiftLeft_16U_6U_32U_return_0_5_sva_2,
          and_dcpl_1532);
      alu_loop_op_else_if_mux_13_itm <= MUX_v_30_2_2((AluIn_data_sva_501[158:129]),
          IntShiftLeft_16U_6U_32U_return_30_1_5_sva_2, and_dcpl_1532);
      alu_loop_op_else_if_mux_12_itm <= MUX_s_1_2_2((AluIn_data_sva_501[159]), IntShiftLeft_16U_6U_32U_return_31_5_sva_2,
          and_dcpl_1532);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_14_itm <= 1'b0;
      alu_loop_op_else_else_if_mux_13_itm <= 30'b0;
      alu_loop_op_else_else_if_mux_12_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_21_cse ) begin
      alu_loop_op_else_else_if_mux_14_itm <= MUX_s_1_2_2((AluIn_data_sva_501[128]),
          IntShiftLeft_16U_6U_32U_return_0_5_sva_2, and_dcpl_1539);
      alu_loop_op_else_else_if_mux_13_itm <= MUX_v_30_2_2((AluIn_data_sva_501[158:129]),
          IntShiftLeft_16U_6U_32U_return_30_1_5_sva_2, and_dcpl_1539);
      alu_loop_op_else_else_if_mux_12_itm <= MUX_s_1_2_2((AluIn_data_sva_501[159]),
          IntShiftLeft_16U_6U_32U_return_31_5_sva_2, and_dcpl_1539);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_if_mux_17_itm <= 1'b0;
      alu_loop_op_else_if_mux_16_itm <= 30'b0;
      alu_loop_op_else_if_mux_15_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_if_and_24_cse ) begin
      alu_loop_op_else_if_mux_17_itm <= MUX_s_1_2_2((AluIn_data_sva_501[160]), IntShiftLeft_16U_6U_32U_return_0_6_sva_2,
          and_dcpl_1546);
      alu_loop_op_else_if_mux_16_itm <= MUX_v_30_2_2((AluIn_data_sva_501[190:161]),
          IntShiftLeft_16U_6U_32U_return_30_1_6_sva_2, and_dcpl_1546);
      alu_loop_op_else_if_mux_15_itm <= MUX_s_1_2_2((AluIn_data_sva_501[191]), IntShiftLeft_16U_6U_32U_return_31_6_sva_2,
          and_dcpl_1546);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_17_itm <= 1'b0;
      alu_loop_op_else_else_if_mux_16_itm <= 30'b0;
      alu_loop_op_else_else_if_mux_15_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_24_cse ) begin
      alu_loop_op_else_else_if_mux_17_itm <= MUX_s_1_2_2((AluIn_data_sva_501[160]),
          IntShiftLeft_16U_6U_32U_return_0_6_sva_2, and_dcpl_1553);
      alu_loop_op_else_else_if_mux_16_itm <= MUX_v_30_2_2((AluIn_data_sva_501[190:161]),
          IntShiftLeft_16U_6U_32U_return_30_1_6_sva_2, and_dcpl_1553);
      alu_loop_op_else_else_if_mux_15_itm <= MUX_s_1_2_2((AluIn_data_sva_501[191]),
          IntShiftLeft_16U_6U_32U_return_31_6_sva_2, and_dcpl_1553);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_if_mux_20_itm <= 1'b0;
      alu_loop_op_else_if_mux_19_itm <= 30'b0;
      alu_loop_op_else_if_mux_18_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_if_and_27_cse ) begin
      alu_loop_op_else_if_mux_20_itm <= MUX_s_1_2_2((AluIn_data_sva_501[192]), IntShiftLeft_16U_6U_32U_return_0_7_sva_2,
          and_dcpl_1560);
      alu_loop_op_else_if_mux_19_itm <= MUX_v_30_2_2((AluIn_data_sva_501[222:193]),
          IntShiftLeft_16U_6U_32U_return_30_1_7_sva_2, and_dcpl_1560);
      alu_loop_op_else_if_mux_18_itm <= MUX_s_1_2_2((AluIn_data_sva_501[223]), IntShiftLeft_16U_6U_32U_return_31_7_sva_2,
          and_dcpl_1560);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_20_itm <= 1'b0;
      alu_loop_op_else_else_if_mux_19_itm <= 30'b0;
      alu_loop_op_else_else_if_mux_18_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_27_cse ) begin
      alu_loop_op_else_else_if_mux_20_itm <= MUX_s_1_2_2((AluIn_data_sva_501[192]),
          IntShiftLeft_16U_6U_32U_return_0_7_sva_2, and_dcpl_1567);
      alu_loop_op_else_else_if_mux_19_itm <= MUX_v_30_2_2((AluIn_data_sva_501[222:193]),
          IntShiftLeft_16U_6U_32U_return_30_1_7_sva_2, and_dcpl_1567);
      alu_loop_op_else_else_if_mux_18_itm <= MUX_s_1_2_2((AluIn_data_sva_501[223]),
          IntShiftLeft_16U_6U_32U_return_31_7_sva_2, and_dcpl_1567);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_if_mux_23_itm <= 1'b0;
      alu_loop_op_else_if_mux_22_itm <= 30'b0;
      alu_loop_op_else_if_mux_21_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_if_and_30_cse ) begin
      alu_loop_op_else_if_mux_23_itm <= MUX_s_1_2_2((AluIn_data_sva_501[224]), IntShiftLeft_16U_6U_32U_return_0_8_sva_2,
          and_dcpl_1574);
      alu_loop_op_else_if_mux_22_itm <= MUX_v_30_2_2((AluIn_data_sva_501[254:225]),
          IntShiftLeft_16U_6U_32U_return_30_1_8_sva_2, and_dcpl_1574);
      alu_loop_op_else_if_mux_21_itm <= MUX_s_1_2_2((AluIn_data_sva_501[255]), IntShiftLeft_16U_6U_32U_return_31_8_sva_2,
          and_dcpl_1574);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_23_itm <= 1'b0;
      alu_loop_op_else_else_if_mux_22_itm <= 30'b0;
      alu_loop_op_else_else_if_mux_21_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_30_cse ) begin
      alu_loop_op_else_else_if_mux_23_itm <= MUX_s_1_2_2((AluIn_data_sva_501[224]),
          IntShiftLeft_16U_6U_32U_return_0_8_sva_2, and_dcpl_1581);
      alu_loop_op_else_else_if_mux_22_itm <= MUX_v_30_2_2((AluIn_data_sva_501[254:225]),
          IntShiftLeft_16U_6U_32U_return_30_1_8_sva_2, and_dcpl_1581);
      alu_loop_op_else_else_if_mux_21_itm <= MUX_s_1_2_2((AluIn_data_sva_501[255]),
          IntShiftLeft_16U_6U_32U_return_31_8_sva_2, and_dcpl_1581);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_if_mux_26_itm <= 1'b0;
      alu_loop_op_else_if_mux_25_itm <= 30'b0;
      alu_loop_op_else_if_mux_24_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_if_and_33_cse ) begin
      alu_loop_op_else_if_mux_26_itm <= MUX_s_1_2_2((AluIn_data_sva_501[256]), IntShiftLeft_16U_6U_32U_return_0_9_sva_2,
          and_dcpl_1588);
      alu_loop_op_else_if_mux_25_itm <= MUX_v_30_2_2((AluIn_data_sva_501[286:257]),
          IntShiftLeft_16U_6U_32U_return_30_1_9_sva_2, and_dcpl_1588);
      alu_loop_op_else_if_mux_24_itm <= MUX_s_1_2_2((AluIn_data_sva_501[287]), IntShiftLeft_16U_6U_32U_return_31_9_sva_2,
          and_dcpl_1588);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_26_itm <= 1'b0;
      alu_loop_op_else_else_if_mux_25_itm <= 30'b0;
      alu_loop_op_else_else_if_mux_24_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_33_cse ) begin
      alu_loop_op_else_else_if_mux_26_itm <= MUX_s_1_2_2((AluIn_data_sva_501[256]),
          IntShiftLeft_16U_6U_32U_return_0_9_sva_2, and_dcpl_1595);
      alu_loop_op_else_else_if_mux_25_itm <= MUX_v_30_2_2((AluIn_data_sva_501[286:257]),
          IntShiftLeft_16U_6U_32U_return_30_1_9_sva_2, and_dcpl_1595);
      alu_loop_op_else_else_if_mux_24_itm <= MUX_s_1_2_2((AluIn_data_sva_501[287]),
          IntShiftLeft_16U_6U_32U_return_31_9_sva_2, and_dcpl_1595);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_if_mux_29_itm <= 1'b0;
      alu_loop_op_else_if_mux_28_itm <= 30'b0;
      alu_loop_op_else_if_mux_27_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_if_and_36_cse ) begin
      alu_loop_op_else_if_mux_29_itm <= MUX_s_1_2_2((AluIn_data_sva_501[288]), IntShiftLeft_16U_6U_32U_return_0_10_sva_2,
          and_dcpl_1602);
      alu_loop_op_else_if_mux_28_itm <= MUX_v_30_2_2((AluIn_data_sva_501[318:289]),
          IntShiftLeft_16U_6U_32U_return_30_1_10_sva_2, and_dcpl_1602);
      alu_loop_op_else_if_mux_27_itm <= MUX_s_1_2_2((AluIn_data_sva_501[319]), IntShiftLeft_16U_6U_32U_return_31_10_sva_2,
          and_dcpl_1602);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_29_itm <= 1'b0;
      alu_loop_op_else_else_if_mux_28_itm <= 30'b0;
      alu_loop_op_else_else_if_mux_27_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_36_cse ) begin
      alu_loop_op_else_else_if_mux_29_itm <= MUX_s_1_2_2((AluIn_data_sva_501[288]),
          IntShiftLeft_16U_6U_32U_return_0_10_sva_2, and_dcpl_1609);
      alu_loop_op_else_else_if_mux_28_itm <= MUX_v_30_2_2((AluIn_data_sva_501[318:289]),
          IntShiftLeft_16U_6U_32U_return_30_1_10_sva_2, and_dcpl_1609);
      alu_loop_op_else_else_if_mux_27_itm <= MUX_s_1_2_2((AluIn_data_sva_501[319]),
          IntShiftLeft_16U_6U_32U_return_31_10_sva_2, and_dcpl_1609);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_if_mux_32_itm <= 1'b0;
      alu_loop_op_else_if_mux_31_itm <= 30'b0;
      alu_loop_op_else_if_mux_30_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_if_and_39_cse ) begin
      alu_loop_op_else_if_mux_32_itm <= MUX_s_1_2_2((AluIn_data_sva_501[320]), IntShiftLeft_16U_6U_32U_return_0_11_sva_2,
          and_dcpl_1616);
      alu_loop_op_else_if_mux_31_itm <= MUX_v_30_2_2((AluIn_data_sva_501[350:321]),
          IntShiftLeft_16U_6U_32U_return_30_1_11_sva_2, and_dcpl_1616);
      alu_loop_op_else_if_mux_30_itm <= MUX_s_1_2_2((AluIn_data_sva_501[351]), IntShiftLeft_16U_6U_32U_return_31_11_sva_2,
          and_dcpl_1616);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_32_itm <= 1'b0;
      alu_loop_op_else_else_if_mux_31_itm <= 30'b0;
      alu_loop_op_else_else_if_mux_30_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_39_cse ) begin
      alu_loop_op_else_else_if_mux_32_itm <= MUX_s_1_2_2((AluIn_data_sva_501[320]),
          IntShiftLeft_16U_6U_32U_return_0_11_sva_2, and_dcpl_1623);
      alu_loop_op_else_else_if_mux_31_itm <= MUX_v_30_2_2((AluIn_data_sva_501[350:321]),
          IntShiftLeft_16U_6U_32U_return_30_1_11_sva_2, and_dcpl_1623);
      alu_loop_op_else_else_if_mux_30_itm <= MUX_s_1_2_2((AluIn_data_sva_501[351]),
          IntShiftLeft_16U_6U_32U_return_31_11_sva_2, and_dcpl_1623);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_if_mux_35_itm <= 1'b0;
      alu_loop_op_else_if_mux_34_itm <= 30'b0;
      alu_loop_op_else_if_mux_33_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_if_and_42_cse ) begin
      alu_loop_op_else_if_mux_35_itm <= MUX_s_1_2_2((AluIn_data_sva_501[352]), IntShiftLeft_16U_6U_32U_return_0_12_sva_2,
          and_dcpl_1630);
      alu_loop_op_else_if_mux_34_itm <= MUX_v_30_2_2((AluIn_data_sva_501[382:353]),
          IntShiftLeft_16U_6U_32U_return_30_1_12_sva_2, and_dcpl_1630);
      alu_loop_op_else_if_mux_33_itm <= MUX_s_1_2_2((AluIn_data_sva_501[383]), IntShiftLeft_16U_6U_32U_return_31_12_sva_2,
          and_dcpl_1630);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_35_itm <= 1'b0;
      alu_loop_op_else_else_if_mux_34_itm <= 30'b0;
      alu_loop_op_else_else_if_mux_33_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_42_cse ) begin
      alu_loop_op_else_else_if_mux_35_itm <= MUX_s_1_2_2((AluIn_data_sva_501[352]),
          IntShiftLeft_16U_6U_32U_return_0_12_sva_2, and_dcpl_1637);
      alu_loop_op_else_else_if_mux_34_itm <= MUX_v_30_2_2((AluIn_data_sva_501[382:353]),
          IntShiftLeft_16U_6U_32U_return_30_1_12_sva_2, and_dcpl_1637);
      alu_loop_op_else_else_if_mux_33_itm <= MUX_s_1_2_2((AluIn_data_sva_501[383]),
          IntShiftLeft_16U_6U_32U_return_31_12_sva_2, and_dcpl_1637);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_if_mux_38_itm <= 1'b0;
      alu_loop_op_else_if_mux_37_itm <= 30'b0;
      alu_loop_op_else_if_mux_36_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_if_and_45_cse ) begin
      alu_loop_op_else_if_mux_38_itm <= MUX_s_1_2_2((AluIn_data_sva_501[384]), IntShiftLeft_16U_6U_32U_return_0_13_sva_2,
          and_dcpl_1644);
      alu_loop_op_else_if_mux_37_itm <= MUX_v_30_2_2((AluIn_data_sva_501[414:385]),
          IntShiftLeft_16U_6U_32U_return_30_1_13_sva_2, and_dcpl_1644);
      alu_loop_op_else_if_mux_36_itm <= MUX_s_1_2_2((AluIn_data_sva_501[415]), IntShiftLeft_16U_6U_32U_return_31_13_sva_2,
          and_dcpl_1644);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_38_itm <= 1'b0;
      alu_loop_op_else_else_if_mux_37_itm <= 30'b0;
      alu_loop_op_else_else_if_mux_36_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_45_cse ) begin
      alu_loop_op_else_else_if_mux_38_itm <= MUX_s_1_2_2((AluIn_data_sva_501[384]),
          IntShiftLeft_16U_6U_32U_return_0_13_sva_2, and_dcpl_1651);
      alu_loop_op_else_else_if_mux_37_itm <= MUX_v_30_2_2((AluIn_data_sva_501[414:385]),
          IntShiftLeft_16U_6U_32U_return_30_1_13_sva_2, and_dcpl_1651);
      alu_loop_op_else_else_if_mux_36_itm <= MUX_s_1_2_2((AluIn_data_sva_501[415]),
          IntShiftLeft_16U_6U_32U_return_31_13_sva_2, and_dcpl_1651);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_if_mux_41_itm <= 1'b0;
      alu_loop_op_else_if_mux_40_itm <= 30'b0;
      alu_loop_op_else_if_mux_39_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_if_and_48_cse ) begin
      alu_loop_op_else_if_mux_41_itm <= MUX_s_1_2_2((AluIn_data_sva_501[416]), IntShiftLeft_16U_6U_32U_return_0_14_sva_2,
          and_dcpl_1658);
      alu_loop_op_else_if_mux_40_itm <= MUX_v_30_2_2((AluIn_data_sva_501[446:417]),
          IntShiftLeft_16U_6U_32U_return_30_1_14_sva_2, and_dcpl_1658);
      alu_loop_op_else_if_mux_39_itm <= MUX_s_1_2_2((AluIn_data_sva_501[447]), IntShiftLeft_16U_6U_32U_return_31_14_sva_2,
          and_dcpl_1658);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_41_itm <= 1'b0;
      alu_loop_op_else_else_if_mux_40_itm <= 30'b0;
      alu_loop_op_else_else_if_mux_39_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_48_cse ) begin
      alu_loop_op_else_else_if_mux_41_itm <= MUX_s_1_2_2((AluIn_data_sva_501[416]),
          IntShiftLeft_16U_6U_32U_return_0_14_sva_2, and_dcpl_1665);
      alu_loop_op_else_else_if_mux_40_itm <= MUX_v_30_2_2((AluIn_data_sva_501[446:417]),
          IntShiftLeft_16U_6U_32U_return_30_1_14_sva_2, and_dcpl_1665);
      alu_loop_op_else_else_if_mux_39_itm <= MUX_s_1_2_2((AluIn_data_sva_501[447]),
          IntShiftLeft_16U_6U_32U_return_31_14_sva_2, and_dcpl_1665);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_if_mux_44_itm <= 1'b0;
      alu_loop_op_else_if_mux_43_itm <= 30'b0;
      alu_loop_op_else_if_mux_42_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_if_and_51_cse ) begin
      alu_loop_op_else_if_mux_44_itm <= MUX_s_1_2_2((AluIn_data_sva_501[448]), IntShiftLeft_16U_6U_32U_return_0_15_sva_2,
          and_dcpl_1672);
      alu_loop_op_else_if_mux_43_itm <= MUX_v_30_2_2((AluIn_data_sva_501[478:449]),
          IntShiftLeft_16U_6U_32U_return_30_1_15_sva_2, and_dcpl_1672);
      alu_loop_op_else_if_mux_42_itm <= MUX_s_1_2_2((AluIn_data_sva_501[479]), IntShiftLeft_16U_6U_32U_return_31_15_sva_2,
          and_dcpl_1672);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_44_itm <= 1'b0;
      alu_loop_op_else_else_if_mux_43_itm <= 30'b0;
      alu_loop_op_else_else_if_mux_42_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_51_cse ) begin
      alu_loop_op_else_else_if_mux_44_itm <= MUX_s_1_2_2((AluIn_data_sva_501[448]),
          IntShiftLeft_16U_6U_32U_return_0_15_sva_2, and_dcpl_1679);
      alu_loop_op_else_else_if_mux_43_itm <= MUX_v_30_2_2((AluIn_data_sva_501[478:449]),
          IntShiftLeft_16U_6U_32U_return_30_1_15_sva_2, and_dcpl_1679);
      alu_loop_op_else_else_if_mux_42_itm <= MUX_s_1_2_2((AluIn_data_sva_501[479]),
          IntShiftLeft_16U_6U_32U_return_31_15_sva_2, and_dcpl_1679);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_if_mux_47_itm <= 1'b0;
      alu_loop_op_else_if_mux_46_itm <= 30'b0;
      alu_loop_op_else_if_mux_45_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_if_and_54_cse ) begin
      alu_loop_op_else_if_mux_47_itm <= MUX_s_1_2_2((AluIn_data_sva_501[480]), IntShiftLeft_16U_6U_32U_return_0_sva_2,
          and_dcpl_1686);
      alu_loop_op_else_if_mux_46_itm <= MUX_v_30_2_2((AluIn_data_sva_501[510:481]),
          IntShiftLeft_16U_6U_32U_return_30_1_sva_2, and_dcpl_1686);
      alu_loop_op_else_if_mux_45_itm <= MUX_s_1_2_2((AluIn_data_sva_501[511]), IntShiftLeft_16U_6U_32U_return_31_sva_2,
          and_dcpl_1686);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_else_else_if_mux_47_itm <= 1'b0;
      alu_loop_op_else_else_if_mux_46_itm <= 30'b0;
      alu_loop_op_else_else_if_mux_45_itm <= 1'b0;
    end
    else if ( alu_loop_op_else_else_if_and_54_cse ) begin
      alu_loop_op_else_else_if_mux_47_itm <= MUX_s_1_2_2((AluIn_data_sva_501[480]),
          IntShiftLeft_16U_6U_32U_return_0_sva_2, and_dcpl_1691);
      alu_loop_op_else_else_if_mux_46_itm <= MUX_v_30_2_2((AluIn_data_sva_501[510:481]),
          IntShiftLeft_16U_6U_32U_return_30_1_sva_2, and_dcpl_1691);
      alu_loop_op_else_else_if_mux_45_itm <= MUX_s_1_2_2((AluIn_data_sva_501[511]),
          IntShiftLeft_16U_6U_32U_return_31_sva_2, and_dcpl_1691);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_12_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_28 & (~ (cfg_precision[0])) & (~ (cfg_alu_algo_1_sva_st_92[0]))
        & and_dcpl_1692 & (~ IsNaN_8U_23U_2_land_12_lpi_1_dfm_st_1)) | and_2163_rgt)
        & (~ mux_1425_itm) ) begin
      IsNaN_8U_23U_1_land_12_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_12_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_1_land_12_lpi_1_dfm, and_2163_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_10_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_29 & (~ (cfg_alu_algo_1_sva_st_92[0])) & (~ IsNaN_8U_23U_2_land_10_lpi_1_dfm_st_1)
        & (cfg_alu_algo_1_sva_st_92[1])) | and_2167_rgt) & (~ mux_1425_itm) ) begin
      IsNaN_8U_23U_1_land_10_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_10_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_1_land_10_lpi_1_dfm, and_2167_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_9_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_29 & and_dcpl_1426 & (~ IsNaN_8U_23U_2_land_9_lpi_1_dfm_st_1))
        | and_2171_rgt) & (~ mux_1425_itm) ) begin
      IsNaN_8U_23U_1_land_9_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_9_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_1_land_9_lpi_1_dfm, and_2171_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_6_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_29 & and_dcpl_1426 & (~ IsNaN_8U_23U_2_land_6_lpi_1_dfm_st_1))
        | and_2175_rgt) & (~ mux_1425_itm) ) begin
      IsNaN_8U_23U_1_land_6_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_6_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_1_land_6_lpi_1_dfm, and_2175_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_4_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_29 & and_dcpl_1426 & (~ IsNaN_8U_23U_2_land_4_lpi_1_dfm_st_1))
        | and_2179_rgt) & (~ mux_1425_itm) ) begin
      IsNaN_8U_23U_1_land_4_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_4_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_1_land_4_lpi_1_dfm, and_2179_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_29 & and_dcpl_1426 & (~ IsNaN_8U_23U_2_land_2_lpi_1_dfm_st_1))
        | and_2183_rgt) & (~ mux_1425_itm) ) begin
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_2_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_1_land_2_lpi_1_dfm, and_2183_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_nan_to_zero_op_sign_1_lpi_1_dfm_4 <= 1'b0;
      alu_nan_to_zero_op_sign_2_lpi_1_dfm_4 <= 1'b0;
      alu_nan_to_zero_op_sign_3_lpi_1_dfm_4 <= 1'b0;
      alu_nan_to_zero_op_sign_4_lpi_1_dfm_4 <= 1'b0;
      alu_nan_to_zero_op_sign_5_lpi_1_dfm_4 <= 1'b0;
      alu_nan_to_zero_op_sign_6_lpi_1_dfm_4 <= 1'b0;
      alu_nan_to_zero_op_sign_7_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( alu_nan_to_zero_op_sign_and_25_cse ) begin
      alu_nan_to_zero_op_sign_1_lpi_1_dfm_4 <= MUX_s_1_2_2(alu_nan_to_zero_op_sign_1_lpi_1_dfm_mx0w0,
          alu_nan_to_zero_op_sign_1_lpi_1_dfm, and_dcpl_23);
      alu_nan_to_zero_op_sign_2_lpi_1_dfm_4 <= MUX_s_1_2_2(alu_nan_to_zero_op_sign_2_lpi_1_dfm_mx0w0,
          alu_nan_to_zero_op_sign_2_lpi_1_dfm, and_dcpl_23);
      alu_nan_to_zero_op_sign_3_lpi_1_dfm_4 <= MUX_s_1_2_2(alu_nan_to_zero_op_sign_3_lpi_1_dfm_mx0w0,
          alu_nan_to_zero_op_sign_3_lpi_1_dfm, and_dcpl_23);
      alu_nan_to_zero_op_sign_4_lpi_1_dfm_4 <= MUX_s_1_2_2(alu_nan_to_zero_op_sign_4_lpi_1_dfm_mx0w0,
          alu_nan_to_zero_op_sign_4_lpi_1_dfm, and_dcpl_23);
      alu_nan_to_zero_op_sign_5_lpi_1_dfm_4 <= MUX_s_1_2_2(alu_nan_to_zero_op_sign_5_lpi_1_dfm_mx0w0,
          alu_nan_to_zero_op_sign_5_lpi_1_dfm, and_dcpl_23);
      alu_nan_to_zero_op_sign_6_lpi_1_dfm_4 <= MUX_s_1_2_2(alu_nan_to_zero_op_sign_6_lpi_1_dfm_mx0w0,
          alu_nan_to_zero_op_sign_6_lpi_1_dfm, and_dcpl_23);
      alu_nan_to_zero_op_sign_7_lpi_1_dfm_4 <= MUX_s_1_2_2(alu_nan_to_zero_op_sign_7_lpi_1_dfm_mx0w0,
          alu_nan_to_zero_op_sign_7_lpi_1_dfm, and_dcpl_23);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_FpCmp_8U_23U_true_else_slc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | io_read_cfg_alu_bypass_rsc_svs_st_5 | (reg_cfg_alu_algo_1_sva_st_93_cse[0])
        | or_dcpl_787)) ) begin
      alu_loop_op_1_FpCmp_8U_23U_true_else_slc_8_svs <= FpCmp_8U_23U_false_else_if_acc_16_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_FpCmp_8U_23U_false_else_slc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~
        (reg_cfg_alu_algo_1_sva_st_93_cse[0])) | or_dcpl_787)) ) begin
      alu_loop_op_1_FpCmp_8U_23U_false_else_slc_8_svs <= FpCmp_8U_23U_false_else_if_acc_16_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_2 <= 1'b0;
      alu_loop_op_10_FpCmp_8U_23U_false_slc_8_1_svs_2 <= 1'b0;
    end
    else if ( FpCmp_8U_23U_false_if_and_48_cse ) begin
      alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_16_itm_8_1,
          alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_st, alu_loop_op_1_FpCmp_8U_23U_true_slc_8_svs_st,
          alu_loop_op_1_FpAdd_8U_23U_is_a_greater_slc_8_svs, {and_dcpl_22 , and_dcpl_34
          , and_dcpl_36 , and_2185_rgt});
      alu_loop_op_10_FpCmp_8U_23U_false_slc_8_1_svs_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_34_itm_8_1,
          alu_loop_op_10_FpCmp_8U_23U_false_slc_8_1_svs_st, alu_loop_op_10_FpCmp_8U_23U_true_slc_8_1_svs_st,
          alu_loop_op_10_FpAdd_8U_23U_is_a_greater_slc_8_1_svs, {and_dcpl_22 , and_dcpl_34
          , and_dcpl_36 , and_2185_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_2_FpCmp_8U_23U_true_else_slc_8_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | or_tmp_39 | (reg_cfg_alu_algo_1_sva_st_93_cse!=2'b00)))
        ) begin
      alu_loop_op_2_FpCmp_8U_23U_true_else_slc_8_1_svs <= FpCmp_8U_23U_false_else_if_acc_18_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_2_FpCmp_8U_23U_false_else_slc_8_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | or_tmp_39 | (reg_cfg_alu_algo_1_sva_st_93_cse!=2'b01)))
        ) begin
      alu_loop_op_2_FpCmp_8U_23U_false_else_slc_8_1_svs <= FpCmp_8U_23U_false_else_if_acc_18_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_2 <= 1'b0;
      alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_2 <= 1'b0;
      alu_loop_op_4_FpCmp_8U_23U_false_slc_8_1_svs_2 <= 1'b0;
      alu_loop_op_5_FpCmp_8U_23U_false_slc_8_svs_2 <= 1'b0;
      alu_loop_op_6_FpCmp_8U_23U_false_slc_8_1_svs_2 <= 1'b0;
      alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_2 <= 1'b0;
      alu_loop_op_9_FpCmp_8U_23U_false_slc_8_svs_2 <= 1'b0;
      alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_2 <= 1'b0;
      alu_loop_op_13_FpCmp_8U_23U_false_slc_8_svs_2 <= 1'b0;
      alu_loop_op_14_FpCmp_8U_23U_false_slc_8_1_svs_2 <= 1'b0;
      alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_2 <= 1'b0;
      alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_2 <= 1'b0;
    end
    else if ( FpCmp_8U_23U_false_if_and_49_cse ) begin
      alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_18_itm_8_1,
          alu_loop_op_2_FpCmp_8U_23U_false_slc_8_1_svs_st, alu_loop_op_2_FpCmp_8U_23U_true_slc_8_1_svs_st,
          reg_alu_loop_op_2_FpAdd_8U_23U_is_a_greater_slc_8_1_svs_cse, {and_dcpl_22
          , and_dcpl_34 , and_dcpl_36 , and_2186_rgt});
      alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_20_itm_8_1,
          alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_st, alu_loop_op_3_FpCmp_8U_23U_true_slc_8_svs_st,
          alu_loop_op_3_FpAdd_8U_23U_is_a_greater_slc_8_svs, {and_dcpl_22 , and_dcpl_34
          , and_dcpl_36 , and_2186_rgt});
      alu_loop_op_4_FpCmp_8U_23U_false_slc_8_1_svs_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_22_itm_8_1,
          alu_loop_op_4_FpCmp_8U_23U_false_slc_8_1_svs_st, alu_loop_op_4_FpCmp_8U_23U_true_slc_8_1_svs_st,
          alu_loop_op_4_FpAdd_8U_23U_is_a_greater_slc_8_1_svs, {and_dcpl_22 , and_dcpl_34
          , and_dcpl_36 , and_2186_rgt});
      alu_loop_op_5_FpCmp_8U_23U_false_slc_8_svs_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_24_itm_8_1,
          alu_loop_op_5_FpCmp_8U_23U_false_slc_8_svs_st, alu_loop_op_5_FpCmp_8U_23U_true_slc_8_svs_st,
          alu_loop_op_5_FpAdd_8U_23U_is_a_greater_slc_8_svs, {and_dcpl_22 , and_dcpl_34
          , and_dcpl_36 , and_2186_rgt});
      alu_loop_op_6_FpCmp_8U_23U_false_slc_8_1_svs_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_26_itm_8_1,
          alu_loop_op_6_FpCmp_8U_23U_false_slc_8_1_svs_st, alu_loop_op_6_FpCmp_8U_23U_true_slc_8_1_svs_st,
          alu_loop_op_6_FpAdd_8U_23U_is_a_greater_slc_8_1_svs, {and_dcpl_22 , and_dcpl_34
          , and_dcpl_36 , and_2186_rgt});
      alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_28_itm_8_1,
          alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_st, alu_loop_op_7_FpCmp_8U_23U_true_slc_8_svs_st,
          alu_loop_op_7_FpAdd_8U_23U_is_a_greater_slc_8_svs, {and_dcpl_22 , and_dcpl_34
          , and_dcpl_36 , and_2186_rgt});
      alu_loop_op_9_FpCmp_8U_23U_false_slc_8_svs_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_32_itm_8_1,
          alu_loop_op_9_FpCmp_8U_23U_false_slc_8_svs_st, alu_loop_op_9_FpCmp_8U_23U_true_slc_8_svs_st,
          alu_loop_op_9_FpAdd_8U_23U_is_a_greater_slc_8_svs, {and_dcpl_22 , and_dcpl_34
          , and_dcpl_36 , and_2186_rgt});
      alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_36_itm_8_1,
          alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_st, alu_loop_op_11_FpCmp_8U_23U_true_slc_8_svs_st,
          alu_loop_op_11_FpAdd_8U_23U_is_a_greater_slc_8_svs, {and_dcpl_22 , and_dcpl_34
          , and_dcpl_36 , and_2186_rgt});
      alu_loop_op_13_FpCmp_8U_23U_false_slc_8_svs_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_40_itm_8_1,
          alu_loop_op_13_FpCmp_8U_23U_false_slc_8_svs_st, alu_loop_op_13_FpCmp_8U_23U_true_slc_8_svs_st,
          alu_loop_op_13_FpAdd_8U_23U_is_a_greater_slc_8_svs, {and_dcpl_22 , and_dcpl_34
          , and_dcpl_36 , and_2186_rgt});
      alu_loop_op_14_FpCmp_8U_23U_false_slc_8_1_svs_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_42_itm_8_1,
          alu_loop_op_14_FpCmp_8U_23U_false_slc_8_1_svs_st, alu_loop_op_14_FpCmp_8U_23U_true_slc_8_1_svs_st,
          alu_loop_op_14_FpAdd_8U_23U_is_a_greater_slc_8_1_svs, {and_dcpl_22 , and_dcpl_34
          , and_dcpl_36 , and_2186_rgt});
      alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_44_itm_8_1,
          alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_st, alu_loop_op_15_FpCmp_8U_23U_true_slc_8_svs_st,
          alu_loop_op_15_FpAdd_8U_23U_is_a_greater_slc_8_svs, {and_dcpl_22 , and_dcpl_34
          , and_dcpl_36 , and_2186_rgt});
      alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_46_itm_8_1,
          alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_st, alu_loop_op_16_FpCmp_8U_23U_true_slc_8_1_svs_st,
          alu_loop_op_16_FpAdd_8U_23U_is_a_greater_slc_8_1_svs, {and_dcpl_22 , and_dcpl_34
          , and_dcpl_36 , and_2186_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_3_FpCmp_8U_23U_true_else_slc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | or_tmp_55 | (reg_cfg_alu_algo_1_sva_st_93_cse!=2'b00)))
        ) begin
      alu_loop_op_3_FpCmp_8U_23U_true_else_slc_8_svs <= FpCmp_8U_23U_false_else_if_acc_20_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_3_FpCmp_8U_23U_false_else_slc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | or_tmp_55 | (reg_cfg_alu_algo_1_sva_st_93_cse!=2'b01)))
        ) begin
      alu_loop_op_3_FpCmp_8U_23U_false_else_slc_8_svs <= FpCmp_8U_23U_false_else_if_acc_20_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_4_FpCmp_8U_23U_true_else_slc_8_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | or_tmp_76 | (reg_cfg_alu_algo_1_sva_st_93_cse!=2'b00)))
        ) begin
      alu_loop_op_4_FpCmp_8U_23U_true_else_slc_8_1_svs <= FpCmp_8U_23U_false_else_if_acc_22_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_4_FpCmp_8U_23U_false_else_slc_8_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | or_tmp_76 | (reg_cfg_alu_algo_1_sva_st_93_cse!=2'b01)))
        ) begin
      alu_loop_op_4_FpCmp_8U_23U_false_else_slc_8_1_svs <= FpCmp_8U_23U_false_else_if_acc_22_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_5_FpCmp_8U_23U_true_else_slc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | or_tmp_97 | (reg_cfg_alu_algo_1_sva_st_93_cse!=2'b00)))
        ) begin
      alu_loop_op_5_FpCmp_8U_23U_true_else_slc_8_svs <= FpCmp_8U_23U_false_else_if_acc_24_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_5_FpCmp_8U_23U_false_else_slc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | or_tmp_97 | (reg_cfg_alu_algo_1_sva_st_93_cse!=2'b01)))
        ) begin
      alu_loop_op_5_FpCmp_8U_23U_false_else_slc_8_svs <= FpCmp_8U_23U_false_else_if_acc_24_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_6_FpCmp_8U_23U_true_else_slc_8_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | io_read_cfg_alu_bypass_rsc_svs_st_5 | (reg_cfg_alu_algo_1_sva_st_93_cse[0])
        | or_dcpl_823)) ) begin
      alu_loop_op_6_FpCmp_8U_23U_true_else_slc_8_1_svs <= FpCmp_8U_23U_false_else_if_acc_26_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_6_FpCmp_8U_23U_false_else_slc_8_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~
        (reg_cfg_alu_algo_1_sva_st_93_cse[0])) | or_dcpl_823)) ) begin
      alu_loop_op_6_FpCmp_8U_23U_false_else_slc_8_1_svs <= FpCmp_8U_23U_false_else_if_acc_26_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_7_FpCmp_8U_23U_true_else_slc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | io_read_cfg_alu_bypass_rsc_svs_st_5 | (reg_cfg_alu_algo_1_sva_st_93_cse[0])
        | or_dcpl_830)) ) begin
      alu_loop_op_7_FpCmp_8U_23U_true_else_slc_8_svs <= FpCmp_8U_23U_false_else_if_acc_28_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_7_FpCmp_8U_23U_false_else_slc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~
        (reg_cfg_alu_algo_1_sva_st_93_cse[0])) | or_dcpl_830)) ) begin
      alu_loop_op_7_FpCmp_8U_23U_false_else_slc_8_svs <= FpCmp_8U_23U_false_else_if_acc_28_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_nan_to_zero_op_sign_8_lpi_1_dfm_3 <= 1'b0;
      alu_nan_to_zero_op_sign_9_lpi_1_dfm_3 <= 1'b0;
      alu_nan_to_zero_op_sign_10_lpi_1_dfm_3 <= 1'b0;
      alu_nan_to_zero_op_sign_11_lpi_1_dfm_3 <= 1'b0;
      alu_nan_to_zero_op_sign_12_lpi_1_dfm_3 <= 1'b0;
      alu_nan_to_zero_op_sign_13_lpi_1_dfm_3 <= 1'b0;
      alu_nan_to_zero_op_sign_14_lpi_1_dfm_3 <= 1'b0;
      alu_nan_to_zero_op_sign_15_lpi_1_dfm_3 <= 1'b0;
      alu_nan_to_zero_op_sign_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( alu_nan_to_zero_op_sign_and_cse ) begin
      alu_nan_to_zero_op_sign_8_lpi_1_dfm_3 <= MUX_s_1_2_2(alu_nan_to_zero_op_sign_8_lpi_1_dfm_mx0w0,
          alu_nan_to_zero_op_sign_8_lpi_1_dfm, and_dcpl_23);
      alu_nan_to_zero_op_sign_9_lpi_1_dfm_3 <= MUX_s_1_2_2(alu_nan_to_zero_op_sign_9_lpi_1_dfm_mx0w0,
          alu_nan_to_zero_op_sign_9_lpi_1_dfm, and_dcpl_23);
      alu_nan_to_zero_op_sign_10_lpi_1_dfm_3 <= MUX_s_1_2_2(alu_nan_to_zero_op_sign_10_lpi_1_dfm_mx0w0,
          alu_nan_to_zero_op_sign_10_lpi_1_dfm, and_dcpl_23);
      alu_nan_to_zero_op_sign_11_lpi_1_dfm_3 <= MUX_s_1_2_2(alu_nan_to_zero_op_sign_11_lpi_1_dfm_mx0w0,
          alu_nan_to_zero_op_sign_11_lpi_1_dfm, and_dcpl_23);
      alu_nan_to_zero_op_sign_12_lpi_1_dfm_3 <= MUX_s_1_2_2(alu_nan_to_zero_op_sign_12_lpi_1_dfm_mx0w0,
          alu_nan_to_zero_op_sign_12_lpi_1_dfm, and_dcpl_23);
      alu_nan_to_zero_op_sign_13_lpi_1_dfm_3 <= MUX_s_1_2_2(alu_nan_to_zero_op_sign_13_lpi_1_dfm_mx0w0,
          alu_nan_to_zero_op_sign_13_lpi_1_dfm, and_dcpl_23);
      alu_nan_to_zero_op_sign_14_lpi_1_dfm_3 <= MUX_s_1_2_2(alu_nan_to_zero_op_sign_14_lpi_1_dfm_mx0w0,
          alu_nan_to_zero_op_sign_14_lpi_1_dfm, and_dcpl_23);
      alu_nan_to_zero_op_sign_15_lpi_1_dfm_3 <= MUX_s_1_2_2(alu_nan_to_zero_op_sign_15_lpi_1_dfm_mx0w0,
          alu_nan_to_zero_op_sign_15_lpi_1_dfm, and_dcpl_23);
      alu_nan_to_zero_op_sign_lpi_1_dfm_3 <= MUX_s_1_2_2(alu_nan_to_zero_op_sign_lpi_1_dfm_mx0w0,
          alu_nan_to_zero_op_sign_lpi_1_dfm, and_dcpl_23);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_8_FpCmp_8U_23U_true_else_slc_8_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | io_read_cfg_alu_bypass_rsc_svs_st_5 | (reg_cfg_alu_algo_1_sva_st_93_cse[0])
        | or_dcpl_837)) ) begin
      alu_loop_op_8_FpCmp_8U_23U_true_else_slc_8_1_svs <= FpCmp_8U_23U_false_else_if_acc_30_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_8_FpCmp_8U_23U_false_else_slc_8_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~
        (reg_cfg_alu_algo_1_sva_st_93_cse[0])) | or_dcpl_837)) ) begin
      alu_loop_op_8_FpCmp_8U_23U_false_else_slc_8_1_svs <= FpCmp_8U_23U_false_else_if_acc_30_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_2 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_22 | and_dcpl_34 | and_dcpl_127 | and_2193_rgt)
        & (~ mux_16_itm) ) begin
      alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_30_itm_8_1,
          alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_st, alu_loop_op_8_FpCmp_8U_23U_true_slc_8_1_svs_st,
          alu_loop_op_8_FpAdd_8U_23U_is_a_greater_slc_8_1_svs, {and_dcpl_22 , and_dcpl_34
          , and_dcpl_127 , and_2193_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_9_FpCmp_8U_23U_true_else_slc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | io_read_cfg_alu_bypass_rsc_svs_st_5 | (reg_cfg_alu_algo_1_sva_st_93_cse[0])
        | or_dcpl_844)) ) begin
      alu_loop_op_9_FpCmp_8U_23U_true_else_slc_8_svs <= FpCmp_8U_23U_false_else_if_acc_32_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_9_FpCmp_8U_23U_false_else_slc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~
        (reg_cfg_alu_algo_1_sva_st_93_cse[0])) | or_dcpl_844)) ) begin
      alu_loop_op_9_FpCmp_8U_23U_false_else_slc_8_svs <= FpCmp_8U_23U_false_else_if_acc_32_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_10_FpCmp_8U_23U_true_else_slc_8_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | io_read_cfg_alu_bypass_rsc_svs_st_5 | (reg_cfg_alu_algo_1_sva_st_93_cse[0])
        | or_dcpl_851)) ) begin
      alu_loop_op_10_FpCmp_8U_23U_true_else_slc_8_1_svs <= FpCmp_8U_23U_false_else_if_acc_34_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_10_FpCmp_8U_23U_false_else_slc_8_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~
        (reg_cfg_alu_algo_1_sva_st_93_cse[0])) | or_dcpl_851)) ) begin
      alu_loop_op_10_FpCmp_8U_23U_false_else_slc_8_1_svs <= FpCmp_8U_23U_false_else_if_acc_34_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_11_FpCmp_8U_23U_true_else_slc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | or_dcpl_859 | (reg_cfg_alu_algo_1_sva_st_93_cse[0])
        | alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_st_2)) ) begin
      alu_loop_op_11_FpCmp_8U_23U_true_else_slc_8_svs <= FpCmp_8U_23U_false_else_if_acc_36_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_11_FpCmp_8U_23U_false_else_slc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | or_dcpl_859 | (~ (reg_cfg_alu_algo_1_sva_st_93_cse[0]))
        | alu_loop_op_11_FpCmp_8U_23U_false_slc_8_svs_st_2)) ) begin
      alu_loop_op_11_FpCmp_8U_23U_false_else_slc_8_svs <= FpCmp_8U_23U_false_else_if_acc_36_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_12_FpCmp_8U_23U_true_else_slc_8_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | or_dcpl_859 | alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_st_2
        | (reg_cfg_alu_algo_1_sva_st_93_cse[0]))) ) begin
      alu_loop_op_12_FpCmp_8U_23U_true_else_slc_8_1_svs <= FpCmp_8U_23U_false_else_if_acc_38_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_12_FpCmp_8U_23U_false_else_slc_8_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | or_dcpl_859 | alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_st_2
        | (~ (reg_cfg_alu_algo_1_sva_st_93_cse[0])))) ) begin
      alu_loop_op_12_FpCmp_8U_23U_false_else_slc_8_1_svs <= FpCmp_8U_23U_false_else_if_acc_38_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_2 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_22 | and_dcpl_34 | and_dcpl_127 | and_2198_rgt)
        & (~ mux_16_itm) ) begin
      alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_2 <= MUX1HOT_s_1_4_2(FpCmp_8U_23U_true_if_acc_38_itm_8_1,
          alu_loop_op_12_FpCmp_8U_23U_false_slc_8_1_svs_st, alu_loop_op_12_FpCmp_8U_23U_true_slc_8_1_svs_st,
          alu_loop_op_12_FpAdd_8U_23U_is_a_greater_slc_8_1_svs, {and_dcpl_22 , and_dcpl_34
          , and_dcpl_127 , and_2198_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_13_FpCmp_8U_23U_true_else_slc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | io_read_cfg_alu_bypass_rsc_svs_st_5 | (reg_cfg_alu_algo_1_sva_st_93_cse[0])
        | or_dcpl_872)) ) begin
      alu_loop_op_13_FpCmp_8U_23U_true_else_slc_8_svs <= FpCmp_8U_23U_false_else_if_acc_40_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_13_FpCmp_8U_23U_false_else_slc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~
        (reg_cfg_alu_algo_1_sva_st_93_cse[0])) | or_dcpl_872)) ) begin
      alu_loop_op_13_FpCmp_8U_23U_false_else_slc_8_svs <= FpCmp_8U_23U_false_else_if_acc_40_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_14_FpCmp_8U_23U_true_else_slc_8_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | io_read_cfg_alu_bypass_rsc_svs_st_5 | (reg_cfg_alu_algo_1_sva_st_93_cse[0])
        | or_dcpl_879)) ) begin
      alu_loop_op_14_FpCmp_8U_23U_true_else_slc_8_1_svs <= FpCmp_8U_23U_false_else_if_acc_42_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_14_FpCmp_8U_23U_false_else_slc_8_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~
        (reg_cfg_alu_algo_1_sva_st_93_cse[0])) | or_dcpl_879)) ) begin
      alu_loop_op_14_FpCmp_8U_23U_false_else_slc_8_1_svs <= FpCmp_8U_23U_false_else_if_acc_42_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_15_FpCmp_8U_23U_true_else_slc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | or_dcpl_859 | alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_st_2
        | (reg_cfg_alu_algo_1_sva_st_93_cse[0]))) ) begin
      alu_loop_op_15_FpCmp_8U_23U_true_else_slc_8_svs <= FpCmp_8U_23U_false_else_if_acc_44_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_15_FpCmp_8U_23U_false_else_slc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | or_dcpl_859 | alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_st_2
        | (~ (reg_cfg_alu_algo_1_sva_st_93_cse[0])))) ) begin
      alu_loop_op_15_FpCmp_8U_23U_false_else_slc_8_svs <= FpCmp_8U_23U_false_else_if_acc_44_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_16_FpCmp_8U_23U_true_else_slc_8_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | io_read_cfg_alu_bypass_rsc_svs_st_5 | (reg_cfg_alu_algo_1_sva_st_93_cse[0])
        | or_dcpl_893)) ) begin
      alu_loop_op_16_FpCmp_8U_23U_true_else_slc_8_1_svs <= FpCmp_8U_23U_false_else_if_acc_46_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_16_FpCmp_8U_23U_false_else_slc_8_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_790 | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~
        (reg_cfg_alu_algo_1_sva_st_93_cse[0])) | or_dcpl_893)) ) begin
      alu_loop_op_16_FpCmp_8U_23U_false_else_slc_8_1_svs <= FpCmp_8U_23U_false_else_if_acc_46_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftLeft_16U_6U_32U_return_0_1_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_1_sva_2 <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_1_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_2_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_2_sva_2 <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_2_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_3_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_3_sva_2 <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_3_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_4_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_4_sva_2 <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_4_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_5_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_5_sva_2 <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_5_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_6_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_6_sva_2 <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_6_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_7_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_7_sva_2 <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_7_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_8_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_8_sva_2 <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_8_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_9_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_9_sva_2 <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_9_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_10_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_10_sva_2 <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_10_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_11_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_11_sva_2 <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_11_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_12_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_12_sva_2 <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_12_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_13_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_13_sva_2 <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_13_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_14_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_14_sva_2 <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_14_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_15_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_15_sva_2 <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_15_sva_2 <= 1'b0;
    end
    else if ( IntShiftLeft_16U_6U_32U_and_48_cse ) begin
      IntShiftLeft_16U_6U_32U_return_0_1_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_0_1_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_0_1_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_30_1_1_sva_2 <= MUX_v_30_2_2(IntShiftLeft_16U_6U_32U_return_30_1_1_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_30_1_1_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_31_1_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_31_1_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_31_1_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_0_2_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_0_2_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_0_2_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_30_1_2_sva_2 <= MUX_v_30_2_2(IntShiftLeft_16U_6U_32U_return_30_1_2_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_30_1_2_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_31_2_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_31_2_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_31_2_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_0_3_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_0_3_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_0_3_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_30_1_3_sva_2 <= MUX_v_30_2_2(IntShiftLeft_16U_6U_32U_return_30_1_3_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_30_1_3_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_31_3_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_31_3_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_31_3_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_0_4_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_0_4_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_0_4_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_30_1_4_sva_2 <= MUX_v_30_2_2(IntShiftLeft_16U_6U_32U_return_30_1_4_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_30_1_4_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_31_4_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_31_4_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_31_4_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_0_5_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_0_5_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_0_5_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_30_1_5_sva_2 <= MUX_v_30_2_2(IntShiftLeft_16U_6U_32U_return_30_1_5_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_30_1_5_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_31_5_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_31_5_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_31_5_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_0_6_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_0_6_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_0_6_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_30_1_6_sva_2 <= MUX_v_30_2_2(IntShiftLeft_16U_6U_32U_return_30_1_6_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_30_1_6_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_31_6_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_31_6_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_31_6_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_0_7_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_0_7_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_0_7_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_30_1_7_sva_2 <= MUX_v_30_2_2(IntShiftLeft_16U_6U_32U_return_30_1_7_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_30_1_7_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_31_7_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_31_7_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_31_7_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_0_8_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_0_8_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_0_8_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_30_1_8_sva_2 <= MUX_v_30_2_2(IntShiftLeft_16U_6U_32U_return_30_1_8_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_30_1_8_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_31_8_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_31_8_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_31_8_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_0_9_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_0_9_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_0_9_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_30_1_9_sva_2 <= MUX_v_30_2_2(IntShiftLeft_16U_6U_32U_return_30_1_9_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_30_1_9_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_31_9_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_31_9_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_31_9_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_0_10_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_0_10_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_0_10_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_30_1_10_sva_2 <= MUX_v_30_2_2(IntShiftLeft_16U_6U_32U_return_30_1_10_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_30_1_10_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_31_10_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_31_10_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_31_10_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_0_11_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_0_11_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_0_11_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_30_1_11_sva_2 <= MUX_v_30_2_2(IntShiftLeft_16U_6U_32U_return_30_1_11_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_30_1_11_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_31_11_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_31_11_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_31_11_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_0_12_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_0_12_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_0_12_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_30_1_12_sva_2 <= MUX_v_30_2_2(IntShiftLeft_16U_6U_32U_return_30_1_12_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_30_1_12_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_31_12_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_31_12_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_31_12_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_0_13_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_0_13_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_0_13_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_30_1_13_sva_2 <= MUX_v_30_2_2(IntShiftLeft_16U_6U_32U_return_30_1_13_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_30_1_13_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_31_13_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_31_13_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_31_13_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_0_14_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_0_14_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_0_14_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_30_1_14_sva_2 <= MUX_v_30_2_2(IntShiftLeft_16U_6U_32U_return_30_1_14_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_30_1_14_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_31_14_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_31_14_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_31_14_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_0_15_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_0_15_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_0_15_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_30_1_15_sva_2 <= MUX_v_30_2_2(IntShiftLeft_16U_6U_32U_return_30_1_15_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_30_1_15_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_31_15_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_31_15_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_31_15_sva, and_dcpl_22);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftLeft_16U_6U_32U_return_0_sva_2 <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_sva_2 <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_sva_2 <= 1'b0;
    end
    else if ( IntShiftLeft_16U_6U_32U_and_93_cse ) begin
      IntShiftLeft_16U_6U_32U_return_0_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_0_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_0_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_30_1_sva_2 <= MUX_v_30_2_2(IntShiftLeft_16U_6U_32U_return_30_1_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_30_1_sva, and_dcpl_22);
      IntShiftLeft_16U_6U_32U_return_31_sva_2 <= MUX_s_1_2_2(IntShiftLeft_16U_6U_32U_return_31_sva_mx0w0,
          IntShiftLeft_16U_6U_32U_return_31_sva, and_dcpl_22);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= 1'b0;
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= 1'b0;
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= 1'b0;
      alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= 1'b0;
      alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= 1'b0;
      alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= 1'b0;
      alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= 1'b0;
      alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= 1'b0;
      alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= 1'b0;
      alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= 1'b0;
      alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= 1'b0;
      alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= 1'b0;
      alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= 1'b0;
      alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= 1'b0;
      alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= 1'b0;
    end
    else if ( IsZero_8U_23U_and_cse ) begin
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= MUX_s_1_2_2(alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0,
          alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm, or_tmp_3479);
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= MUX_s_1_2_2(alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0,
          alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm, or_tmp_3479);
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= MUX_s_1_2_2(alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0,
          alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm, or_tmp_3479);
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= MUX_s_1_2_2(alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0,
          alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm, or_tmp_3479);
      alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= MUX_s_1_2_2(alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0,
          alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_or_itm, or_tmp_3479);
      alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= MUX_s_1_2_2(alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0,
          alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_or_itm, or_tmp_3479);
      alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= MUX_s_1_2_2(alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0,
          alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_or_itm, or_tmp_3479);
      alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= MUX_s_1_2_2(alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0,
          alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_or_itm, or_tmp_3479);
      alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= MUX_s_1_2_2(alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0,
          alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_or_itm, or_tmp_3479);
      alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= MUX_s_1_2_2(alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0,
          alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_or_itm, or_tmp_3479);
      alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= MUX_s_1_2_2(alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0,
          alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_or_itm, or_tmp_3479);
      alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= MUX_s_1_2_2(alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0,
          alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_or_itm, or_tmp_3479);
      alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= MUX_s_1_2_2(alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0,
          alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_or_itm, or_tmp_3479);
      alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= MUX_s_1_2_2(alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0,
          alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_or_itm, or_tmp_3479);
      alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= MUX_s_1_2_2(alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0,
          alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_or_itm, or_tmp_3479);
      alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_or_itm_1 <= MUX_s_1_2_2(alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0,
          alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_or_itm, or_tmp_3479);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_algo_1_sva_st_31 <= 2'b0;
    end
    else if ( core_wen & (~(and_dcpl_21 | or_dcpl_3 | (fsm_output[0]))) ) begin
      cfg_alu_algo_1_sva_st_31 <= cfg_alu_algo_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_393 | or_dcpl_699)) ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm <= IsNaN_8U_23U_3_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_2_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_393 | or_dcpl_785)) ) begin
      IsNaN_8U_23U_1_land_2_lpi_1_dfm <= IsNaN_8U_23U_3_land_2_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_393 | or_dcpl_696)) ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm <= IsNaN_8U_23U_3_land_3_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_4_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_393 | or_dcpl_783)) ) begin
      IsNaN_8U_23U_1_land_4_lpi_1_dfm <= IsNaN_8U_23U_3_land_4_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_5_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_393 | or_dcpl_694)) ) begin
      IsNaN_8U_23U_1_land_5_lpi_1_dfm <= IsNaN_8U_23U_3_land_5_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_6_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_393 | or_dcpl_780)) ) begin
      IsNaN_8U_23U_1_land_6_lpi_1_dfm <= IsNaN_8U_23U_3_land_6_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_7_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_393 | or_dcpl_692)) ) begin
      IsNaN_8U_23U_1_land_7_lpi_1_dfm <= IsNaN_8U_23U_3_land_7_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_8_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_13 | (cfg_precision[0]) | (cfg_alu_algo_1_sva_st_92!=2'b10)
        | IsNaN_8U_23U_2_land_8_lpi_1_dfm_st_1 | (~ and_89_tmp))) ) begin
      IsNaN_8U_23U_1_land_8_lpi_1_dfm <= IsNaN_8U_23U_3_land_8_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_9_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_393 | or_dcpl_777)) ) begin
      IsNaN_8U_23U_1_land_9_lpi_1_dfm <= IsNaN_8U_23U_3_land_9_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_10_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_393 | or_dcpl_775)) ) begin
      IsNaN_8U_23U_1_land_10_lpi_1_dfm <= IsNaN_8U_23U_3_land_10_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_11_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_393 | or_dcpl_688)) ) begin
      IsNaN_8U_23U_1_land_11_lpi_1_dfm <= IsNaN_8U_23U_3_land_11_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_12_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_13 | (cfg_precision[0]) | (cfg_alu_algo_1_sva_st_92!=2'b10)
        | (~ and_89_tmp) | IsNaN_8U_23U_2_land_12_lpi_1_dfm_st_1)) ) begin
      IsNaN_8U_23U_1_land_12_lpi_1_dfm <= IsNaN_8U_23U_3_land_12_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_13_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_393 | or_dcpl_686)) ) begin
      IsNaN_8U_23U_1_land_13_lpi_1_dfm <= IsNaN_8U_23U_3_land_13_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_14_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_393 | or_dcpl_683)) ) begin
      IsNaN_8U_23U_1_land_14_lpi_1_dfm <= IsNaN_8U_23U_3_land_14_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_15_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_393 | or_dcpl_681)) ) begin
      IsNaN_8U_23U_1_land_15_lpi_1_dfm <= IsNaN_8U_23U_3_land_15_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_393 | or_dcpl_679)) ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm <= IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftLeft_16U_6U_32U_return_31_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_sva <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_15_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_15_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_15_sva <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_14_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_14_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_14_sva <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_13_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_13_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_13_sva <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_12_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_12_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_12_sva <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_11_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_11_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_11_sva <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_10_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_10_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_10_sva <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_9_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_9_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_9_sva <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_8_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_8_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_8_sva <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_7_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_7_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_7_sva <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_6_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_6_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_6_sva <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_5_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_5_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_5_sva <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_4_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_4_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_4_sva <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_3_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_3_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_3_sva <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_2_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_2_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_2_sva <= 30'b0;
      IntShiftLeft_16U_6U_32U_return_31_1_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_0_1_sva <= 1'b0;
      IntShiftLeft_16U_6U_32U_return_30_1_1_sva <= 30'b0;
    end
    else if ( IntShiftLeft_16U_6U_32U_and_cse ) begin
      IntShiftLeft_16U_6U_32U_return_31_sva <= IntShiftLeft_16U_6U_32U_return_31_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_0_sva <= IntShiftLeft_16U_6U_32U_return_0_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_30_1_sva <= IntShiftLeft_16U_6U_32U_return_30_1_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_31_15_sva <= IntShiftLeft_16U_6U_32U_return_31_15_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_0_15_sva <= IntShiftLeft_16U_6U_32U_return_0_15_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_30_1_15_sva <= IntShiftLeft_16U_6U_32U_return_30_1_15_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_31_14_sva <= IntShiftLeft_16U_6U_32U_return_31_14_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_0_14_sva <= IntShiftLeft_16U_6U_32U_return_0_14_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_30_1_14_sva <= IntShiftLeft_16U_6U_32U_return_30_1_14_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_31_13_sva <= IntShiftLeft_16U_6U_32U_return_31_13_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_0_13_sva <= IntShiftLeft_16U_6U_32U_return_0_13_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_30_1_13_sva <= IntShiftLeft_16U_6U_32U_return_30_1_13_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_31_12_sva <= IntShiftLeft_16U_6U_32U_return_31_12_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_0_12_sva <= IntShiftLeft_16U_6U_32U_return_0_12_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_30_1_12_sva <= IntShiftLeft_16U_6U_32U_return_30_1_12_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_31_11_sva <= IntShiftLeft_16U_6U_32U_return_31_11_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_0_11_sva <= IntShiftLeft_16U_6U_32U_return_0_11_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_30_1_11_sva <= IntShiftLeft_16U_6U_32U_return_30_1_11_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_31_10_sva <= IntShiftLeft_16U_6U_32U_return_31_10_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_0_10_sva <= IntShiftLeft_16U_6U_32U_return_0_10_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_30_1_10_sva <= IntShiftLeft_16U_6U_32U_return_30_1_10_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_31_9_sva <= IntShiftLeft_16U_6U_32U_return_31_9_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_0_9_sva <= IntShiftLeft_16U_6U_32U_return_0_9_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_30_1_9_sva <= IntShiftLeft_16U_6U_32U_return_30_1_9_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_31_8_sva <= IntShiftLeft_16U_6U_32U_return_31_8_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_0_8_sva <= IntShiftLeft_16U_6U_32U_return_0_8_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_30_1_8_sva <= IntShiftLeft_16U_6U_32U_return_30_1_8_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_31_7_sva <= IntShiftLeft_16U_6U_32U_return_31_7_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_0_7_sva <= IntShiftLeft_16U_6U_32U_return_0_7_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_30_1_7_sva <= IntShiftLeft_16U_6U_32U_return_30_1_7_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_31_6_sva <= IntShiftLeft_16U_6U_32U_return_31_6_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_0_6_sva <= IntShiftLeft_16U_6U_32U_return_0_6_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_30_1_6_sva <= IntShiftLeft_16U_6U_32U_return_30_1_6_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_31_5_sva <= IntShiftLeft_16U_6U_32U_return_31_5_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_0_5_sva <= IntShiftLeft_16U_6U_32U_return_0_5_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_30_1_5_sva <= IntShiftLeft_16U_6U_32U_return_30_1_5_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_31_4_sva <= IntShiftLeft_16U_6U_32U_return_31_4_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_0_4_sva <= IntShiftLeft_16U_6U_32U_return_0_4_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_30_1_4_sva <= IntShiftLeft_16U_6U_32U_return_30_1_4_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_31_3_sva <= IntShiftLeft_16U_6U_32U_return_31_3_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_0_3_sva <= IntShiftLeft_16U_6U_32U_return_0_3_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_30_1_3_sva <= IntShiftLeft_16U_6U_32U_return_30_1_3_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_31_2_sva <= IntShiftLeft_16U_6U_32U_return_31_2_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_0_2_sva <= IntShiftLeft_16U_6U_32U_return_0_2_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_30_1_2_sva <= IntShiftLeft_16U_6U_32U_return_30_1_2_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_31_1_sva <= IntShiftLeft_16U_6U_32U_return_31_1_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_0_1_sva <= IntShiftLeft_16U_6U_32U_return_0_1_sva_mx0w0;
      IntShiftLeft_16U_6U_32U_return_30_1_1_sva <= IntShiftLeft_16U_6U_32U_return_30_1_1_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_4_land_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_4_land_15_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_4_land_14_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_4_land_13_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_4_land_12_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_4_land_11_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_4_land_10_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_4_land_9_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_4_land_8_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_4_land_7_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_4_land_6_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_4_land_5_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_4_land_4_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_4_land_3_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_4_land_2_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_4_land_1_lpi_1_dfm_4 <= 1'b0;
      cfg_alu_algo_1_sva_1 <= 2'b0;
      cfg_alu_shift_value_1_sva_1 <= 6'b0;
    end
    else if ( cfg_alu_src_and_cse ) begin
      IsNaN_8U_23U_4_land_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_4_land_15_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_15_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_4_land_14_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_14_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_4_land_13_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_13_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_4_land_12_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_12_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_4_land_11_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_11_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_4_land_10_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_10_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_4_land_9_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_9_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_4_land_8_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_8_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_4_land_7_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_7_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_4_land_6_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_6_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_4_land_5_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_5_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_4_land_4_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_4_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_4_land_3_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_3_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_4_land_2_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_2_lpi_1_dfm_mx1w0;
      IsNaN_8U_23U_4_land_1_lpi_1_dfm_4 <= IsNaN_8U_23U_2_land_1_lpi_1_dfm_mx1w0;
      cfg_alu_algo_1_sva_1 <= cfg_alu_algo_rsci_d;
      cfg_alu_shift_value_1_sva_1 <= cfg_alu_shift_value_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= 1'b0;
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= 1'b0;
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= 1'b0;
      alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= 1'b0;
      alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= 1'b0;
      alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= 1'b0;
      alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= 1'b0;
      alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= 1'b0;
      alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= 1'b0;
      alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= 1'b0;
      alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= 1'b0;
      alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= 1'b0;
      alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= 1'b0;
      alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= 1'b0;
      alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= 1'b0;
    end
    else if ( IsZero_8U_23U_and_16_cse ) begin
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
      alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= alu_loop_op_5_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
      alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= alu_loop_op_6_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
      alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= alu_loop_op_7_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
      alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= alu_loop_op_8_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
      alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= alu_loop_op_9_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
      alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= alu_loop_op_10_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
      alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= alu_loop_op_11_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
      alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= alu_loop_op_12_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
      alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= alu_loop_op_13_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
      alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= alu_loop_op_14_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
      alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= alu_loop_op_15_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
      alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_or_itm <= alu_loop_op_16_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp_2 <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp_2 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_cse ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_6_tmp_2;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_6_tmp_2;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_6_tmp_2;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_6_tmp_2;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_6_tmp_2;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_6_tmp_2;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_6_tmp_2;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_6_tmp_2;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_6_tmp_2;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_6_tmp_2;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_6_tmp_2;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_6_tmp_2;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_6_tmp_2;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_6_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_tmp_2 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_95_ssc ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_tmp_2 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_94_ssc ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_tmp_2 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_93_ssc ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_tmp_2 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_92_ssc ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_tmp_2 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_91_ssc ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_tmp_2 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_90_ssc ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_tmp_2 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_89_ssc ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_tmp_2 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_88_ssc ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_tmp_2 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_87_ssc ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_tmp_2 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_86_ssc ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_tmp_2 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_85_ssc ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_tmp_2 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_84_ssc ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_tmp_2 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_83_ssc ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_tmp_2 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_82_ssc ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_tmp_2 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_81_ssc ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_tmp <= 10'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_tmp_1 <= 3'b0;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_tmp_2 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_80_ssc ) begin
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_tmp <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_tmp_1 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp_1;
      reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_tmp_2 <= reg_FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_tmp_2;
    end
  end
  assign FpAlu_8U_23U_mux1h_1039_nl = MUX1HOT_v_22_3_2((FpAdd_8U_23U_o_mant_1_lpi_1_dfm_2_mx0[22:1]),
      (FpCmp_8U_23U_true_o_22_0_1_lpi_1_dfm_6[22:1]), (FpCmp_8U_23U_false_o_22_0_1_lpi_1_dfm_6[22:1]),
      {FpAlu_8U_23U_nor_dfs_79 , FpAlu_8U_23U_equal_tmp_235 , FpAlu_8U_23U_equal_tmp_239});
  assign FpAlu_8U_23U_not_80_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_3_nl = MUX_v_22_2_2(22'b0000000000000000000000, (FpAlu_8U_23U_mux1h_1039_nl),
      (FpAlu_8U_23U_not_80_nl));
  assign FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_15_nl = MUX_v_4_2_2(FpAdd_8U_23U_o_expo_1_lpi_1_dfm_2_7_4,
      (FpAdd_8U_23U_o_expo_1_sva_4[7:4]), FpAdd_8U_23U_and_51_ssc);
  assign FpAlu_8U_23U_nor_16_nl = ~(MUX_v_4_2_2((FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_15_nl),
      4'b1111, FpAdd_8U_23U_and_113_ssc));
  assign FpAlu_8U_23U_FpAlu_8U_23U_nor_16_nl = ~(MUX_v_4_2_2((FpAlu_8U_23U_nor_16_nl),
      4'b1111, FpAlu_8U_23U_equal_tmp_237));
  assign and_4125_nl = nor_7_ssc & (~(or_dcpl_1047 | and_dcpl_1796));
  assign FpAlu_8U_23U_mux1h_1036_nl = MUX1HOT_v_22_3_2((FpAdd_8U_23U_o_mant_2_lpi_1_dfm_2_mx0[22:1]),
      (FpCmp_8U_23U_true_o_22_0_2_lpi_1_dfm_6[22:1]), (FpCmp_8U_23U_false_o_22_0_2_lpi_1_dfm_6[22:1]),
      {FpAlu_8U_23U_nor_dfs_79 , FpAlu_8U_23U_equal_tmp_235 , FpAlu_8U_23U_equal_tmp_239});
  assign FpAlu_8U_23U_not_82_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_7_nl = MUX_v_22_2_2(22'b0000000000000000000000, (FpAlu_8U_23U_mux1h_1036_nl),
      (FpAlu_8U_23U_not_82_nl));
  assign FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_14_nl = MUX_v_4_2_2(FpAdd_8U_23U_o_expo_2_lpi_1_dfm_2_7_4,
      (FpAdd_8U_23U_o_expo_2_sva_4[7:4]), FpAdd_8U_23U_and_55_ssc);
  assign FpAlu_8U_23U_nor_15_nl = ~(MUX_v_4_2_2((FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_14_nl),
      4'b1111, FpAdd_8U_23U_and_115_ssc));
  assign FpAlu_8U_23U_FpAlu_8U_23U_nor_15_nl = ~(MUX_v_4_2_2((FpAlu_8U_23U_nor_15_nl),
      4'b1111, FpAlu_8U_23U_equal_tmp_237));
  assign and_4119_nl = nor_7_ssc & (~(or_dcpl_1052 | and_dcpl_1804));
  assign FpAlu_8U_23U_mux1h_1033_nl = MUX1HOT_v_22_3_2((FpAdd_8U_23U_o_mant_3_lpi_1_dfm_2_mx0[22:1]),
      (FpCmp_8U_23U_true_o_22_0_3_lpi_1_dfm_6[22:1]), (FpCmp_8U_23U_false_o_22_0_3_lpi_1_dfm_6[22:1]),
      {FpAlu_8U_23U_nor_dfs_79 , FpAlu_8U_23U_equal_tmp_235 , FpAlu_8U_23U_equal_tmp_239});
  assign FpAlu_8U_23U_not_84_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_11_nl = MUX_v_22_2_2(22'b0000000000000000000000, (FpAlu_8U_23U_mux1h_1033_nl),
      (FpAlu_8U_23U_not_84_nl));
  assign FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_13_nl = MUX_v_4_2_2(FpAdd_8U_23U_o_expo_3_lpi_1_dfm_2_7_4,
      (FpAdd_8U_23U_o_expo_3_sva_4[7:4]), FpAdd_8U_23U_and_59_ssc);
  assign FpAlu_8U_23U_nor_14_nl = ~(MUX_v_4_2_2((FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_13_nl),
      4'b1111, FpAdd_8U_23U_and_117_ssc));
  assign FpAlu_8U_23U_FpAlu_8U_23U_nor_14_nl = ~(MUX_v_4_2_2((FpAlu_8U_23U_nor_14_nl),
      4'b1111, FpAlu_8U_23U_equal_tmp_237));
  assign and_4113_nl = nor_7_ssc & (~(or_dcpl_1057 | and_dcpl_1812));
  assign FpAlu_8U_23U_mux1h_1030_nl = MUX1HOT_v_22_3_2((FpAdd_8U_23U_o_mant_4_lpi_1_dfm_2_mx0[22:1]),
      (FpCmp_8U_23U_true_o_22_0_4_lpi_1_dfm_6[22:1]), (FpCmp_8U_23U_false_o_22_0_4_lpi_1_dfm_6[22:1]),
      {FpAlu_8U_23U_nor_dfs_79 , FpAlu_8U_23U_equal_tmp_235 , FpAlu_8U_23U_equal_tmp_239});
  assign FpAlu_8U_23U_not_86_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_15_nl = MUX_v_22_2_2(22'b0000000000000000000000, (FpAlu_8U_23U_mux1h_1030_nl),
      (FpAlu_8U_23U_not_86_nl));
  assign FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_12_nl = MUX_v_4_2_2(FpAdd_8U_23U_o_expo_4_lpi_1_dfm_2_7_4,
      (FpAdd_8U_23U_o_expo_4_sva_4[7:4]), FpAdd_8U_23U_and_63_ssc);
  assign FpAlu_8U_23U_nor_13_nl = ~(MUX_v_4_2_2((FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_12_nl),
      4'b1111, FpAdd_8U_23U_and_119_ssc));
  assign FpAlu_8U_23U_FpAlu_8U_23U_nor_13_nl = ~(MUX_v_4_2_2((FpAlu_8U_23U_nor_13_nl),
      4'b1111, FpAlu_8U_23U_equal_tmp_237));
  assign and_4107_nl = nor_7_ssc & (~(or_dcpl_1062 | and_dcpl_1820));
  assign FpAlu_8U_23U_mux1h_1027_nl = MUX1HOT_v_22_3_2((FpAdd_8U_23U_o_mant_5_lpi_1_dfm_2_mx0[22:1]),
      (FpCmp_8U_23U_true_o_22_0_5_lpi_1_dfm_6[22:1]), (FpCmp_8U_23U_false_o_22_0_5_lpi_1_dfm_6[22:1]),
      {FpAlu_8U_23U_nor_dfs_79 , FpAlu_8U_23U_equal_tmp_235 , FpAlu_8U_23U_equal_tmp_239});
  assign FpAlu_8U_23U_not_88_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_19_nl = MUX_v_22_2_2(22'b0000000000000000000000, (FpAlu_8U_23U_mux1h_1027_nl),
      (FpAlu_8U_23U_not_88_nl));
  assign FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_11_nl = MUX_v_4_2_2(FpAdd_8U_23U_o_expo_5_lpi_1_dfm_2_7_4,
      (FpAdd_8U_23U_o_expo_5_sva_4[7:4]), FpAdd_8U_23U_and_67_ssc);
  assign FpAlu_8U_23U_nor_12_nl = ~(MUX_v_4_2_2((FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_11_nl),
      4'b1111, FpAdd_8U_23U_and_121_ssc));
  assign FpAlu_8U_23U_FpAlu_8U_23U_nor_12_nl = ~(MUX_v_4_2_2((FpAlu_8U_23U_nor_12_nl),
      4'b1111, FpAlu_8U_23U_equal_tmp_237));
  assign and_4101_nl = nor_7_ssc & (~(or_dcpl_1067 | and_dcpl_1828));
  assign FpAlu_8U_23U_mux1h_292_nl = MUX1HOT_v_22_3_2((FpAdd_8U_23U_o_mant_6_lpi_1_dfm_2_mx0[22:1]),
      (FpCmp_8U_23U_true_o_22_0_6_lpi_1_dfm_6[22:1]), (FpCmp_8U_23U_false_o_22_0_6_lpi_1_dfm_6[22:1]),
      {FpAlu_8U_23U_nor_dfs_79 , FpAlu_8U_23U_equal_tmp_235 , FpAlu_8U_23U_equal_tmp_239});
  assign FpAlu_8U_23U_not_90_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_23_nl = MUX_v_22_2_2(22'b0000000000000000000000, (FpAlu_8U_23U_mux1h_292_nl),
      (FpAlu_8U_23U_not_90_nl));
  assign FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_10_nl = MUX_v_4_2_2(FpAdd_8U_23U_o_expo_6_lpi_1_dfm_2_7_4,
      (FpAdd_8U_23U_o_expo_6_sva_4[7:4]), FpAdd_8U_23U_and_71_ssc);
  assign FpAlu_8U_23U_nor_11_nl = ~(MUX_v_4_2_2((FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_10_nl),
      4'b1111, FpAdd_8U_23U_and_123_ssc));
  assign FpAlu_8U_23U_FpAlu_8U_23U_nor_11_nl = ~(MUX_v_4_2_2((FpAlu_8U_23U_nor_11_nl),
      4'b1111, FpAlu_8U_23U_equal_tmp_237));
  assign and_4095_nl = nor_7_ssc & (~(or_dcpl_1072 | and_dcpl_1836));
  assign FpAlu_8U_23U_mux1h_344_nl = MUX1HOT_v_22_3_2((FpAdd_8U_23U_o_mant_7_lpi_1_dfm_2_mx0[22:1]),
      (FpCmp_8U_23U_true_o_22_0_7_lpi_1_dfm_6[22:1]), (FpCmp_8U_23U_false_o_22_0_7_lpi_1_dfm_6[22:1]),
      {FpAlu_8U_23U_nor_dfs_79 , FpAlu_8U_23U_equal_tmp_235 , FpAlu_8U_23U_equal_tmp_239});
  assign FpAlu_8U_23U_not_92_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_27_nl = MUX_v_22_2_2(22'b0000000000000000000000, (FpAlu_8U_23U_mux1h_344_nl),
      (FpAlu_8U_23U_not_92_nl));
  assign FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_9_nl = MUX_v_4_2_2(FpAdd_8U_23U_o_expo_7_lpi_1_dfm_2_7_4,
      (FpAdd_8U_23U_o_expo_7_sva_4[7:4]), FpAdd_8U_23U_and_75_ssc);
  assign FpAlu_8U_23U_nor_10_nl = ~(MUX_v_4_2_2((FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_9_nl),
      4'b1111, FpAdd_8U_23U_and_125_ssc));
  assign FpAlu_8U_23U_FpAlu_8U_23U_nor_10_nl = ~(MUX_v_4_2_2((FpAlu_8U_23U_nor_10_nl),
      4'b1111, FpAlu_8U_23U_equal_tmp_237));
  assign and_4089_nl = nor_7_ssc & (~(or_dcpl_1077 | and_dcpl_1844));
  assign FpAlu_8U_23U_mux1h_396_nl = MUX1HOT_v_22_3_2((FpAdd_8U_23U_o_mant_8_lpi_1_dfm_2_mx0[22:1]),
      (FpCmp_8U_23U_true_o_22_0_8_lpi_1_dfm_6[22:1]), (FpCmp_8U_23U_false_o_22_0_8_lpi_1_dfm_6[22:1]),
      {FpAlu_8U_23U_nor_dfs_79 , FpAlu_8U_23U_equal_tmp_235 , FpAlu_8U_23U_equal_tmp_239});
  assign FpAlu_8U_23U_not_94_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_31_nl = MUX_v_22_2_2(22'b0000000000000000000000, (FpAlu_8U_23U_mux1h_396_nl),
      (FpAlu_8U_23U_not_94_nl));
  assign FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_8_nl = MUX_v_4_2_2(FpAdd_8U_23U_o_expo_8_lpi_1_dfm_2_7_4,
      (FpAdd_8U_23U_o_expo_8_sva_4[7:4]), FpAdd_8U_23U_and_79_ssc);
  assign FpAlu_8U_23U_nor_9_nl = ~(MUX_v_4_2_2((FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_8_nl),
      4'b1111, FpAdd_8U_23U_and_127_ssc));
  assign FpAlu_8U_23U_FpAlu_8U_23U_nor_9_nl = ~(MUX_v_4_2_2((FpAlu_8U_23U_nor_9_nl),
      4'b1111, FpAlu_8U_23U_equal_tmp_237));
  assign and_4083_nl = nor_7_ssc & (~(or_dcpl_1082 | and_dcpl_1852));
  assign FpAlu_8U_23U_mux1h_448_nl = MUX1HOT_v_22_3_2((FpAdd_8U_23U_o_mant_9_lpi_1_dfm_2_mx0[22:1]),
      (FpCmp_8U_23U_true_o_22_0_9_lpi_1_dfm_6[22:1]), (FpCmp_8U_23U_false_o_22_0_9_lpi_1_dfm_6[22:1]),
      {FpAlu_8U_23U_nor_dfs_79 , FpAlu_8U_23U_equal_tmp_235 , FpAlu_8U_23U_equal_tmp_239});
  assign FpAlu_8U_23U_not_96_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_35_nl = MUX_v_22_2_2(22'b0000000000000000000000, (FpAlu_8U_23U_mux1h_448_nl),
      (FpAlu_8U_23U_not_96_nl));
  assign FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_7_nl = MUX_v_4_2_2(FpAdd_8U_23U_o_expo_9_lpi_1_dfm_2_7_4,
      (FpAdd_8U_23U_o_expo_9_sva_4[7:4]), FpAdd_8U_23U_and_83_ssc);
  assign FpAlu_8U_23U_nor_8_nl = ~(MUX_v_4_2_2((FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_7_nl),
      4'b1111, FpAdd_8U_23U_and_129_ssc));
  assign FpAlu_8U_23U_FpAlu_8U_23U_nor_8_nl = ~(MUX_v_4_2_2((FpAlu_8U_23U_nor_8_nl),
      4'b1111, FpAlu_8U_23U_equal_tmp_237));
  assign and_4077_nl = nor_7_ssc & (~(or_dcpl_1087 | and_dcpl_1860));
  assign FpAlu_8U_23U_mux1h_500_nl = MUX1HOT_v_22_3_2((FpAdd_8U_23U_o_mant_10_lpi_1_dfm_2_mx0[22:1]),
      (FpCmp_8U_23U_true_o_22_0_10_lpi_1_dfm_6[22:1]), (FpCmp_8U_23U_false_o_22_0_10_lpi_1_dfm_6[22:1]),
      {FpAlu_8U_23U_nor_dfs_79 , FpAlu_8U_23U_equal_tmp_235 , FpAlu_8U_23U_equal_tmp_239});
  assign FpAlu_8U_23U_not_98_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_39_nl = MUX_v_22_2_2(22'b0000000000000000000000, (FpAlu_8U_23U_mux1h_500_nl),
      (FpAlu_8U_23U_not_98_nl));
  assign FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_6_nl = MUX_v_4_2_2(FpAdd_8U_23U_o_expo_10_lpi_1_dfm_2_7_4,
      (FpAdd_8U_23U_o_expo_10_sva_4[7:4]), FpAdd_8U_23U_and_87_ssc);
  assign FpAlu_8U_23U_nor_7_nl = ~(MUX_v_4_2_2((FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_6_nl),
      4'b1111, FpAdd_8U_23U_and_131_ssc));
  assign FpAlu_8U_23U_FpAlu_8U_23U_nor_7_nl = ~(MUX_v_4_2_2((FpAlu_8U_23U_nor_7_nl),
      4'b1111, FpAlu_8U_23U_equal_tmp_237));
  assign and_4071_nl = nor_7_ssc & (~(or_dcpl_1092 | and_dcpl_1868));
  assign FpAlu_8U_23U_mux1h_552_nl = MUX1HOT_v_22_3_2((FpAdd_8U_23U_o_mant_11_lpi_1_dfm_2_mx0[22:1]),
      (FpCmp_8U_23U_true_o_22_0_11_lpi_1_dfm_6[22:1]), (FpCmp_8U_23U_false_o_22_0_11_lpi_1_dfm_6[22:1]),
      {FpAlu_8U_23U_nor_dfs_79 , FpAlu_8U_23U_equal_tmp_235 , FpAlu_8U_23U_equal_tmp_239});
  assign FpAlu_8U_23U_not_100_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_43_nl = MUX_v_22_2_2(22'b0000000000000000000000, (FpAlu_8U_23U_mux1h_552_nl),
      (FpAlu_8U_23U_not_100_nl));
  assign FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_5_nl = MUX_v_4_2_2(FpAdd_8U_23U_o_expo_11_lpi_1_dfm_2_7_4,
      (FpAdd_8U_23U_o_expo_11_sva_4[7:4]), FpAdd_8U_23U_and_91_ssc);
  assign FpAlu_8U_23U_nor_6_nl = ~(MUX_v_4_2_2((FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_5_nl),
      4'b1111, FpAdd_8U_23U_and_133_ssc));
  assign FpAlu_8U_23U_FpAlu_8U_23U_nor_6_nl = ~(MUX_v_4_2_2((FpAlu_8U_23U_nor_6_nl),
      4'b1111, FpAlu_8U_23U_equal_tmp_237));
  assign and_4065_nl = nor_7_ssc & (~(or_dcpl_1097 | and_dcpl_1876));
  assign FpAlu_8U_23U_mux1h_604_nl = MUX1HOT_v_22_3_2((FpAdd_8U_23U_o_mant_12_lpi_1_dfm_2_mx0[22:1]),
      (FpCmp_8U_23U_true_o_22_0_12_lpi_1_dfm_6[22:1]), (FpCmp_8U_23U_false_o_22_0_12_lpi_1_dfm_6[22:1]),
      {FpAlu_8U_23U_nor_dfs_79 , FpAlu_8U_23U_equal_tmp_235 , FpAlu_8U_23U_equal_tmp_239});
  assign FpAlu_8U_23U_not_102_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_47_nl = MUX_v_22_2_2(22'b0000000000000000000000, (FpAlu_8U_23U_mux1h_604_nl),
      (FpAlu_8U_23U_not_102_nl));
  assign FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_4_nl = MUX_v_4_2_2(FpAdd_8U_23U_o_expo_12_lpi_1_dfm_2_7_4,
      (FpAdd_8U_23U_o_expo_12_sva_4[7:4]), FpAdd_8U_23U_and_95_ssc);
  assign FpAlu_8U_23U_nor_5_nl = ~(MUX_v_4_2_2((FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_4_nl),
      4'b1111, FpAdd_8U_23U_and_135_ssc));
  assign FpAlu_8U_23U_FpAlu_8U_23U_nor_5_nl = ~(MUX_v_4_2_2((FpAlu_8U_23U_nor_5_nl),
      4'b1111, FpAlu_8U_23U_equal_tmp_237));
  assign and_4059_nl = nor_7_ssc & (~(or_dcpl_1102 | and_dcpl_1884));
  assign FpAlu_8U_23U_mux1h_656_nl = MUX1HOT_v_22_3_2((FpAdd_8U_23U_o_mant_13_lpi_1_dfm_2_mx0[22:1]),
      (FpCmp_8U_23U_true_o_22_0_13_lpi_1_dfm_6[22:1]), (FpCmp_8U_23U_false_o_22_0_13_lpi_1_dfm_6[22:1]),
      {FpAlu_8U_23U_nor_dfs_79 , FpAlu_8U_23U_equal_tmp_235 , FpAlu_8U_23U_equal_tmp_239});
  assign FpAlu_8U_23U_not_104_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_51_nl = MUX_v_22_2_2(22'b0000000000000000000000, (FpAlu_8U_23U_mux1h_656_nl),
      (FpAlu_8U_23U_not_104_nl));
  assign FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_3_nl = MUX_v_4_2_2(FpAdd_8U_23U_o_expo_13_lpi_1_dfm_2_7_4,
      (FpAdd_8U_23U_o_expo_13_sva_4[7:4]), FpAdd_8U_23U_and_99_ssc);
  assign FpAlu_8U_23U_nor_4_nl = ~(MUX_v_4_2_2((FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_3_nl),
      4'b1111, FpAdd_8U_23U_and_137_ssc));
  assign FpAlu_8U_23U_FpAlu_8U_23U_nor_4_nl = ~(MUX_v_4_2_2((FpAlu_8U_23U_nor_4_nl),
      4'b1111, FpAlu_8U_23U_equal_tmp_237));
  assign and_4053_nl = nor_7_ssc & (~(or_dcpl_1107 | and_dcpl_1892));
  assign FpAlu_8U_23U_mux1h_708_nl = MUX1HOT_v_22_3_2((FpAdd_8U_23U_o_mant_14_lpi_1_dfm_2_mx0[22:1]),
      (FpCmp_8U_23U_true_o_22_0_14_lpi_1_dfm_6[22:1]), (FpCmp_8U_23U_false_o_22_0_14_lpi_1_dfm_6[22:1]),
      {FpAlu_8U_23U_nor_dfs_79 , FpAlu_8U_23U_equal_tmp_235 , FpAlu_8U_23U_equal_tmp_239});
  assign FpAlu_8U_23U_not_106_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_55_nl = MUX_v_22_2_2(22'b0000000000000000000000, (FpAlu_8U_23U_mux1h_708_nl),
      (FpAlu_8U_23U_not_106_nl));
  assign FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_2_nl = MUX_v_4_2_2(FpAdd_8U_23U_o_expo_14_lpi_1_dfm_2_7_4,
      (FpAdd_8U_23U_o_expo_14_sva_4[7:4]), FpAdd_8U_23U_and_103_ssc);
  assign FpAlu_8U_23U_nor_3_nl = ~(MUX_v_4_2_2((FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_2_nl),
      4'b1111, FpAdd_8U_23U_and_139_ssc));
  assign FpAlu_8U_23U_FpAlu_8U_23U_nor_3_nl = ~(MUX_v_4_2_2((FpAlu_8U_23U_nor_3_nl),
      4'b1111, FpAlu_8U_23U_equal_tmp_237));
  assign and_4047_nl = nor_7_ssc & (~(or_dcpl_1112 | and_dcpl_1900));
  assign FpAlu_8U_23U_mux1h_760_nl = MUX1HOT_v_22_3_2((FpAdd_8U_23U_o_mant_15_lpi_1_dfm_2_mx0[22:1]),
      (FpCmp_8U_23U_true_o_22_0_15_lpi_1_dfm_6[22:1]), (FpCmp_8U_23U_false_o_22_0_15_lpi_1_dfm_6[22:1]),
      {FpAlu_8U_23U_nor_dfs_79 , FpAlu_8U_23U_equal_tmp_235 , FpAlu_8U_23U_equal_tmp_239});
  assign FpAlu_8U_23U_not_108_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_59_nl = MUX_v_22_2_2(22'b0000000000000000000000, (FpAlu_8U_23U_mux1h_760_nl),
      (FpAlu_8U_23U_not_108_nl));
  assign FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_1_nl = MUX_v_4_2_2(FpAdd_8U_23U_o_expo_15_lpi_1_dfm_2_7_4,
      (FpAdd_8U_23U_o_expo_15_sva_4[7:4]), FpAdd_8U_23U_and_107_ssc);
  assign FpAlu_8U_23U_nor_2_nl = ~(MUX_v_4_2_2((FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_1_nl),
      4'b1111, FpAdd_8U_23U_and_141_ssc));
  assign FpAlu_8U_23U_FpAlu_8U_23U_nor_2_nl = ~(MUX_v_4_2_2((FpAlu_8U_23U_nor_2_nl),
      4'b1111, FpAlu_8U_23U_equal_tmp_237));
  assign and_4041_nl = nor_7_ssc & (~(or_dcpl_1117 | and_dcpl_1908));
  assign FpAlu_8U_23U_mux1h_1004_nl = MUX1HOT_v_22_3_2((FpAdd_8U_23U_o_mant_lpi_1_dfm_2_mx0[22:1]),
      (FpCmp_8U_23U_true_o_22_0_lpi_1_dfm_6[22:1]), (FpCmp_8U_23U_false_o_22_0_lpi_1_dfm_6[22:1]),
      {FpAlu_8U_23U_nor_dfs_79 , FpAlu_8U_23U_equal_tmp_235 , FpAlu_8U_23U_equal_tmp_239});
  assign FpAlu_8U_23U_not_110_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_63_nl = MUX_v_22_2_2(22'b0000000000000000000000, (FpAlu_8U_23U_mux1h_1004_nl),
      (FpAlu_8U_23U_not_110_nl));
  assign FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_nl = MUX_v_4_2_2(FpAdd_8U_23U_o_expo_lpi_1_dfm_2_7_4,
      (FpAdd_8U_23U_o_expo_sva_4[7:4]), FpAdd_8U_23U_and_111_ssc);
  assign FpAlu_8U_23U_nor_1_nl = ~(MUX_v_4_2_2((FpAdd_8U_23U_FpAdd_8U_23U_FpAdd_8U_23U_mux_nl),
      4'b1111, FpAdd_8U_23U_and_143_ssc));
  assign FpAlu_8U_23U_FpAlu_8U_23U_nor_1_nl = ~(MUX_v_4_2_2((FpAlu_8U_23U_nor_1_nl),
      4'b1111, FpAlu_8U_23U_equal_tmp_237));
  assign and_4035_nl = nor_7_ssc & (~(or_dcpl_1122 | and_dcpl_1916));
  assign FpAlu_8U_23U_and_610_nl = (~(FpAdd_8U_23U_and_32_tmp | FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0))
      & alu_loop_op_if_alu_loop_op_if_nor_cse & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_611_nl = FpAdd_8U_23U_and_51_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_612_nl = FpAdd_8U_23U_and_113_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_mux1h_1040_nl = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_11,
      FpAdd_8U_23U_o_expo_1_lpi_1_dfm_2_3_0, (FpAdd_8U_23U_o_expo_1_sva_4[3:0]),
      4'b1110, {FpAlu_8U_23U_or_863_cse , (FpAlu_8U_23U_and_610_nl) , (FpAlu_8U_23U_and_611_nl)
      , (FpAlu_8U_23U_and_612_nl)});
  assign FpAlu_8U_23U_not_114_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_2_nl = MUX_v_4_2_2(4'b0000, (FpAlu_8U_23U_mux1h_1040_nl),
      (FpAlu_8U_23U_not_114_nl));
  assign and_4128_nl = nor_7_ssc & (~ or_dcpl_1047);
  assign or_5091_nl = io_read_cfg_alu_bypass_rsc_svs_7 | FpAlu_8U_23U_or_831_itm_4
      | FpAlu_8U_23U_equal_tmp_237 | (cfg_precision!=2'b10) | FpAlu_8U_23U_nor_dfs_79
      | reg_FpAlu_8U_23U_or_752_cse;
  assign nand_nl = ~(((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_1_lpi_1_dfm_10)
      & (cfg_precision[1]) & (~(FpAlu_8U_23U_or_831_itm_4 | FpAlu_8U_23U_equal_tmp_237
      | (cfg_precision[0]))));
  assign mux_1569_nl = MUX_s_1_2_2((nand_nl), (or_5091_nl), or_dcpl_1047);
  assign FpAlu_8U_23U_and_615_nl = (~(FpAdd_8U_23U_and_33_tmp | FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0))
      & alu_loop_op_if_alu_loop_op_if_nor_1_cse & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_616_nl = FpAdd_8U_23U_and_55_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_617_nl = FpAdd_8U_23U_and_115_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_mux1h_1037_nl = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_11,
      FpAdd_8U_23U_o_expo_2_lpi_1_dfm_2_3_0, (FpAdd_8U_23U_o_expo_2_sva_4[3:0]),
      4'b1110, {FpAlu_8U_23U_or_864_cse , (FpAlu_8U_23U_and_615_nl) , (FpAlu_8U_23U_and_616_nl)
      , (FpAlu_8U_23U_and_617_nl)});
  assign FpAlu_8U_23U_not_115_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_6_nl = MUX_v_4_2_2(4'b0000, (FpAlu_8U_23U_mux1h_1037_nl),
      (FpAlu_8U_23U_not_115_nl));
  assign and_4122_nl = nor_7_ssc & (~ or_dcpl_1052);
  assign or_5097_nl = io_read_cfg_alu_bypass_rsc_svs_7 | FpAlu_8U_23U_or_833_itm_4
      | FpAlu_8U_23U_equal_tmp_237 | (cfg_precision!=2'b10) | FpAlu_8U_23U_nor_dfs_79
      | reg_FpAlu_8U_23U_or_755_cse;
  assign nand_429_nl = ~(((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_2_lpi_1_dfm_10)
      & (cfg_precision[1]) & (~(FpAlu_8U_23U_or_833_itm_4 | FpAlu_8U_23U_equal_tmp_237
      | (cfg_precision[0]))));
  assign mux_1572_nl = MUX_s_1_2_2((nand_429_nl), (or_5097_nl), or_dcpl_1052);
  assign FpAlu_8U_23U_and_620_nl = (~(FpAdd_8U_23U_and_34_tmp | FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0))
      & alu_loop_op_if_alu_loop_op_if_nor_2_cse & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_621_nl = FpAdd_8U_23U_and_59_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_622_nl = FpAdd_8U_23U_and_117_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_mux1h_1034_nl = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_11,
      FpAdd_8U_23U_o_expo_3_lpi_1_dfm_2_3_0, (FpAdd_8U_23U_o_expo_3_sva_4[3:0]),
      4'b1110, {FpAlu_8U_23U_or_865_cse , (FpAlu_8U_23U_and_620_nl) , (FpAlu_8U_23U_and_621_nl)
      , (FpAlu_8U_23U_and_622_nl)});
  assign FpAlu_8U_23U_not_116_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_10_nl = MUX_v_4_2_2(4'b0000, (FpAlu_8U_23U_mux1h_1034_nl),
      (FpAlu_8U_23U_not_116_nl));
  assign and_4116_nl = nor_7_ssc & (~ or_dcpl_1057);
  assign or_5103_nl = io_read_cfg_alu_bypass_rsc_svs_7 | FpAlu_8U_23U_or_835_itm_4
      | FpAlu_8U_23U_equal_tmp_237 | (cfg_precision!=2'b10) | FpAlu_8U_23U_nor_dfs_79
      | reg_FpAlu_8U_23U_or_758_cse;
  assign nand_430_nl = ~(((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_3_lpi_1_dfm_10)
      & (cfg_precision[1]) & (~(FpAlu_8U_23U_or_835_itm_4 | FpAlu_8U_23U_equal_tmp_237
      | (cfg_precision[0]))));
  assign mux_1575_nl = MUX_s_1_2_2((nand_430_nl), (or_5103_nl), or_dcpl_1057);
  assign FpAlu_8U_23U_and_625_nl = (~(FpAdd_8U_23U_and_35_tmp | FpAdd_8U_23U_is_inf_4_lpi_1_dfm_2_mx0))
      & alu_loop_op_if_alu_loop_op_if_nor_3_cse & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_626_nl = FpAdd_8U_23U_and_63_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_627_nl = FpAdd_8U_23U_and_119_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_mux1h_1031_nl = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_11,
      FpAdd_8U_23U_o_expo_4_lpi_1_dfm_2_3_0, (FpAdd_8U_23U_o_expo_4_sva_4[3:0]),
      4'b1110, {FpAlu_8U_23U_or_866_cse , (FpAlu_8U_23U_and_625_nl) , (FpAlu_8U_23U_and_626_nl)
      , (FpAlu_8U_23U_and_627_nl)});
  assign FpAlu_8U_23U_not_117_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_14_nl = MUX_v_4_2_2(4'b0000, (FpAlu_8U_23U_mux1h_1031_nl),
      (FpAlu_8U_23U_not_117_nl));
  assign and_4110_nl = nor_7_ssc & (~ or_dcpl_1062);
  assign or_5109_nl = io_read_cfg_alu_bypass_rsc_svs_7 | FpAlu_8U_23U_or_837_itm_4
      | FpAlu_8U_23U_equal_tmp_237 | (cfg_precision!=2'b10) | FpAlu_8U_23U_nor_dfs_79
      | reg_FpAlu_8U_23U_or_761_cse;
  assign nand_431_nl = ~(((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_4_lpi_1_dfm_10)
      & (cfg_precision[1]) & (~(FpAlu_8U_23U_or_837_itm_4 | FpAlu_8U_23U_equal_tmp_237
      | (cfg_precision[0]))));
  assign mux_1578_nl = MUX_s_1_2_2((nand_431_nl), (or_5109_nl), or_dcpl_1062);
  assign FpAlu_8U_23U_and_630_nl = (~(FpAdd_8U_23U_and_36_tmp | FpAdd_8U_23U_is_inf_5_lpi_1_dfm_2_mx0))
      & alu_loop_op_if_alu_loop_op_if_nor_4_cse & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_631_nl = FpAdd_8U_23U_and_67_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_632_nl = FpAdd_8U_23U_and_121_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_mux1h_1028_nl = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_11,
      FpAdd_8U_23U_o_expo_5_lpi_1_dfm_2_3_0, (FpAdd_8U_23U_o_expo_5_sva_4[3:0]),
      4'b1110, {FpAlu_8U_23U_or_867_cse , (FpAlu_8U_23U_and_630_nl) , (FpAlu_8U_23U_and_631_nl)
      , (FpAlu_8U_23U_and_632_nl)});
  assign FpAlu_8U_23U_not_118_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_18_nl = MUX_v_4_2_2(4'b0000, (FpAlu_8U_23U_mux1h_1028_nl),
      (FpAlu_8U_23U_not_118_nl));
  assign and_4104_nl = nor_7_ssc & (~ or_dcpl_1067);
  assign or_5115_nl = io_read_cfg_alu_bypass_rsc_svs_7 | FpAlu_8U_23U_or_839_itm_4
      | FpAlu_8U_23U_equal_tmp_237 | (cfg_precision!=2'b10) | FpAlu_8U_23U_nor_dfs_79
      | reg_FpAlu_8U_23U_or_764_cse;
  assign nand_432_nl = ~(((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_5_lpi_1_dfm_10)
      & (cfg_precision[1]) & (~(FpAlu_8U_23U_or_839_itm_4 | FpAlu_8U_23U_equal_tmp_237
      | (cfg_precision[0]))));
  assign mux_1581_nl = MUX_s_1_2_2((nand_432_nl), (or_5115_nl), or_dcpl_1067);
  assign FpAlu_8U_23U_and_635_nl = (~(FpAdd_8U_23U_and_37_tmp | FpAdd_8U_23U_is_inf_6_lpi_1_dfm_2_mx0))
      & alu_loop_op_if_alu_loop_op_if_nor_5_cse & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_636_nl = FpAdd_8U_23U_and_71_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_637_nl = FpAdd_8U_23U_and_123_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_mux1h_1025_nl = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_11,
      FpAdd_8U_23U_o_expo_6_lpi_1_dfm_2_3_0, (FpAdd_8U_23U_o_expo_6_sva_4[3:0]),
      4'b1110, {FpAlu_8U_23U_or_868_cse , (FpAlu_8U_23U_and_635_nl) , (FpAlu_8U_23U_and_636_nl)
      , (FpAlu_8U_23U_and_637_nl)});
  assign FpAlu_8U_23U_not_119_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_22_nl = MUX_v_4_2_2(4'b0000, (FpAlu_8U_23U_mux1h_1025_nl),
      (FpAlu_8U_23U_not_119_nl));
  assign and_4098_nl = nor_7_ssc & (~ or_dcpl_1072);
  assign or_5121_nl = io_read_cfg_alu_bypass_rsc_svs_7 | FpAlu_8U_23U_or_841_itm_4
      | FpAlu_8U_23U_equal_tmp_237 | (cfg_precision!=2'b10) | FpAlu_8U_23U_nor_dfs_79
      | reg_FpAlu_8U_23U_or_767_cse;
  assign nand_433_nl = ~(((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_6_lpi_1_dfm_10)
      & (cfg_precision[1]) & (~(FpAlu_8U_23U_or_841_itm_4 | FpAlu_8U_23U_equal_tmp_237
      | (cfg_precision[0]))));
  assign mux_1584_nl = MUX_s_1_2_2((nand_433_nl), (or_5121_nl), or_dcpl_1072);
  assign FpAlu_8U_23U_and_640_nl = (~(FpAdd_8U_23U_and_38_tmp | FpAdd_8U_23U_is_inf_7_lpi_1_dfm_2_mx0))
      & alu_loop_op_if_alu_loop_op_if_nor_6_cse & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_641_nl = FpAdd_8U_23U_and_75_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_642_nl = FpAdd_8U_23U_and_125_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_mux1h_1023_nl = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_11,
      FpAdd_8U_23U_o_expo_7_lpi_1_dfm_2_3_0, (FpAdd_8U_23U_o_expo_7_sva_4[3:0]),
      4'b1110, {FpAlu_8U_23U_or_869_cse , (FpAlu_8U_23U_and_640_nl) , (FpAlu_8U_23U_and_641_nl)
      , (FpAlu_8U_23U_and_642_nl)});
  assign FpAlu_8U_23U_not_120_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_26_nl = MUX_v_4_2_2(4'b0000, (FpAlu_8U_23U_mux1h_1023_nl),
      (FpAlu_8U_23U_not_120_nl));
  assign and_4092_nl = nor_7_ssc & (~ or_dcpl_1077);
  assign or_5127_nl = io_read_cfg_alu_bypass_rsc_svs_7 | FpAlu_8U_23U_or_843_itm_4
      | FpAlu_8U_23U_equal_tmp_237 | (cfg_precision!=2'b10) | FpAlu_8U_23U_nor_dfs_79
      | reg_FpAlu_8U_23U_or_770_cse;
  assign nand_434_nl = ~(((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_7_lpi_1_dfm_10)
      & (cfg_precision[1]) & (~(FpAlu_8U_23U_or_843_itm_4 | FpAlu_8U_23U_equal_tmp_237
      | (cfg_precision[0]))));
  assign mux_1587_nl = MUX_s_1_2_2((nand_434_nl), (or_5127_nl), or_dcpl_1077);
  assign FpAlu_8U_23U_and_645_nl = (~(FpAdd_8U_23U_and_39_tmp | FpAdd_8U_23U_is_inf_8_lpi_1_dfm_2_mx0))
      & alu_loop_op_if_alu_loop_op_if_nor_7_cse & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_646_nl = FpAdd_8U_23U_and_79_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_647_nl = FpAdd_8U_23U_and_127_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_mux1h_1021_nl = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_11,
      FpAdd_8U_23U_o_expo_8_lpi_1_dfm_2_3_0, (FpAdd_8U_23U_o_expo_8_sva_4[3:0]),
      4'b1110, {FpAlu_8U_23U_or_870_cse , (FpAlu_8U_23U_and_645_nl) , (FpAlu_8U_23U_and_646_nl)
      , (FpAlu_8U_23U_and_647_nl)});
  assign FpAlu_8U_23U_not_121_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_30_nl = MUX_v_4_2_2(4'b0000, (FpAlu_8U_23U_mux1h_1021_nl),
      (FpAlu_8U_23U_not_121_nl));
  assign and_4086_nl = nor_7_ssc & (~ or_dcpl_1082);
  assign or_5133_nl = io_read_cfg_alu_bypass_rsc_svs_7 | FpAlu_8U_23U_or_845_itm_4
      | FpAlu_8U_23U_equal_tmp_237 | (cfg_precision!=2'b10) | FpAlu_8U_23U_nor_dfs_79
      | reg_FpAlu_8U_23U_or_773_cse;
  assign nand_435_nl = ~(((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_8_lpi_1_dfm_10)
      & (cfg_precision[1]) & (~(FpAlu_8U_23U_or_845_itm_4 | FpAlu_8U_23U_equal_tmp_237
      | (cfg_precision[0]))));
  assign mux_1590_nl = MUX_s_1_2_2((nand_435_nl), (or_5133_nl), or_dcpl_1082);
  assign FpAlu_8U_23U_and_650_nl = (~(FpAdd_8U_23U_and_40_tmp | FpAdd_8U_23U_is_inf_9_lpi_1_dfm_2_mx0))
      & alu_loop_op_if_alu_loop_op_if_nor_8_cse & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_651_nl = FpAdd_8U_23U_and_83_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_652_nl = FpAdd_8U_23U_and_129_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_mux1h_1019_nl = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_11,
      FpAdd_8U_23U_o_expo_9_lpi_1_dfm_2_3_0, (FpAdd_8U_23U_o_expo_9_sva_4[3:0]),
      4'b1110, {FpAlu_8U_23U_or_871_cse , (FpAlu_8U_23U_and_650_nl) , (FpAlu_8U_23U_and_651_nl)
      , (FpAlu_8U_23U_and_652_nl)});
  assign FpAlu_8U_23U_not_122_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_34_nl = MUX_v_4_2_2(4'b0000, (FpAlu_8U_23U_mux1h_1019_nl),
      (FpAlu_8U_23U_not_122_nl));
  assign and_4080_nl = nor_7_ssc & (~ or_dcpl_1087);
  assign or_5139_nl = io_read_cfg_alu_bypass_rsc_svs_7 | FpAlu_8U_23U_or_847_itm_4
      | FpAlu_8U_23U_equal_tmp_237 | (cfg_precision!=2'b10) | FpAlu_8U_23U_nor_dfs_79
      | reg_FpAlu_8U_23U_or_776_cse;
  assign nand_436_nl = ~(((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_9_lpi_1_dfm_10)
      & (cfg_precision[1]) & (~(FpAlu_8U_23U_or_847_itm_4 | FpAlu_8U_23U_equal_tmp_237
      | (cfg_precision[0]))));
  assign mux_1593_nl = MUX_s_1_2_2((nand_436_nl), (or_5139_nl), or_dcpl_1087);
  assign FpAlu_8U_23U_and_655_nl = (~(FpAdd_8U_23U_and_41_tmp | FpAdd_8U_23U_is_inf_10_lpi_1_dfm_2_mx0))
      & alu_loop_op_if_alu_loop_op_if_nor_9_cse & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_656_nl = FpAdd_8U_23U_and_87_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_657_nl = FpAdd_8U_23U_and_131_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_mux1h_1017_nl = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_11,
      FpAdd_8U_23U_o_expo_10_lpi_1_dfm_2_3_0, (FpAdd_8U_23U_o_expo_10_sva_4[3:0]),
      4'b1110, {FpAlu_8U_23U_or_872_cse , (FpAlu_8U_23U_and_655_nl) , (FpAlu_8U_23U_and_656_nl)
      , (FpAlu_8U_23U_and_657_nl)});
  assign FpAlu_8U_23U_not_123_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_38_nl = MUX_v_4_2_2(4'b0000, (FpAlu_8U_23U_mux1h_1017_nl),
      (FpAlu_8U_23U_not_123_nl));
  assign and_4074_nl = nor_7_ssc & (~ or_dcpl_1092);
  assign or_5145_nl = io_read_cfg_alu_bypass_rsc_svs_7 | FpAlu_8U_23U_or_849_itm_4
      | FpAlu_8U_23U_equal_tmp_237 | (cfg_precision!=2'b10) | FpAlu_8U_23U_nor_dfs_79
      | reg_FpAlu_8U_23U_or_779_cse;
  assign nand_437_nl = ~(((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_10_lpi_1_dfm_10)
      & (cfg_precision[1]) & (~(FpAlu_8U_23U_or_849_itm_4 | FpAlu_8U_23U_equal_tmp_237
      | (cfg_precision[0]))));
  assign mux_1596_nl = MUX_s_1_2_2((nand_437_nl), (or_5145_nl), or_dcpl_1092);
  assign FpAlu_8U_23U_and_660_nl = (~(FpAdd_8U_23U_and_42_tmp | FpAdd_8U_23U_is_inf_11_lpi_1_dfm_2_mx0))
      & alu_loop_op_if_alu_loop_op_if_nor_10_cse & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_661_nl = FpAdd_8U_23U_and_91_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_662_nl = FpAdd_8U_23U_and_133_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_mux1h_1015_nl = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_11,
      FpAdd_8U_23U_o_expo_11_lpi_1_dfm_2_3_0, (FpAdd_8U_23U_o_expo_11_sva_4[3:0]),
      4'b1110, {FpAlu_8U_23U_or_873_cse , (FpAlu_8U_23U_and_660_nl) , (FpAlu_8U_23U_and_661_nl)
      , (FpAlu_8U_23U_and_662_nl)});
  assign FpAlu_8U_23U_not_124_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_42_nl = MUX_v_4_2_2(4'b0000, (FpAlu_8U_23U_mux1h_1015_nl),
      (FpAlu_8U_23U_not_124_nl));
  assign and_4068_nl = nor_7_ssc & (~ or_dcpl_1097);
  assign or_5151_nl = io_read_cfg_alu_bypass_rsc_svs_7 | FpAlu_8U_23U_or_851_itm_4
      | FpAlu_8U_23U_equal_tmp_237 | (cfg_precision!=2'b10) | FpAlu_8U_23U_nor_dfs_79
      | reg_FpAlu_8U_23U_or_782_cse;
  assign nand_438_nl = ~(((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_11_lpi_1_dfm_10)
      & (cfg_precision[1]) & (~(FpAlu_8U_23U_or_851_itm_4 | FpAlu_8U_23U_equal_tmp_237
      | (cfg_precision[0]))));
  assign mux_1599_nl = MUX_s_1_2_2((nand_438_nl), (or_5151_nl), or_dcpl_1097);
  assign FpAlu_8U_23U_and_665_nl = (~(FpAdd_8U_23U_and_43_tmp | FpAdd_8U_23U_is_inf_12_lpi_1_dfm_2_mx0))
      & alu_loop_op_if_alu_loop_op_if_nor_11_cse & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_666_nl = FpAdd_8U_23U_and_95_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_667_nl = FpAdd_8U_23U_and_135_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_mux1h_1013_nl = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_11,
      FpAdd_8U_23U_o_expo_12_lpi_1_dfm_2_3_0, (FpAdd_8U_23U_o_expo_12_sva_4[3:0]),
      4'b1110, {FpAlu_8U_23U_or_874_cse , (FpAlu_8U_23U_and_665_nl) , (FpAlu_8U_23U_and_666_nl)
      , (FpAlu_8U_23U_and_667_nl)});
  assign FpAlu_8U_23U_not_125_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_46_nl = MUX_v_4_2_2(4'b0000, (FpAlu_8U_23U_mux1h_1013_nl),
      (FpAlu_8U_23U_not_125_nl));
  assign and_4062_nl = nor_7_ssc & (~ or_dcpl_1102);
  assign or_5157_nl = io_read_cfg_alu_bypass_rsc_svs_7 | FpAlu_8U_23U_or_853_itm_4
      | FpAlu_8U_23U_equal_tmp_237 | (cfg_precision!=2'b10) | FpAlu_8U_23U_nor_dfs_79
      | reg_FpAlu_8U_23U_or_785_cse;
  assign nand_439_nl = ~(((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_12_lpi_1_dfm_10)
      & (cfg_precision[1]) & (~(FpAlu_8U_23U_or_853_itm_4 | FpAlu_8U_23U_equal_tmp_237
      | (cfg_precision[0]))));
  assign mux_1602_nl = MUX_s_1_2_2((nand_439_nl), (or_5157_nl), or_dcpl_1102);
  assign FpAlu_8U_23U_and_670_nl = (~(FpAdd_8U_23U_and_44_tmp | FpAdd_8U_23U_is_inf_13_lpi_1_dfm_2_mx0))
      & alu_loop_op_if_alu_loop_op_if_nor_12_cse & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_671_nl = FpAdd_8U_23U_and_99_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_672_nl = FpAdd_8U_23U_and_137_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_mux1h_1011_nl = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_11,
      FpAdd_8U_23U_o_expo_13_lpi_1_dfm_2_3_0, (FpAdd_8U_23U_o_expo_13_sva_4[3:0]),
      4'b1110, {FpAlu_8U_23U_or_875_cse , (FpAlu_8U_23U_and_670_nl) , (FpAlu_8U_23U_and_671_nl)
      , (FpAlu_8U_23U_and_672_nl)});
  assign FpAlu_8U_23U_not_126_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_50_nl = MUX_v_4_2_2(4'b0000, (FpAlu_8U_23U_mux1h_1011_nl),
      (FpAlu_8U_23U_not_126_nl));
  assign and_4056_nl = nor_7_ssc & (~ or_dcpl_1107);
  assign or_5163_nl = io_read_cfg_alu_bypass_rsc_svs_7 | FpAlu_8U_23U_or_855_itm_4
      | FpAlu_8U_23U_equal_tmp_237 | (cfg_precision!=2'b10) | FpAlu_8U_23U_nor_dfs_79
      | reg_FpAlu_8U_23U_or_788_cse;
  assign nand_440_nl = ~(((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_13_lpi_1_dfm_10)
      & (cfg_precision[1]) & (~(FpAlu_8U_23U_or_855_itm_4 | FpAlu_8U_23U_equal_tmp_237
      | (cfg_precision[0]))));
  assign mux_1605_nl = MUX_s_1_2_2((nand_440_nl), (or_5163_nl), or_dcpl_1107);
  assign FpAlu_8U_23U_and_675_nl = (~(FpAdd_8U_23U_and_45_tmp | FpAdd_8U_23U_is_inf_14_lpi_1_dfm_2_mx0))
      & alu_loop_op_if_alu_loop_op_if_nor_13_cse & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_676_nl = FpAdd_8U_23U_and_103_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_677_nl = FpAdd_8U_23U_and_139_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_mux1h_1009_nl = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_11,
      FpAdd_8U_23U_o_expo_14_lpi_1_dfm_2_3_0, (FpAdd_8U_23U_o_expo_14_sva_4[3:0]),
      4'b1110, {FpAlu_8U_23U_or_876_cse , (FpAlu_8U_23U_and_675_nl) , (FpAlu_8U_23U_and_676_nl)
      , (FpAlu_8U_23U_and_677_nl)});
  assign FpAlu_8U_23U_not_127_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_54_nl = MUX_v_4_2_2(4'b0000, (FpAlu_8U_23U_mux1h_1009_nl),
      (FpAlu_8U_23U_not_127_nl));
  assign and_4050_nl = nor_7_ssc & (~ or_dcpl_1112);
  assign or_5169_nl = io_read_cfg_alu_bypass_rsc_svs_7 | FpAlu_8U_23U_or_857_itm_4
      | FpAlu_8U_23U_equal_tmp_237 | (cfg_precision!=2'b10) | FpAlu_8U_23U_nor_dfs_79
      | reg_FpAlu_8U_23U_or_791_cse;
  assign nand_441_nl = ~(((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_14_lpi_1_dfm_10)
      & (cfg_precision[1]) & (~(FpAlu_8U_23U_or_857_itm_4 | FpAlu_8U_23U_equal_tmp_237
      | (cfg_precision[0]))));
  assign mux_1608_nl = MUX_s_1_2_2((nand_441_nl), (or_5169_nl), or_dcpl_1112);
  assign FpAlu_8U_23U_and_680_nl = (~(FpAdd_8U_23U_and_46_tmp | FpAdd_8U_23U_is_inf_15_lpi_1_dfm_2_mx0))
      & alu_loop_op_if_alu_loop_op_if_nor_14_cse & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_681_nl = FpAdd_8U_23U_and_107_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_682_nl = FpAdd_8U_23U_and_141_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_mux1h_1007_nl = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_11,
      FpAdd_8U_23U_o_expo_15_lpi_1_dfm_2_3_0, (FpAdd_8U_23U_o_expo_15_sva_4[3:0]),
      4'b1110, {FpAlu_8U_23U_or_877_cse , (FpAlu_8U_23U_and_680_nl) , (FpAlu_8U_23U_and_681_nl)
      , (FpAlu_8U_23U_and_682_nl)});
  assign FpAlu_8U_23U_not_128_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_58_nl = MUX_v_4_2_2(4'b0000, (FpAlu_8U_23U_mux1h_1007_nl),
      (FpAlu_8U_23U_not_128_nl));
  assign and_4044_nl = nor_7_ssc & (~ or_dcpl_1117);
  assign or_5175_nl = io_read_cfg_alu_bypass_rsc_svs_7 | FpAlu_8U_23U_or_859_itm_4
      | FpAlu_8U_23U_equal_tmp_237 | (cfg_precision!=2'b10) | FpAlu_8U_23U_nor_dfs_79
      | reg_FpAlu_8U_23U_or_794_cse;
  assign nand_442_nl = ~(((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_15_lpi_1_dfm_10)
      & (cfg_precision[1]) & (~(FpAlu_8U_23U_or_859_itm_4 | FpAlu_8U_23U_equal_tmp_237
      | (cfg_precision[0]))));
  assign mux_1611_nl = MUX_s_1_2_2((nand_442_nl), (or_5175_nl), or_dcpl_1117);
  assign FpAlu_8U_23U_and_685_nl = (~(FpAdd_8U_23U_and_47_tmp | FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0))
      & alu_loop_op_if_alu_loop_op_if_nor_15_cse & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_686_nl = FpAdd_8U_23U_and_111_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_and_687_nl = FpAdd_8U_23U_and_143_ssc & FpAlu_8U_23U_nor_dfs_79;
  assign FpAlu_8U_23U_mux1h_1005_nl = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_11,
      FpAdd_8U_23U_o_expo_lpi_1_dfm_2_3_0, (FpAdd_8U_23U_o_expo_sva_4[3:0]), 4'b1110,
      {FpAlu_8U_23U_or_878_cse , (FpAlu_8U_23U_and_685_nl) , (FpAlu_8U_23U_and_686_nl)
      , (FpAlu_8U_23U_and_687_nl)});
  assign FpAlu_8U_23U_not_129_nl = ~ FpAlu_8U_23U_equal_tmp_237;
  assign FpAlu_8U_23U_and_62_nl = MUX_v_4_2_2(4'b0000, (FpAlu_8U_23U_mux1h_1005_nl),
      (FpAlu_8U_23U_not_129_nl));
  assign and_4038_nl = nor_7_ssc & (~ or_dcpl_1122);
  assign or_5181_nl = io_read_cfg_alu_bypass_rsc_svs_7 | FpAlu_8U_23U_or_861_itm_4
      | FpAlu_8U_23U_equal_tmp_237 | (cfg_precision!=2'b10) | FpAlu_8U_23U_nor_dfs_79
      | reg_FpAlu_8U_23U_or_797_cse;
  assign nand_443_nl = ~(((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_lpi_1_dfm_10)
      & (cfg_precision[1]) & (~(FpAlu_8U_23U_or_861_itm_4 | FpAlu_8U_23U_equal_tmp_237
      | (cfg_precision[0]))));
  assign mux_1614_nl = MUX_s_1_2_2((nand_443_nl), (or_5181_nl), or_dcpl_1122);
  assign and_492_nl = (or_22_cse | FpCmp_8U_23U_true_if_acc_16_itm_8_1) & and_89_tmp;
  assign and_509_nl = (or_22_cse | FpCmp_8U_23U_true_if_acc_18_itm_8_1) & and_89_tmp;
  assign and_522_nl = (or_22_cse | FpCmp_8U_23U_true_if_acc_20_itm_8_1) & and_89_tmp;
  assign and_535_nl = (or_22_cse | FpCmp_8U_23U_true_if_acc_22_itm_8_1) & and_89_tmp;
  assign and_548_nl = (or_22_cse | FpCmp_8U_23U_true_if_acc_24_itm_8_1) & and_89_tmp;
  assign and_561_nl = (or_22_cse | FpCmp_8U_23U_true_if_acc_26_itm_8_1) & and_89_tmp;
  assign and_574_nl = (or_22_cse | FpCmp_8U_23U_true_if_acc_28_itm_8_1) & and_89_tmp;
  assign and_587_nl = (or_22_cse | FpCmp_8U_23U_true_if_acc_30_itm_8_1) & and_89_tmp;
  assign and_600_nl = (or_22_cse | FpCmp_8U_23U_true_if_acc_32_itm_8_1) & and_89_tmp;
  assign and_613_nl = (or_22_cse | FpCmp_8U_23U_true_if_acc_34_itm_8_1) & and_89_tmp;
  assign and_626_nl = (or_22_cse | FpCmp_8U_23U_true_if_acc_36_itm_8_1) & and_89_tmp;
  assign and_639_nl = (or_22_cse | FpCmp_8U_23U_true_if_acc_38_itm_8_1) & and_89_tmp;
  assign and_652_nl = (or_22_cse | FpCmp_8U_23U_true_if_acc_40_itm_8_1) & and_89_tmp;
  assign and_665_nl = (or_22_cse | FpCmp_8U_23U_true_if_acc_42_itm_8_1) & and_89_tmp;
  assign and_678_nl = (or_22_cse | FpCmp_8U_23U_true_if_acc_44_itm_8_1) & and_89_tmp;
  assign and_691_nl = (or_22_cse | FpCmp_8U_23U_true_if_acc_46_itm_8_1) & and_89_tmp;
  assign or_35_nl = (~((~ FpCmp_8U_23U_true_if_acc_18_itm_8_1) | (cfg_precision!=2'b10)))
      | io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign mux_17_nl = MUX_s_1_2_2((or_35_nl), or_tmp_24, reg_alu_loop_op_2_FpAdd_8U_23U_is_a_greater_slc_8_1_svs_cse);
  assign nor_2052_nl = ~((cfg_alu_algo_1_sva_st_92!=2'b10) | (mux_17_nl));
  assign nor_2053_nl = ~((reg_cfg_alu_algo_1_sva_st_93_cse!=2'b10) | alu_loop_op_2_FpAdd_8U_23U_is_a_greater_slc_8_1_svs_st_2
      | (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (~ main_stage_v_2));
  assign mux_18_nl = MUX_s_1_2_2((nor_2053_nl), (nor_2052_nl), and_89_tmp);
  assign mux_170_nl = MUX_s_1_2_2(mux_157_cse, or_338_cse, cfg_alu_algo_1_sva_st_204[0]);
  assign or_359_nl = (cfg_alu_algo_1_sva_st_204[0]) | (~ reg_chn_alu_out_rsci_ld_core_psct_cse)
      | chn_alu_out_rsci_bawt | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign mux_171_nl = MUX_s_1_2_2((or_359_nl), (mux_170_nl), reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign or_361_nl = (reg_cfg_alu_algo_1_sva_st_93_cse!=2'b10) | or_tmp_327;
  assign mux_172_nl = MUX_s_1_2_2((or_361_nl), (mux_171_nl), cfg_alu_algo_1_sva_st_204[1]);
  assign nor_1745_nl = ~((~((~((~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_8) | IsNaN_8U_23U_land_1_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_831_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign mux_383_nl = MUX_s_1_2_2(nor_1748_cse, (nor_1745_nl), nor_326_cse);
  assign mux_384_nl = MUX_s_1_2_2(nor_1748_cse, (mux_383_nl), FpAlu_8U_23U_nor_dfs_48);
  assign nor_1751_nl = ~((~(IsNaN_8U_23U_land_1_lpi_1_dfm_10 | (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_9)
      | (~ FpAlu_8U_23U_nor_dfs_79))) | FpAlu_8U_23U_or_831_itm_4);
  assign nor_1752_nl = ~(FpAlu_8U_23U_nor_dfs_79 | FpAlu_8U_23U_or_831_itm_4);
  assign mux_385_nl = MUX_s_1_2_2((nor_1752_nl), (nor_1751_nl), nor_327_cse);
  assign nor_1750_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      FpAlu_8U_23U_equal_tmp_237 | (mux_385_nl));
  assign mux_386_nl = MUX_s_1_2_2((nor_1750_nl), (mux_384_nl), or_cse_2);
  assign nor_1739_nl = ~((~ FpAdd_8U_23U_mux_2_tmp_49) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1740_nl = ~((~ alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm)
      | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign mux_389_nl = MUX_s_1_2_2((nor_1740_nl), (nor_1739_nl), nor_333_cse);
  assign nor_1741_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2)));
  assign mux_390_nl = MUX_s_1_2_2((nor_1741_nl), (mux_389_nl), or_cse_2);
  assign nor_1731_nl = ~((((~ FpAlu_8U_23U_nor_dfs_48) | IsNaN_8U_23U_land_1_lpi_1_dfm_9
      | IsNaN_8U_23U_3_land_1_lpi_1_dfm_7) & FpAlu_8U_23U_equal_tmp_146) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1732_nl = ~((((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_1_lpi_1_dfm_10
      | IsNaN_8U_23U_land_1_lpi_1_dfm_st_5) & FpAlu_8U_23U_equal_tmp_237) | (~ main_stage_v_4)
      | io_read_cfg_alu_bypass_rsc_svs_7 | (cfg_alu_algo_1_sva_st_205!=2'b10));
  assign mux_397_nl = MUX_s_1_2_2((nor_1732_nl), (nor_1731_nl), or_cse_2);
  assign nor_1726_nl = ~((~((~((cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48)
      | (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_8) | IsNaN_8U_23U_land_1_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_831_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1729_nl = ~((~((~((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_1_lpi_1_dfm_10
      | (cfg_alu_algo_1_sva_st_205!=2'b10) | (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_831_itm_4)) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign mux_404_nl = MUX_s_1_2_2((nor_1729_nl), (nor_1726_nl), or_cse_2);
  assign nor_1717_nl = ~((~((~((~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_8) | IsNaN_8U_23U_land_2_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_833_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign mux_405_nl = MUX_s_1_2_2(nor_1720_cse, (nor_1717_nl), nor_326_cse);
  assign mux_406_nl = MUX_s_1_2_2(nor_1720_cse, (mux_405_nl), FpAlu_8U_23U_nor_dfs_48);
  assign nor_1722_nl = ~((~((~(IsNaN_8U_23U_land_2_lpi_1_dfm_10 | (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_833_itm_4)) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign mux_407_nl = MUX_s_1_2_2(nor_1724_cse, (nor_1722_nl), nor_327_cse);
  assign mux_408_nl = MUX_s_1_2_2(nor_1724_cse, (mux_407_nl), FpAlu_8U_23U_nor_dfs_79);
  assign mux_409_nl = MUX_s_1_2_2((mux_408_nl), (mux_406_nl), or_cse_2);
  assign nor_1711_nl = ~((~ FpAdd_8U_23U_mux_18_tmp_49) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1712_nl = ~((~ alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm)
      | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign mux_412_nl = MUX_s_1_2_2((nor_1712_nl), (nor_1711_nl), nor_333_cse);
  assign nor_1713_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2)));
  assign mux_413_nl = MUX_s_1_2_2((nor_1713_nl), (mux_412_nl), or_cse_2);
  assign nor_1704_nl = ~((((~ FpAlu_8U_23U_nor_dfs_48) | IsNaN_8U_23U_land_2_lpi_1_dfm_9
      | IsNaN_8U_23U_2_land_2_lpi_1_dfm_8) & FpAlu_8U_23U_equal_tmp_146) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1705_nl = ~((((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_2_lpi_1_dfm_10
      | IsNaN_8U_23U_land_2_lpi_1_dfm_st_5) & FpAlu_8U_23U_equal_tmp_237) | (~ main_stage_v_4)
      | io_read_cfg_alu_bypass_rsc_svs_7 | (cfg_alu_algo_1_sva_st_205!=2'b10));
  assign mux_419_nl = MUX_s_1_2_2((nor_1705_nl), (nor_1704_nl), or_cse_2);
  assign nor_1699_nl = ~((~((~((cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48)
      | (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_8) | IsNaN_8U_23U_land_2_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_833_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1702_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      FpAlu_8U_23U_equal_tmp_237 | (~((~((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_2_lpi_1_dfm_10
      | (cfg_alu_algo_1_sva_st_205!=2'b10) | (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_833_itm_4)));
  assign mux_425_nl = MUX_s_1_2_2((nor_1702_nl), (nor_1699_nl), or_cse_2);
  assign nor_1690_nl = ~((~((~((~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_8) | IsNaN_8U_23U_land_3_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_835_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign mux_426_nl = MUX_s_1_2_2(nor_1693_cse, (nor_1690_nl), nor_326_cse);
  assign mux_427_nl = MUX_s_1_2_2(nor_1693_cse, (mux_426_nl), FpAlu_8U_23U_nor_dfs_48);
  assign nor_1695_nl = ~((~((~(IsNaN_8U_23U_land_3_lpi_1_dfm_10 | (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_835_itm_4)) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign mux_428_nl = MUX_s_1_2_2(nor_1697_cse, (nor_1695_nl), nor_327_cse);
  assign mux_429_nl = MUX_s_1_2_2(nor_1697_cse, (mux_428_nl), FpAlu_8U_23U_nor_dfs_79);
  assign mux_430_nl = MUX_s_1_2_2((mux_429_nl), (mux_427_nl), or_cse_2);
  assign nor_1684_nl = ~((~ FpAdd_8U_23U_mux_34_tmp_49) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1685_nl = ~((~ alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm)
      | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign mux_433_nl = MUX_s_1_2_2((nor_1685_nl), (nor_1684_nl), nor_333_cse);
  assign nor_1686_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2)));
  assign mux_434_nl = MUX_s_1_2_2((nor_1686_nl), (mux_433_nl), or_cse_2);
  assign nor_1677_nl = ~((((~ FpAlu_8U_23U_nor_dfs_48) | IsNaN_8U_23U_land_3_lpi_1_dfm_9
      | IsNaN_8U_23U_3_land_3_lpi_1_dfm_7) & FpAlu_8U_23U_equal_tmp_146) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1678_nl = ~((((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_3_lpi_1_dfm_10
      | IsNaN_8U_23U_land_3_lpi_1_dfm_st_5) & FpAlu_8U_23U_equal_tmp_237) | (~ main_stage_v_4)
      | io_read_cfg_alu_bypass_rsc_svs_7 | (cfg_alu_algo_1_sva_st_205!=2'b10));
  assign mux_440_nl = MUX_s_1_2_2((nor_1678_nl), (nor_1677_nl), or_cse_2);
  assign nor_1672_nl = ~((~((~((cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48)
      | (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_8) | IsNaN_8U_23U_land_3_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_835_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1675_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      FpAlu_8U_23U_equal_tmp_237 | (~((~((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_3_lpi_1_dfm_10
      | (cfg_alu_algo_1_sva_st_205!=2'b10) | (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_835_itm_4)));
  assign mux_446_nl = MUX_s_1_2_2((nor_1675_nl), (nor_1672_nl), or_cse_2);
  assign nor_1663_nl = ~((~((~((~ IsNaN_8U_23U_1_land_4_lpi_1_dfm_8) | IsNaN_8U_23U_land_4_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_837_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign mux_447_nl = MUX_s_1_2_2(nor_1666_cse, (nor_1663_nl), nor_326_cse);
  assign mux_448_nl = MUX_s_1_2_2(nor_1666_cse, (mux_447_nl), FpAlu_8U_23U_nor_dfs_48);
  assign nor_1668_nl = ~((~((~(IsNaN_8U_23U_land_4_lpi_1_dfm_10 | (~ IsNaN_8U_23U_1_land_4_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_837_itm_4)) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign mux_449_nl = MUX_s_1_2_2(nor_1670_cse, (nor_1668_nl), nor_327_cse);
  assign mux_450_nl = MUX_s_1_2_2(nor_1670_cse, (mux_449_nl), FpAlu_8U_23U_nor_dfs_79);
  assign mux_451_nl = MUX_s_1_2_2((mux_450_nl), (mux_448_nl), or_cse_2);
  assign nor_1657_nl = ~((~ FpAdd_8U_23U_mux_50_tmp_49) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1658_nl = ~((~ alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm)
      | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign mux_454_nl = MUX_s_1_2_2((nor_1658_nl), (nor_1657_nl), nor_333_cse);
  assign nor_1659_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2)));
  assign mux_455_nl = MUX_s_1_2_2((nor_1659_nl), (mux_454_nl), or_cse_2);
  assign nor_1650_nl = ~((((~ FpAlu_8U_23U_nor_dfs_48) | IsNaN_8U_23U_land_4_lpi_1_dfm_9
      | IsNaN_8U_23U_2_land_4_lpi_1_dfm_8) & FpAlu_8U_23U_equal_tmp_146) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1651_nl = ~((((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_4_lpi_1_dfm_10
      | IsNaN_8U_23U_land_4_lpi_1_dfm_st_5) & FpAlu_8U_23U_equal_tmp_237) | (~ main_stage_v_4)
      | io_read_cfg_alu_bypass_rsc_svs_7 | (cfg_alu_algo_1_sva_st_205!=2'b10));
  assign mux_461_nl = MUX_s_1_2_2((nor_1651_nl), (nor_1650_nl), or_cse_2);
  assign nor_1645_nl = ~((~((~((cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48)
      | (~ IsNaN_8U_23U_1_land_4_lpi_1_dfm_8) | IsNaN_8U_23U_land_4_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_837_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1648_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      FpAlu_8U_23U_equal_tmp_237 | (~((~((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_4_lpi_1_dfm_10
      | (cfg_alu_algo_1_sva_st_205!=2'b10) | (~ IsNaN_8U_23U_1_land_4_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_837_itm_4)));
  assign mux_467_nl = MUX_s_1_2_2((nor_1648_nl), (nor_1645_nl), or_cse_2);
  assign nor_1636_nl = ~((~((~((~ IsNaN_8U_23U_1_land_5_lpi_1_dfm_8) | IsNaN_8U_23U_land_5_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_839_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign mux_468_nl = MUX_s_1_2_2(nor_1639_cse, (nor_1636_nl), nor_326_cse);
  assign mux_469_nl = MUX_s_1_2_2(nor_1639_cse, (mux_468_nl), FpAlu_8U_23U_nor_dfs_48);
  assign nor_1641_nl = ~((~((~(IsNaN_8U_23U_land_5_lpi_1_dfm_10 | (~ IsNaN_8U_23U_1_land_5_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_839_itm_4)) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign mux_470_nl = MUX_s_1_2_2(nor_1643_cse, (nor_1641_nl), nor_327_cse);
  assign mux_471_nl = MUX_s_1_2_2(nor_1643_cse, (mux_470_nl), FpAlu_8U_23U_nor_dfs_79);
  assign mux_472_nl = MUX_s_1_2_2((mux_471_nl), (mux_469_nl), or_cse_2);
  assign nor_1630_nl = ~((~ FpAdd_8U_23U_mux_66_tmp_49) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1631_nl = ~((~ alu_loop_op_5_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm)
      | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign mux_475_nl = MUX_s_1_2_2((nor_1631_nl), (nor_1630_nl), nor_333_cse);
  assign nor_1632_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & alu_loop_op_5_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2)));
  assign mux_476_nl = MUX_s_1_2_2((nor_1632_nl), (mux_475_nl), or_cse_2);
  assign nor_1623_nl = ~((((~ FpAlu_8U_23U_nor_dfs_48) | IsNaN_8U_23U_land_5_lpi_1_dfm_9
      | IsNaN_8U_23U_2_land_5_lpi_1_dfm_8) & FpAlu_8U_23U_equal_tmp_146) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1624_nl = ~((((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_5_lpi_1_dfm_10
      | IsNaN_8U_23U_land_5_lpi_1_dfm_st_5) & FpAlu_8U_23U_equal_tmp_237) | (~ main_stage_v_4)
      | io_read_cfg_alu_bypass_rsc_svs_7 | (cfg_alu_algo_1_sva_st_205!=2'b10));
  assign mux_482_nl = MUX_s_1_2_2((nor_1624_nl), (nor_1623_nl), or_cse_2);
  assign nor_1618_nl = ~((~((~((cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48)
      | (~ IsNaN_8U_23U_1_land_5_lpi_1_dfm_8) | IsNaN_8U_23U_land_5_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_839_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1621_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      FpAlu_8U_23U_equal_tmp_237 | (~((~((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_5_lpi_1_dfm_10
      | (cfg_alu_algo_1_sva_st_205!=2'b10) | (~ IsNaN_8U_23U_1_land_5_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_839_itm_4)));
  assign mux_488_nl = MUX_s_1_2_2((nor_1621_nl), (nor_1618_nl), or_cse_2);
  assign nor_1609_nl = ~((~((~((~ IsNaN_8U_23U_1_land_6_lpi_1_dfm_8) | IsNaN_8U_23U_land_6_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_841_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign mux_489_nl = MUX_s_1_2_2(nor_1612_cse, (nor_1609_nl), nor_326_cse);
  assign mux_490_nl = MUX_s_1_2_2(nor_1612_cse, (mux_489_nl), FpAlu_8U_23U_nor_dfs_48);
  assign nor_1614_nl = ~((~((~(IsNaN_8U_23U_land_6_lpi_1_dfm_10 | (~ IsNaN_8U_23U_1_land_6_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_841_itm_4)) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign mux_491_nl = MUX_s_1_2_2(nor_1616_cse, (nor_1614_nl), nor_327_cse);
  assign mux_492_nl = MUX_s_1_2_2(nor_1616_cse, (mux_491_nl), FpAlu_8U_23U_nor_dfs_79);
  assign mux_493_nl = MUX_s_1_2_2((mux_492_nl), (mux_490_nl), or_cse_2);
  assign nor_1603_nl = ~((~ FpAdd_8U_23U_mux_82_tmp_49) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1604_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204[0]) | (~((cfg_alu_algo_1_sva_st_204[1]) & alu_loop_op_6_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm)));
  assign mux_496_nl = MUX_s_1_2_2((nor_1604_nl), (nor_1603_nl), nor_333_cse);
  assign nor_1605_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & alu_loop_op_6_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2)));
  assign mux_497_nl = MUX_s_1_2_2((nor_1605_nl), (mux_496_nl), or_cse_2);
  assign nor_1596_nl = ~((((~ FpAlu_8U_23U_nor_dfs_48) | IsNaN_8U_23U_land_6_lpi_1_dfm_9
      | IsNaN_8U_23U_2_land_6_lpi_1_dfm_8) & FpAlu_8U_23U_equal_tmp_146) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1597_nl = ~((((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_6_lpi_1_dfm_10
      | IsNaN_8U_23U_land_6_lpi_1_dfm_st_5) & FpAlu_8U_23U_equal_tmp_237) | (~ main_stage_v_4)
      | io_read_cfg_alu_bypass_rsc_svs_7 | (cfg_alu_algo_1_sva_st_205!=2'b10));
  assign mux_503_nl = MUX_s_1_2_2((nor_1597_nl), (nor_1596_nl), or_cse_2);
  assign nor_1591_nl = ~((~((~((cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48)
      | (~ IsNaN_8U_23U_1_land_6_lpi_1_dfm_8) | IsNaN_8U_23U_land_6_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_841_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1594_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      FpAlu_8U_23U_equal_tmp_237 | (~((~((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_6_lpi_1_dfm_10
      | (cfg_alu_algo_1_sva_st_205!=2'b10) | (~ IsNaN_8U_23U_1_land_6_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_841_itm_4)));
  assign mux_509_nl = MUX_s_1_2_2((nor_1594_nl), (nor_1591_nl), or_cse_2);
  assign nor_1582_nl = ~((~((~((~ IsNaN_8U_23U_1_land_7_lpi_1_dfm_8) | IsNaN_8U_23U_land_7_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_843_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign mux_510_nl = MUX_s_1_2_2(nor_1585_cse, (nor_1582_nl), nor_326_cse);
  assign mux_511_nl = MUX_s_1_2_2(nor_1585_cse, (mux_510_nl), FpAlu_8U_23U_nor_dfs_48);
  assign nor_1587_nl = ~((~((~(IsNaN_8U_23U_land_7_lpi_1_dfm_10 | (~ IsNaN_8U_23U_1_land_7_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_843_itm_4)) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign mux_512_nl = MUX_s_1_2_2(nor_1589_cse, (nor_1587_nl), nor_327_cse);
  assign mux_513_nl = MUX_s_1_2_2(nor_1589_cse, (mux_512_nl), FpAlu_8U_23U_nor_dfs_79);
  assign mux_514_nl = MUX_s_1_2_2((mux_513_nl), (mux_511_nl), or_cse_2);
  assign nor_1577_nl = ~((~ FpAdd_8U_23U_mux_98_tmp_49) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1578_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204[0]) | (~((cfg_alu_algo_1_sva_st_204[1]) & alu_loop_op_7_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm)));
  assign mux_517_nl = MUX_s_1_2_2((nor_1578_nl), (nor_1577_nl), nor_333_cse);
  assign nor_1579_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & alu_loop_op_7_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2)));
  assign mux_518_nl = MUX_s_1_2_2((nor_1579_nl), (mux_517_nl), or_cse_2);
  assign nor_1570_nl = ~((((~ FpAlu_8U_23U_nor_dfs_48) | IsNaN_8U_23U_land_7_lpi_1_dfm_9
      | IsNaN_8U_23U_3_land_7_lpi_1_dfm_7) & FpAlu_8U_23U_equal_tmp_146) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1571_nl = ~((((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_7_lpi_1_dfm_10
      | IsNaN_8U_23U_land_7_lpi_1_dfm_st_5) & FpAlu_8U_23U_equal_tmp_237) | (~ main_stage_v_4)
      | io_read_cfg_alu_bypass_rsc_svs_7 | (cfg_alu_algo_1_sva_st_205!=2'b10));
  assign mux_524_nl = MUX_s_1_2_2((nor_1571_nl), (nor_1570_nl), or_cse_2);
  assign nor_1565_nl = ~((~((~((cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48)
      | (~ IsNaN_8U_23U_1_land_7_lpi_1_dfm_8) | IsNaN_8U_23U_land_7_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_843_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1568_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      FpAlu_8U_23U_equal_tmp_237 | (~((~((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_7_lpi_1_dfm_10
      | (cfg_alu_algo_1_sva_st_205!=2'b10) | (~ IsNaN_8U_23U_1_land_7_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_843_itm_4)));
  assign mux_530_nl = MUX_s_1_2_2((nor_1568_nl), (nor_1565_nl), or_cse_2);
  assign nor_1556_nl = ~((~((~((~ IsNaN_8U_23U_1_land_8_lpi_1_dfm_8) | IsNaN_8U_23U_land_8_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_845_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign mux_531_nl = MUX_s_1_2_2(nor_1559_cse, (nor_1556_nl), nor_326_cse);
  assign mux_532_nl = MUX_s_1_2_2(nor_1559_cse, (mux_531_nl), FpAlu_8U_23U_nor_dfs_48);
  assign nor_1561_nl = ~((~((~(IsNaN_8U_23U_land_8_lpi_1_dfm_10 | (~ IsNaN_8U_23U_1_land_8_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_845_itm_4)) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign mux_533_nl = MUX_s_1_2_2(nor_1563_cse, (nor_1561_nl), nor_327_cse);
  assign mux_534_nl = MUX_s_1_2_2(nor_1563_cse, (mux_533_nl), FpAlu_8U_23U_nor_dfs_79);
  assign mux_535_nl = MUX_s_1_2_2((mux_534_nl), (mux_532_nl), or_cse_2);
  assign nor_1551_nl = ~((~ FpAdd_8U_23U_mux_114_tmp_49) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1552_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204[0]) | (~((cfg_alu_algo_1_sva_st_204[1]) & alu_loop_op_8_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm)));
  assign mux_538_nl = MUX_s_1_2_2((nor_1552_nl), (nor_1551_nl), nor_333_cse);
  assign nor_1553_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & alu_loop_op_8_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2)));
  assign mux_539_nl = MUX_s_1_2_2((nor_1553_nl), (mux_538_nl), or_cse_2);
  assign nor_1544_nl = ~((((~ FpAlu_8U_23U_nor_dfs_48) | IsNaN_8U_23U_land_8_lpi_1_dfm_9
      | IsNaN_8U_23U_3_land_8_lpi_1_dfm_7) & FpAlu_8U_23U_equal_tmp_146) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1545_nl = ~((((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_8_lpi_1_dfm_10
      | IsNaN_8U_23U_land_8_lpi_1_dfm_st_5) & FpAlu_8U_23U_equal_tmp_237) | (~ main_stage_v_4)
      | io_read_cfg_alu_bypass_rsc_svs_7 | (cfg_alu_algo_1_sva_st_205!=2'b10));
  assign mux_545_nl = MUX_s_1_2_2((nor_1545_nl), (nor_1544_nl), or_cse_2);
  assign nor_1539_nl = ~((~((~((cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48)
      | (~ IsNaN_8U_23U_1_land_8_lpi_1_dfm_8) | IsNaN_8U_23U_land_8_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_845_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1542_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      FpAlu_8U_23U_equal_tmp_237 | (~((~((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_8_lpi_1_dfm_10
      | (cfg_alu_algo_1_sva_st_205!=2'b10) | (~ IsNaN_8U_23U_1_land_8_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_845_itm_4)));
  assign mux_551_nl = MUX_s_1_2_2((nor_1542_nl), (nor_1539_nl), or_cse_2);
  assign nor_1530_nl = ~((~((~((~ IsNaN_8U_23U_1_land_9_lpi_1_dfm_8) | IsNaN_8U_23U_land_9_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_847_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign mux_552_nl = MUX_s_1_2_2(nor_1533_cse, (nor_1530_nl), nor_326_cse);
  assign mux_553_nl = MUX_s_1_2_2(nor_1533_cse, (mux_552_nl), FpAlu_8U_23U_nor_dfs_48);
  assign nor_1535_nl = ~((~((~(IsNaN_8U_23U_land_9_lpi_1_dfm_10 | (~ IsNaN_8U_23U_1_land_9_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_847_itm_4)) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign mux_554_nl = MUX_s_1_2_2(nor_1537_cse, (nor_1535_nl), nor_327_cse);
  assign mux_555_nl = MUX_s_1_2_2(nor_1537_cse, (mux_554_nl), FpAlu_8U_23U_nor_dfs_79);
  assign mux_556_nl = MUX_s_1_2_2((mux_555_nl), (mux_553_nl), or_cse_2);
  assign nor_1525_nl = ~((~ FpAdd_8U_23U_mux_130_tmp_49) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1526_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204[0]) | (~((cfg_alu_algo_1_sva_st_204[1]) & alu_loop_op_9_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm)));
  assign mux_559_nl = MUX_s_1_2_2((nor_1526_nl), (nor_1525_nl), nor_333_cse);
  assign nor_1527_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & alu_loop_op_9_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2)));
  assign mux_560_nl = MUX_s_1_2_2((nor_1527_nl), (mux_559_nl), or_cse_2);
  assign nor_1518_nl = ~((((~ FpAlu_8U_23U_nor_dfs_48) | IsNaN_8U_23U_land_9_lpi_1_dfm_9
      | IsNaN_8U_23U_2_land_9_lpi_1_dfm_8) & FpAlu_8U_23U_equal_tmp_146) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1519_nl = ~((((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_9_lpi_1_dfm_10
      | IsNaN_8U_23U_land_9_lpi_1_dfm_st_5) & FpAlu_8U_23U_equal_tmp_237) | (~ main_stage_v_4)
      | io_read_cfg_alu_bypass_rsc_svs_7 | (cfg_alu_algo_1_sva_st_205!=2'b10));
  assign mux_566_nl = MUX_s_1_2_2((nor_1519_nl), (nor_1518_nl), or_cse_2);
  assign nor_1513_nl = ~((~((~((cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48)
      | (~ IsNaN_8U_23U_1_land_9_lpi_1_dfm_8) | IsNaN_8U_23U_land_9_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_847_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1516_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      FpAlu_8U_23U_equal_tmp_237 | (~((~((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_9_lpi_1_dfm_10
      | (cfg_alu_algo_1_sva_st_205!=2'b10) | (~ IsNaN_8U_23U_1_land_9_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_847_itm_4)));
  assign mux_572_nl = MUX_s_1_2_2((nor_1516_nl), (nor_1513_nl), or_cse_2);
  assign nor_1504_nl = ~((~((~((~ IsNaN_8U_23U_1_land_10_lpi_1_dfm_8) | IsNaN_8U_23U_land_10_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_849_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign mux_573_nl = MUX_s_1_2_2(nor_1507_cse, (nor_1504_nl), nor_326_cse);
  assign mux_574_nl = MUX_s_1_2_2(nor_1507_cse, (mux_573_nl), FpAlu_8U_23U_nor_dfs_48);
  assign nor_1509_nl = ~((~((~(IsNaN_8U_23U_land_10_lpi_1_dfm_10 | (~ IsNaN_8U_23U_1_land_10_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_849_itm_4)) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign mux_575_nl = MUX_s_1_2_2(nor_1511_cse, (nor_1509_nl), nor_327_cse);
  assign mux_576_nl = MUX_s_1_2_2(nor_1511_cse, (mux_575_nl), FpAlu_8U_23U_nor_dfs_79);
  assign mux_577_nl = MUX_s_1_2_2((mux_576_nl), (mux_574_nl), or_cse_2);
  assign nor_1499_nl = ~((~ FpAdd_8U_23U_mux_146_tmp_49) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1500_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204[0]) | (~((cfg_alu_algo_1_sva_st_204[1]) & alu_loop_op_10_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm)));
  assign mux_580_nl = MUX_s_1_2_2((nor_1500_nl), (nor_1499_nl), nor_333_cse);
  assign nor_1501_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & alu_loop_op_10_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2)));
  assign mux_581_nl = MUX_s_1_2_2((nor_1501_nl), (mux_580_nl), or_cse_2);
  assign nor_1492_nl = ~((((~ FpAlu_8U_23U_nor_dfs_48) | IsNaN_8U_23U_land_10_lpi_1_dfm_9
      | IsNaN_8U_23U_2_land_10_lpi_1_dfm_8) & FpAlu_8U_23U_equal_tmp_146) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1493_nl = ~((((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_10_lpi_1_dfm_10
      | IsNaN_8U_23U_land_10_lpi_1_dfm_st_5) & FpAlu_8U_23U_equal_tmp_237) | (~ main_stage_v_4)
      | io_read_cfg_alu_bypass_rsc_svs_7 | (cfg_alu_algo_1_sva_st_205!=2'b10));
  assign mux_587_nl = MUX_s_1_2_2((nor_1493_nl), (nor_1492_nl), or_cse_2);
  assign nor_1487_nl = ~((~((~((cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48)
      | (~ IsNaN_8U_23U_1_land_10_lpi_1_dfm_8) | IsNaN_8U_23U_land_10_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_849_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1490_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      FpAlu_8U_23U_equal_tmp_237 | (~((~((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_10_lpi_1_dfm_10
      | (cfg_alu_algo_1_sva_st_205!=2'b10) | (~ IsNaN_8U_23U_1_land_10_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_849_itm_4)));
  assign mux_593_nl = MUX_s_1_2_2((nor_1490_nl), (nor_1487_nl), or_cse_2);
  assign nor_1478_nl = ~((~((~((~ IsNaN_8U_23U_1_land_11_lpi_1_dfm_8) | IsNaN_8U_23U_land_11_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_851_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign mux_594_nl = MUX_s_1_2_2(nor_1481_cse, (nor_1478_nl), nor_326_cse);
  assign mux_595_nl = MUX_s_1_2_2(nor_1481_cse, (mux_594_nl), FpAlu_8U_23U_nor_dfs_48);
  assign nor_1483_nl = ~((~((~(IsNaN_8U_23U_land_11_lpi_1_dfm_10 | (~ IsNaN_8U_23U_1_land_11_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_851_itm_4)) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign mux_596_nl = MUX_s_1_2_2(nor_1485_cse, (nor_1483_nl), nor_327_cse);
  assign mux_597_nl = MUX_s_1_2_2(nor_1485_cse, (mux_596_nl), FpAlu_8U_23U_nor_dfs_79);
  assign mux_598_nl = MUX_s_1_2_2((mux_597_nl), (mux_595_nl), or_cse_2);
  assign nor_1473_nl = ~((~ FpAdd_8U_23U_mux_162_tmp_49) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1474_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204[0]) | (~((cfg_alu_algo_1_sva_st_204[1]) & alu_loop_op_11_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm)));
  assign mux_601_nl = MUX_s_1_2_2((nor_1474_nl), (nor_1473_nl), nor_333_cse);
  assign nor_1475_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & alu_loop_op_11_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2)));
  assign mux_602_nl = MUX_s_1_2_2((nor_1475_nl), (mux_601_nl), or_cse_2);
  assign nor_1466_nl = ~((((~ FpAlu_8U_23U_nor_dfs_48) | IsNaN_8U_23U_land_11_lpi_1_dfm_9
      | IsNaN_8U_23U_2_land_11_lpi_1_dfm_8) & FpAlu_8U_23U_equal_tmp_146) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1467_nl = ~((((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_11_lpi_1_dfm_10
      | IsNaN_8U_23U_land_11_lpi_1_dfm_st_5) & FpAlu_8U_23U_equal_tmp_237) | (~ main_stage_v_4)
      | io_read_cfg_alu_bypass_rsc_svs_7 | (cfg_alu_algo_1_sva_st_205!=2'b10));
  assign mux_608_nl = MUX_s_1_2_2((nor_1467_nl), (nor_1466_nl), or_cse_2);
  assign nor_1461_nl = ~((~((~((cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48)
      | (~ IsNaN_8U_23U_1_land_11_lpi_1_dfm_8) | IsNaN_8U_23U_land_11_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_851_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1464_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      FpAlu_8U_23U_equal_tmp_237 | (~((~((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_11_lpi_1_dfm_10
      | (cfg_alu_algo_1_sva_st_205!=2'b10) | (~ IsNaN_8U_23U_1_land_11_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_851_itm_4)));
  assign mux_614_nl = MUX_s_1_2_2((nor_1464_nl), (nor_1461_nl), or_cse_2);
  assign nor_1452_nl = ~((~((~((~ IsNaN_8U_23U_1_land_12_lpi_1_dfm_8) | IsNaN_8U_23U_land_12_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_853_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign mux_615_nl = MUX_s_1_2_2(nor_1455_cse, (nor_1452_nl), nor_326_cse);
  assign mux_616_nl = MUX_s_1_2_2(nor_1455_cse, (mux_615_nl), FpAlu_8U_23U_nor_dfs_48);
  assign nor_1457_nl = ~((~((~(IsNaN_8U_23U_land_12_lpi_1_dfm_10 | (~ IsNaN_8U_23U_1_land_12_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_853_itm_4)) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign mux_617_nl = MUX_s_1_2_2(nor_1459_cse, (nor_1457_nl), nor_327_cse);
  assign mux_618_nl = MUX_s_1_2_2(nor_1459_cse, (mux_617_nl), FpAlu_8U_23U_nor_dfs_79);
  assign mux_619_nl = MUX_s_1_2_2((mux_618_nl), (mux_616_nl), or_cse_2);
  assign nor_1447_nl = ~((~ FpAdd_8U_23U_mux_178_tmp_49) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1448_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204[0]) | (~((cfg_alu_algo_1_sva_st_204[1]) & alu_loop_op_12_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm)));
  assign mux_622_nl = MUX_s_1_2_2((nor_1448_nl), (nor_1447_nl), nor_333_cse);
  assign nor_1449_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & alu_loop_op_12_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2)));
  assign mux_623_nl = MUX_s_1_2_2((nor_1449_nl), (mux_622_nl), or_cse_2);
  assign nor_1440_nl = ~((((~ FpAlu_8U_23U_nor_dfs_48) | IsNaN_8U_23U_land_12_lpi_1_dfm_9
      | IsNaN_8U_23U_2_land_12_lpi_1_dfm_8) & FpAlu_8U_23U_equal_tmp_146) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1441_nl = ~((((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_12_lpi_1_dfm_10
      | IsNaN_8U_23U_land_12_lpi_1_dfm_st_5) & FpAlu_8U_23U_equal_tmp_237) | (~ main_stage_v_4)
      | io_read_cfg_alu_bypass_rsc_svs_7 | (cfg_alu_algo_1_sva_st_205!=2'b10));
  assign mux_629_nl = MUX_s_1_2_2((nor_1441_nl), (nor_1440_nl), or_cse_2);
  assign nor_1435_nl = ~((~((~((cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48)
      | (~ IsNaN_8U_23U_1_land_12_lpi_1_dfm_8) | IsNaN_8U_23U_land_12_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_853_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1438_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      FpAlu_8U_23U_equal_tmp_237 | (~((~((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_12_lpi_1_dfm_10
      | (cfg_alu_algo_1_sva_st_205!=2'b10) | (~ IsNaN_8U_23U_1_land_12_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_853_itm_4)));
  assign mux_635_nl = MUX_s_1_2_2((nor_1438_nl), (nor_1435_nl), or_cse_2);
  assign nor_1426_nl = ~((~((~((~ IsNaN_8U_23U_1_land_13_lpi_1_dfm_8) | IsNaN_8U_23U_land_13_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_855_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign mux_636_nl = MUX_s_1_2_2(nor_1429_cse, (nor_1426_nl), nor_326_cse);
  assign mux_637_nl = MUX_s_1_2_2(nor_1429_cse, (mux_636_nl), FpAlu_8U_23U_nor_dfs_48);
  assign nor_1431_nl = ~((~((~(IsNaN_8U_23U_land_13_lpi_1_dfm_10 | (~ IsNaN_8U_23U_1_land_13_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_855_itm_4)) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign mux_638_nl = MUX_s_1_2_2(nor_1433_cse, (nor_1431_nl), nor_327_cse);
  assign mux_639_nl = MUX_s_1_2_2(nor_1433_cse, (mux_638_nl), FpAlu_8U_23U_nor_dfs_79);
  assign mux_640_nl = MUX_s_1_2_2((mux_639_nl), (mux_637_nl), or_cse_2);
  assign nor_1421_nl = ~((~ FpAdd_8U_23U_mux_194_tmp_49) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1422_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204[0]) | (~((cfg_alu_algo_1_sva_st_204[1]) & alu_loop_op_13_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm)));
  assign mux_643_nl = MUX_s_1_2_2((nor_1422_nl), (nor_1421_nl), nor_333_cse);
  assign nor_1423_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & alu_loop_op_13_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2)));
  assign mux_644_nl = MUX_s_1_2_2((nor_1423_nl), (mux_643_nl), or_cse_2);
  assign nor_1414_nl = ~((((~ FpAlu_8U_23U_nor_dfs_48) | IsNaN_8U_23U_land_13_lpi_1_dfm_9
      | IsNaN_8U_23U_2_land_13_lpi_1_dfm_8) & FpAlu_8U_23U_equal_tmp_146) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1415_nl = ~((((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_13_lpi_1_dfm_10
      | IsNaN_8U_23U_land_13_lpi_1_dfm_st_5) & FpAlu_8U_23U_equal_tmp_237) | (~ main_stage_v_4)
      | io_read_cfg_alu_bypass_rsc_svs_7 | (cfg_alu_algo_1_sva_st_205!=2'b10));
  assign mux_650_nl = MUX_s_1_2_2((nor_1415_nl), (nor_1414_nl), or_cse_2);
  assign nor_1409_nl = ~((~((~((cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48)
      | (~ IsNaN_8U_23U_1_land_13_lpi_1_dfm_8) | IsNaN_8U_23U_land_13_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_855_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1412_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      FpAlu_8U_23U_equal_tmp_237 | (~((~((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_13_lpi_1_dfm_10
      | (cfg_alu_algo_1_sva_st_205!=2'b10) | (~ IsNaN_8U_23U_1_land_13_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_855_itm_4)));
  assign mux_656_nl = MUX_s_1_2_2((nor_1412_nl), (nor_1409_nl), or_cse_2);
  assign nor_1400_nl = ~((~((~((~ IsNaN_8U_23U_1_land_14_lpi_1_dfm_8) | IsNaN_8U_23U_land_14_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_857_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign mux_657_nl = MUX_s_1_2_2(nor_1403_cse, (nor_1400_nl), nor_326_cse);
  assign mux_658_nl = MUX_s_1_2_2(nor_1403_cse, (mux_657_nl), FpAlu_8U_23U_nor_dfs_48);
  assign nor_1405_nl = ~((~((~(IsNaN_8U_23U_land_14_lpi_1_dfm_10 | (~ IsNaN_8U_23U_1_land_14_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_857_itm_4)) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign mux_659_nl = MUX_s_1_2_2(nor_1407_cse, (nor_1405_nl), nor_327_cse);
  assign mux_660_nl = MUX_s_1_2_2(nor_1407_cse, (mux_659_nl), FpAlu_8U_23U_nor_dfs_79);
  assign mux_661_nl = MUX_s_1_2_2((mux_660_nl), (mux_658_nl), or_cse_2);
  assign nor_1395_nl = ~((~ FpAdd_8U_23U_mux_210_tmp_49) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1396_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204[0]) | (~((cfg_alu_algo_1_sva_st_204[1]) & alu_loop_op_14_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm)));
  assign mux_664_nl = MUX_s_1_2_2((nor_1396_nl), (nor_1395_nl), nor_333_cse);
  assign nor_1397_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & alu_loop_op_14_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2)));
  assign mux_665_nl = MUX_s_1_2_2((nor_1397_nl), (mux_664_nl), or_cse_2);
  assign nor_1388_nl = ~((((~ FpAlu_8U_23U_nor_dfs_48) | IsNaN_8U_23U_land_14_lpi_1_dfm_9
      | IsNaN_8U_23U_2_land_14_lpi_1_dfm_8) & FpAlu_8U_23U_equal_tmp_146) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1389_nl = ~((((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_14_lpi_1_dfm_10
      | IsNaN_8U_23U_land_14_lpi_1_dfm_st_5) & FpAlu_8U_23U_equal_tmp_237) | (~ main_stage_v_4)
      | io_read_cfg_alu_bypass_rsc_svs_7 | (cfg_alu_algo_1_sva_st_205!=2'b10));
  assign mux_671_nl = MUX_s_1_2_2((nor_1389_nl), (nor_1388_nl), or_cse_2);
  assign nor_1383_nl = ~((~((~((cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48)
      | (~ IsNaN_8U_23U_1_land_14_lpi_1_dfm_8) | IsNaN_8U_23U_land_14_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_857_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1386_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      FpAlu_8U_23U_equal_tmp_237 | (~((~((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_14_lpi_1_dfm_10
      | (cfg_alu_algo_1_sva_st_205!=2'b10) | (~ IsNaN_8U_23U_1_land_14_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_857_itm_4)));
  assign mux_677_nl = MUX_s_1_2_2((nor_1386_nl), (nor_1383_nl), or_cse_2);
  assign nor_1375_nl = ~((~((~((~ IsNaN_8U_23U_1_land_15_lpi_1_dfm_8) | IsNaN_8U_23U_land_15_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_859_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign mux_678_nl = MUX_s_1_2_2(nor_1378_cse, (nor_1375_nl), nor_326_cse);
  assign mux_679_nl = MUX_s_1_2_2(nor_1378_cse, (mux_678_nl), FpAlu_8U_23U_nor_dfs_48);
  assign nor_1381_nl = ~((~(IsNaN_8U_23U_land_15_lpi_1_dfm_10 | (~ IsNaN_8U_23U_1_land_15_lpi_1_dfm_9)
      | (~ FpAlu_8U_23U_nor_dfs_79))) | FpAlu_8U_23U_or_859_itm_4);
  assign nor_1382_nl = ~(FpAlu_8U_23U_nor_dfs_79 | FpAlu_8U_23U_or_859_itm_4);
  assign mux_680_nl = MUX_s_1_2_2((nor_1382_nl), (nor_1381_nl), nor_327_cse);
  assign nor_1380_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      FpAlu_8U_23U_equal_tmp_237 | (mux_680_nl));
  assign mux_681_nl = MUX_s_1_2_2((nor_1380_nl), (mux_679_nl), or_cse_2);
  assign nor_1370_nl = ~((~ FpAdd_8U_23U_mux_226_tmp_49) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1371_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204[0]) | (~((cfg_alu_algo_1_sva_st_204[1]) & alu_loop_op_15_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm)));
  assign mux_684_nl = MUX_s_1_2_2((nor_1371_nl), (nor_1370_nl), nor_333_cse);
  assign nor_1372_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & alu_loop_op_15_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2)));
  assign mux_685_nl = MUX_s_1_2_2((nor_1372_nl), (mux_684_nl), or_cse_2);
  assign nor_1363_nl = ~((((~ FpAlu_8U_23U_nor_dfs_48) | IsNaN_8U_23U_land_15_lpi_1_dfm_9
      | IsNaN_8U_23U_3_land_15_lpi_1_dfm_7) & FpAlu_8U_23U_equal_tmp_146) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1364_nl = ~((((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_15_lpi_1_dfm_10
      | IsNaN_8U_23U_land_15_lpi_1_dfm_st_5) & FpAlu_8U_23U_equal_tmp_237) | (~ main_stage_v_4)
      | io_read_cfg_alu_bypass_rsc_svs_7 | (cfg_alu_algo_1_sva_st_205!=2'b10));
  assign mux_691_nl = MUX_s_1_2_2((nor_1364_nl), (nor_1363_nl), or_cse_2);
  assign nor_1358_nl = ~((~((~((cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48)
      | (~ IsNaN_8U_23U_1_land_15_lpi_1_dfm_8) | IsNaN_8U_23U_land_15_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_859_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1361_nl = ~((~((~((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_15_lpi_1_dfm_10
      | (cfg_alu_algo_1_sva_st_205!=2'b10) | (~ IsNaN_8U_23U_1_land_15_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_859_itm_4)) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign mux_697_nl = MUX_s_1_2_2((nor_1361_nl), (nor_1358_nl), or_cse_2);
  assign nor_1350_nl = ~((~((~((~ IsNaN_8U_23U_1_land_lpi_1_dfm_8) | IsNaN_8U_23U_land_lpi_1_dfm_9))
      | FpAlu_8U_23U_or_861_itm_3)) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | FpAlu_8U_23U_equal_tmp_146);
  assign mux_698_nl = MUX_s_1_2_2(nor_1353_cse, (nor_1350_nl), nor_326_cse);
  assign mux_699_nl = MUX_s_1_2_2(nor_1353_cse, (mux_698_nl), FpAlu_8U_23U_nor_dfs_48);
  assign nor_1356_nl = ~((~(IsNaN_8U_23U_land_lpi_1_dfm_10 | (~ IsNaN_8U_23U_1_land_lpi_1_dfm_9)
      | (~ FpAlu_8U_23U_nor_dfs_79))) | FpAlu_8U_23U_or_861_itm_4);
  assign nor_1357_nl = ~(FpAlu_8U_23U_nor_dfs_79 | FpAlu_8U_23U_or_861_itm_4);
  assign mux_700_nl = MUX_s_1_2_2((nor_1357_nl), (nor_1356_nl), nor_327_cse);
  assign nor_1355_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      FpAlu_8U_23U_equal_tmp_237 | (mux_700_nl));
  assign mux_701_nl = MUX_s_1_2_2((nor_1355_nl), (mux_699_nl), or_cse_2);
  assign nor_1345_nl = ~((~ FpAdd_8U_23U_mux_242_tmp_49) | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1346_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_204[0]) | (~((cfg_alu_algo_1_sva_st_204[1]) & alu_loop_op_16_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm)));
  assign mux_704_nl = MUX_s_1_2_2((nor_1346_nl), (nor_1345_nl), nor_333_cse);
  assign nor_1347_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7 |
      (cfg_alu_algo_1_sva_st_205[0]) | (~((cfg_alu_algo_1_sva_st_205[1]) & alu_loop_op_16_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2)));
  assign mux_705_nl = MUX_s_1_2_2((nor_1347_nl), (mux_704_nl), or_cse_2);
  assign nor_1338_nl = ~((((~ FpAlu_8U_23U_nor_dfs_48) | IsNaN_8U_23U_land_lpi_1_dfm_9
      | IsNaN_8U_23U_3_land_lpi_1_dfm_7) & FpAlu_8U_23U_equal_tmp_146) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_204!=2'b10));
  assign nor_1339_nl = ~((((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_lpi_1_dfm_10
      | IsNaN_8U_23U_land_lpi_1_dfm_st_5) & FpAlu_8U_23U_equal_tmp_237) | (~ main_stage_v_4)
      | io_read_cfg_alu_bypass_rsc_svs_7 | (cfg_alu_algo_1_sva_st_205!=2'b10));
  assign mux_711_nl = MUX_s_1_2_2((nor_1339_nl), (nor_1338_nl), or_cse_2);
  assign nor_1333_nl = ~((~((~((cfg_alu_algo_1_sva_st_204!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_48)
      | (~ IsNaN_8U_23U_1_land_lpi_1_dfm_8) | IsNaN_8U_23U_land_lpi_1_dfm_9)) | FpAlu_8U_23U_or_861_itm_3))
      | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6 | FpAlu_8U_23U_equal_tmp_146);
  assign nor_1336_nl = ~((~((~((~ FpAlu_8U_23U_nor_dfs_79) | IsNaN_8U_23U_land_lpi_1_dfm_10
      | (cfg_alu_algo_1_sva_st_205!=2'b10) | (~ IsNaN_8U_23U_1_land_lpi_1_dfm_9)))
      | FpAlu_8U_23U_or_861_itm_4)) | (~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_7
      | FpAlu_8U_23U_equal_tmp_237);
  assign mux_717_nl = MUX_s_1_2_2((nor_1336_nl), (nor_1333_nl), or_cse_2);
  assign or_1929_nl = alu_loop_op_16_FpCmp_8U_23U_false_slc_8_1_svs_st_2 | (~ FpAlu_8U_23U_nor_dfs)
      | IsNaN_8U_23U_land_lpi_1_dfm_8 | (reg_cfg_alu_algo_1_sva_st_93_cse[0]) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign mux_806_nl = MUX_s_1_2_2(or_tmp_1915, (or_1929_nl), FpAlu_8U_23U_equal_tmp_1);
  assign mux_808_nl = MUX_s_1_2_2(mux_807_cse, (mux_806_nl), reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign mux_809_nl = MUX_s_1_2_2((mux_808_nl), mux_805_cse, nor_333_cse);
  assign or_1934_nl = IsNaN_8U_23U_land_lpi_1_dfm_9 | (~ FpAlu_8U_23U_nor_dfs_48)
      | IsNaN_8U_23U_3_land_lpi_1_dfm_7 | io_read_cfg_alu_bypass_rsc_svs_st_6 | (~
      main_stage_v_3);
  assign mux_810_nl = MUX_s_1_2_2(or_1935_cse, (or_1934_nl), FpAlu_8U_23U_equal_tmp_146);
  assign or_1936_nl = (cfg_alu_algo_1_sva_st_204[0]) | (mux_810_nl);
  assign mux_812_nl = MUX_s_1_2_2(mux_811_cse, (or_1936_nl), cfg_alu_algo_1_sva_st_204[1]);
  assign mux_813_nl = MUX_s_1_2_2((mux_812_nl), (mux_809_nl), or_cse_2);
  assign nor_1308_nl = ~(((alu_loop_op_15_FpCmp_8U_23U_false_slc_8_svs_st_2 | (~
      FpAlu_8U_23U_nor_dfs) | IsNaN_8U_23U_land_15_lpi_1_dfm_8) & FpAlu_8U_23U_equal_tmp_1)
      | (reg_cfg_alu_algo_1_sva_st_93_cse[0]) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (~ main_stage_v_2));
  assign mux_820_nl = MUX_s_1_2_2(mux_819_cse, (nor_1308_nl), reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign mux_821_nl = MUX_s_1_2_2((mux_820_nl), mux_818_cse, nor_333_cse);
  assign nor_1311_nl = ~(IsNaN_8U_23U_land_15_lpi_1_dfm_9 | (~ FpAlu_8U_23U_nor_dfs_48)
      | IsNaN_8U_23U_3_land_15_lpi_1_dfm_7 | (cfg_alu_algo_1_sva_st_204[0]) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign mux_822_nl = MUX_s_1_2_2(nor_1312_cse, (nor_1311_nl), FpAlu_8U_23U_equal_tmp_146);
  assign mux_824_nl = MUX_s_1_2_2(mux_823_cse, (mux_822_nl), cfg_alu_algo_1_sva_st_204[1]);
  assign mux_825_nl = MUX_s_1_2_2((mux_824_nl), (mux_821_nl), or_cse_2);
  assign nor_1271_nl = ~(((alu_loop_op_8_FpCmp_8U_23U_false_slc_8_1_svs_st_2 | (~
      FpAlu_8U_23U_nor_dfs) | IsNaN_8U_23U_land_8_lpi_1_dfm_8) & FpAlu_8U_23U_equal_tmp_1)
      | (reg_cfg_alu_algo_1_sva_st_93_cse[0]) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (~ main_stage_v_2));
  assign mux_852_nl = MUX_s_1_2_2(mux_819_cse, (nor_1271_nl), reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign mux_853_nl = MUX_s_1_2_2((mux_852_nl), mux_818_cse, nor_333_cse);
  assign or_2030_nl = IsNaN_8U_23U_land_8_lpi_1_dfm_9 | (~ FpAlu_8U_23U_nor_dfs_48)
      | IsNaN_8U_23U_3_land_8_lpi_1_dfm_7 | io_read_cfg_alu_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign mux_854_nl = MUX_s_1_2_2(or_1935_cse, (or_2030_nl), FpAlu_8U_23U_equal_tmp_146);
  assign nor_1274_nl = ~((cfg_alu_algo_1_sva_st_204[0]) | (mux_854_nl));
  assign mux_856_nl = MUX_s_1_2_2(mux_823_cse, (nor_1274_nl), cfg_alu_algo_1_sva_st_204[1]);
  assign mux_857_nl = MUX_s_1_2_2((mux_856_nl), (mux_853_nl), or_cse_2);
  assign or_2051_nl = (~ FpAlu_8U_23U_nor_dfs) | alu_loop_op_7_FpCmp_8U_23U_false_slc_8_svs_st_2
      | IsNaN_8U_23U_land_7_lpi_1_dfm_8 | (reg_cfg_alu_algo_1_sva_st_93_cse[0]) |
      io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign mux_863_nl = MUX_s_1_2_2(or_tmp_1915, (or_2051_nl), FpAlu_8U_23U_equal_tmp_1);
  assign mux_865_nl = MUX_s_1_2_2(mux_807_cse, (mux_863_nl), reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign mux_866_nl = MUX_s_1_2_2((mux_865_nl), mux_805_cse, nor_333_cse);
  assign or_2056_nl = IsNaN_8U_23U_land_7_lpi_1_dfm_9 | (~ FpAlu_8U_23U_nor_dfs_48)
      | IsNaN_8U_23U_3_land_7_lpi_1_dfm_7 | io_read_cfg_alu_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign mux_867_nl = MUX_s_1_2_2(or_1935_cse, (or_2056_nl), FpAlu_8U_23U_equal_tmp_146);
  assign or_2058_nl = (cfg_alu_algo_1_sva_st_204[0]) | (mux_867_nl);
  assign mux_869_nl = MUX_s_1_2_2(mux_811_cse, (or_2058_nl), cfg_alu_algo_1_sva_st_204[1]);
  assign mux_870_nl = MUX_s_1_2_2((mux_869_nl), (mux_866_nl), or_cse_2);
  assign nor_1239_nl = ~(alu_loop_op_3_FpCmp_8U_23U_false_slc_8_svs_st_2 | (~ FpAlu_8U_23U_nor_dfs)
      | IsNaN_8U_23U_land_3_lpi_1_dfm_8 | (reg_cfg_alu_algo_1_sva_st_93_cse[0]) |
      io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign nor_1240_nl = ~((reg_cfg_alu_algo_1_sva_st_93_cse[0]) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (~ main_stage_v_2));
  assign mux_885_nl = MUX_s_1_2_2((nor_1240_nl), (nor_1239_nl), FpAlu_8U_23U_equal_tmp_1);
  assign nor_1241_nl = ~((~(FpAlu_8U_23U_equal_tmp | (reg_cfg_alu_algo_1_sva_st_93_cse[0])))
      | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign nor_1243_nl = ~((~ FpAlu_8U_23U_equal_tmp) | (reg_cfg_alu_algo_1_sva_st_93_cse[0])
      | io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_886_nl = MUX_s_1_2_2((nor_1243_nl), (nor_1241_nl), FpAlu_8U_23U_equal_tmp_2);
  assign mux_887_nl = MUX_s_1_2_2((mux_886_nl), (mux_885_nl), reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign mux_888_nl = MUX_s_1_2_2((mux_887_nl), mux_818_cse, nor_333_cse);
  assign nor_1244_nl = ~(IsNaN_8U_23U_land_3_lpi_1_dfm_9 | (~ FpAlu_8U_23U_nor_dfs_48)
      | IsNaN_8U_23U_3_land_3_lpi_1_dfm_7 | (cfg_alu_algo_1_sva_st_204[0]) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign mux_889_nl = MUX_s_1_2_2(nor_1312_cse, (nor_1244_nl), FpAlu_8U_23U_equal_tmp_146);
  assign mux_891_nl = MUX_s_1_2_2(mux_823_cse, (mux_889_nl), cfg_alu_algo_1_sva_st_204[1]);
  assign mux_892_nl = MUX_s_1_2_2((mux_891_nl), (mux_888_nl), or_cse_2);
  assign or_2132_nl = (~ FpAlu_8U_23U_nor_dfs) | alu_loop_op_1_FpCmp_8U_23U_false_slc_8_svs_st_2
      | IsNaN_8U_23U_land_1_lpi_1_dfm_8 | (reg_cfg_alu_algo_1_sva_st_93_cse[0]) |
      io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign mux_901_nl = MUX_s_1_2_2(or_tmp_1915, (or_2132_nl), FpAlu_8U_23U_equal_tmp_1);
  assign mux_903_nl = MUX_s_1_2_2(mux_807_cse, (mux_901_nl), reg_cfg_alu_algo_1_sva_st_93_cse[1]);
  assign mux_904_nl = MUX_s_1_2_2((mux_903_nl), mux_805_cse, nor_333_cse);
  assign or_2137_nl = (~ FpAlu_8U_23U_equal_tmp_148) | (cfg_alu_algo_1_sva_st_204[1])
      | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign or_2138_nl = IsNaN_8U_23U_land_1_lpi_1_dfm_9 | (~ FpAlu_8U_23U_nor_dfs_48)
      | IsNaN_8U_23U_3_land_1_lpi_1_dfm_7 | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign mux_905_nl = MUX_s_1_2_2(or_1935_cse, (or_2138_nl), FpAlu_8U_23U_equal_tmp_146);
  assign mux_906_nl = MUX_s_1_2_2(or_1938_cse, (mux_905_nl), cfg_alu_algo_1_sva_st_204[1]);
  assign mux_907_nl = MUX_s_1_2_2((mux_906_nl), (or_2137_nl), cfg_alu_algo_1_sva_st_204[0]);
  assign mux_908_nl = MUX_s_1_2_2((mux_907_nl), (mux_904_nl), or_cse_2);
  assign nl_AluOut_data_15_sva_7 = conv_s2s_32_33(AluIn_data_sva_501[511:480]) +
      conv_s2s_32_33({IntShiftLeft_16U_6U_32U_return_31_sva_2 , IntShiftLeft_16U_6U_32U_return_30_1_sva_2
      , IntShiftLeft_16U_6U_32U_return_0_sva_2});
  assign nl_AluOut_data_14_sva_7 = conv_s2s_32_33(AluIn_data_sva_501[479:448]) +
      conv_s2s_32_33({IntShiftLeft_16U_6U_32U_return_31_15_sva_2 , IntShiftLeft_16U_6U_32U_return_30_1_15_sva_2
      , IntShiftLeft_16U_6U_32U_return_0_15_sva_2});
  assign nl_AluOut_data_13_sva_7 = conv_s2s_32_33(AluIn_data_sva_501[447:416]) +
      conv_s2s_32_33({IntShiftLeft_16U_6U_32U_return_31_14_sva_2 , IntShiftLeft_16U_6U_32U_return_30_1_14_sva_2
      , IntShiftLeft_16U_6U_32U_return_0_14_sva_2});
  assign nl_AluOut_data_12_sva_7 = conv_s2s_32_33(AluIn_data_sva_501[415:384]) +
      conv_s2s_32_33({IntShiftLeft_16U_6U_32U_return_31_13_sva_2 , IntShiftLeft_16U_6U_32U_return_30_1_13_sva_2
      , IntShiftLeft_16U_6U_32U_return_0_13_sva_2});
  assign nl_AluOut_data_11_sva_7 = conv_s2s_32_33(AluIn_data_sva_501[383:352]) +
      conv_s2s_32_33({IntShiftLeft_16U_6U_32U_return_31_12_sva_2 , IntShiftLeft_16U_6U_32U_return_30_1_12_sva_2
      , IntShiftLeft_16U_6U_32U_return_0_12_sva_2});
  assign nl_AluOut_data_10_sva_7 = conv_s2s_32_33(AluIn_data_sva_501[351:320]) +
      conv_s2s_32_33({IntShiftLeft_16U_6U_32U_return_31_11_sva_2 , IntShiftLeft_16U_6U_32U_return_30_1_11_sva_2
      , IntShiftLeft_16U_6U_32U_return_0_11_sva_2});
  assign nl_AluOut_data_9_sva_7 = conv_s2s_32_33(AluIn_data_sva_501[319:288]) +
      conv_s2s_32_33({IntShiftLeft_16U_6U_32U_return_31_10_sva_2 , IntShiftLeft_16U_6U_32U_return_30_1_10_sva_2
      , IntShiftLeft_16U_6U_32U_return_0_10_sva_2});
  assign nl_AluOut_data_8_sva_7 = conv_s2s_32_33(AluIn_data_sva_501[287:256]) +
      conv_s2s_32_33({IntShiftLeft_16U_6U_32U_return_31_9_sva_2 , IntShiftLeft_16U_6U_32U_return_30_1_9_sva_2
      , IntShiftLeft_16U_6U_32U_return_0_9_sva_2});
  assign nl_AluOut_data_7_sva_7 = conv_s2s_32_33(AluIn_data_sva_501[255:224]) +
      conv_s2s_32_33({IntShiftLeft_16U_6U_32U_return_31_8_sva_2 , IntShiftLeft_16U_6U_32U_return_30_1_8_sva_2
      , IntShiftLeft_16U_6U_32U_return_0_8_sva_2});
  assign nl_AluOut_data_6_sva_7 = conv_s2s_32_33(AluIn_data_sva_501[223:192]) +
      conv_s2s_32_33({IntShiftLeft_16U_6U_32U_return_31_7_sva_2 , IntShiftLeft_16U_6U_32U_return_30_1_7_sva_2
      , IntShiftLeft_16U_6U_32U_return_0_7_sva_2});
  assign nl_AluOut_data_5_sva_7 = conv_s2s_32_33(AluIn_data_sva_501[191:160]) +
      conv_s2s_32_33({IntShiftLeft_16U_6U_32U_return_31_6_sva_2 , IntShiftLeft_16U_6U_32U_return_30_1_6_sva_2
      , IntShiftLeft_16U_6U_32U_return_0_6_sva_2});
  assign nl_AluOut_data_4_sva_7 = conv_s2s_32_33(AluIn_data_sva_501[159:128]) +
      conv_s2s_32_33({IntShiftLeft_16U_6U_32U_return_31_5_sva_2 , IntShiftLeft_16U_6U_32U_return_30_1_5_sva_2
      , IntShiftLeft_16U_6U_32U_return_0_5_sva_2});
  assign nl_AluOut_data_3_sva_7 = conv_s2s_32_33(AluIn_data_sva_501[127:96]) + conv_s2s_32_33({IntShiftLeft_16U_6U_32U_return_31_4_sva_2
      , IntShiftLeft_16U_6U_32U_return_30_1_4_sva_2 , IntShiftLeft_16U_6U_32U_return_0_4_sva_2});
  assign nl_AluOut_data_2_sva_7 = conv_s2s_32_33(AluIn_data_sva_501[95:64]) + conv_s2s_32_33({IntShiftLeft_16U_6U_32U_return_31_3_sva_2
      , IntShiftLeft_16U_6U_32U_return_30_1_3_sva_2 , IntShiftLeft_16U_6U_32U_return_0_3_sva_2});
  assign nl_AluOut_data_1_sva_7 = conv_s2s_32_33(AluIn_data_sva_501[63:32]) + conv_s2s_32_33({IntShiftLeft_16U_6U_32U_return_31_2_sva_2
      , IntShiftLeft_16U_6U_32U_return_30_1_2_sva_2 , IntShiftLeft_16U_6U_32U_return_0_2_sva_2});
  assign nl_AluOut_data_0_sva_7 = conv_s2s_32_33(AluIn_data_sva_501[31:0]) + conv_s2s_32_33({IntShiftLeft_16U_6U_32U_return_31_1_sva_2
      , IntShiftLeft_16U_6U_32U_return_30_1_1_sva_2 , IntShiftLeft_16U_6U_32U_return_0_1_sva_2});
  assign IsNaN_8U_23U_3_aelse_or_nl = and_1318_cse | and_1307_cse;
  assign nor_931_nl = ~((~ FpCmp_8U_23U_true_if_acc_18_itm_8_1) | (cfg_precision!=2'b10)
      | io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign mux_1358_nl = MUX_s_1_2_2((nor_931_nl), or_tmp_24, reg_alu_loop_op_2_FpAdd_8U_23U_is_a_greater_slc_8_1_svs_cse);
  assign or_2821_nl = (~ and_89_tmp) | (cfg_alu_algo_1_sva_st_92!=2'b10);
  assign mux_1359_nl = MUX_s_1_2_2((mux_1358_nl), reg_alu_loop_op_2_FpAdd_8U_23U_is_a_greater_slc_8_1_svs_cse,
      or_2821_nl);
  assign and_1917_nl = (or_dcpl_14 | or_dcpl_295 | IsNaN_8U_23U_2_land_8_lpi_1_dfm_st_1)
      & and_89_tmp;
  assign FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_16_nl = ~((fsm_output[1])
      & (FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49]));
  assign FpAdd_8U_23U_if_3_if_mux_64_nl = MUX_v_6_2_2(6'b1, (~ IntLeadZero_49U_leading_sign_49_0_rtn_1_sva_2),
      FpNormalize_8U_49U_else_and_tmp);
  assign nl_acc_nl = ({FpAdd_8U_23U_qr_2_lpi_1_dfm_5_7_4_1 , FpAdd_8U_23U_qr_2_lpi_1_dfm_5_3_0_1
      , (FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_16_nl)}) + conv_s2u_8_9({FpNormalize_8U_49U_else_and_tmp
      , (FpAdd_8U_23U_if_3_if_mux_64_nl) , 1'b1});
  assign acc_nl = nl_acc_nl[8:0];
  assign z_out = readslicef_9_8_1((acc_nl));
  assign FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_17_nl = ~((fsm_output[1])
      & (FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49]));
  assign FpAdd_8U_23U_if_3_if_mux_65_nl = MUX_v_6_2_2(6'b1, (~ IntLeadZero_49U_leading_sign_49_0_rtn_2_sva_2),
      FpNormalize_8U_49U_else_and_tmp_1);
  assign nl_acc_1_nl = ({FpAdd_8U_23U_qr_3_lpi_1_dfm_5_7_4_1 , FpAdd_8U_23U_qr_3_lpi_1_dfm_5_3_0_1
      , (FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_17_nl)}) + conv_s2u_8_9({FpNormalize_8U_49U_else_and_tmp_1
      , (FpAdd_8U_23U_if_3_if_mux_65_nl) , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[8:0];
  assign z_out_1 = readslicef_9_8_1((acc_1_nl));
  assign FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_18_nl = ~((fsm_output[1])
      & (FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49]));
  assign FpAdd_8U_23U_if_3_if_mux_66_nl = MUX_v_6_2_2(6'b1, (~ IntLeadZero_49U_leading_sign_49_0_rtn_3_sva_2),
      FpNormalize_8U_49U_else_and_tmp_2);
  assign nl_acc_2_nl = ({FpAdd_8U_23U_qr_4_lpi_1_dfm_5_7_4_1 , FpAdd_8U_23U_qr_4_lpi_1_dfm_5_3_0_1
      , (FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_18_nl)}) + conv_s2u_8_9({FpNormalize_8U_49U_else_and_tmp_2
      , (FpAdd_8U_23U_if_3_if_mux_66_nl) , 1'b1});
  assign acc_2_nl = nl_acc_2_nl[8:0];
  assign z_out_2 = readslicef_9_8_1((acc_2_nl));
  assign FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_19_nl = ~((fsm_output[1])
      & (FpAdd_8U_23U_int_mant_p1_4_lpi_1_dfm_5[49]));
  assign FpAdd_8U_23U_if_3_if_mux_67_nl = MUX_v_6_2_2(6'b1, (~ IntLeadZero_49U_leading_sign_49_0_rtn_4_sva_2),
      FpNormalize_8U_49U_else_and_tmp_3);
  assign nl_acc_3_nl = ({FpAdd_8U_23U_qr_5_lpi_1_dfm_5_7_4_1 , FpAdd_8U_23U_qr_5_lpi_1_dfm_5_3_0_1
      , (FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_19_nl)}) + conv_s2u_8_9({FpNormalize_8U_49U_else_and_tmp_3
      , (FpAdd_8U_23U_if_3_if_mux_67_nl) , 1'b1});
  assign acc_3_nl = nl_acc_3_nl[8:0];
  assign z_out_3 = readslicef_9_8_1((acc_3_nl));
  assign FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_20_nl = ~((fsm_output[1])
      & (FpAdd_8U_23U_int_mant_p1_5_lpi_1_dfm_5[49]));
  assign FpAdd_8U_23U_if_3_if_mux_68_nl = MUX_v_6_2_2(6'b1, (~ IntLeadZero_49U_leading_sign_49_0_rtn_5_sva_2),
      FpNormalize_8U_49U_else_and_tmp_4);
  assign nl_acc_4_nl = ({FpAdd_8U_23U_qr_6_lpi_1_dfm_5_7_4_1 , FpAdd_8U_23U_qr_6_lpi_1_dfm_5_3_0_1
      , (FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_20_nl)}) + conv_s2u_8_9({FpNormalize_8U_49U_else_and_tmp_4
      , (FpAdd_8U_23U_if_3_if_mux_68_nl) , 1'b1});
  assign acc_4_nl = nl_acc_4_nl[8:0];
  assign z_out_4 = readslicef_9_8_1((acc_4_nl));
  assign FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_21_nl = ~((fsm_output[1])
      & (FpAdd_8U_23U_int_mant_p1_6_lpi_1_dfm_5[49]));
  assign FpAdd_8U_23U_if_3_if_mux_69_nl = MUX_v_6_2_2(6'b1, (~ IntLeadZero_49U_leading_sign_49_0_rtn_6_sva_2),
      FpNormalize_8U_49U_else_and_tmp_5);
  assign nl_acc_5_nl = ({FpAdd_8U_23U_qr_7_lpi_1_dfm_5_7_4_1 , FpAdd_8U_23U_qr_7_lpi_1_dfm_5_3_0_1
      , (FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_21_nl)}) + conv_s2u_8_9({FpNormalize_8U_49U_else_and_tmp_5
      , (FpAdd_8U_23U_if_3_if_mux_69_nl) , 1'b1});
  assign acc_5_nl = nl_acc_5_nl[8:0];
  assign z_out_5 = readslicef_9_8_1((acc_5_nl));
  assign FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_22_nl = ~((fsm_output[1])
      & (FpAdd_8U_23U_int_mant_p1_7_lpi_1_dfm_5[49]));
  assign FpAdd_8U_23U_if_3_if_mux_70_nl = MUX_v_6_2_2(6'b1, (~ IntLeadZero_49U_leading_sign_49_0_rtn_7_sva_2),
      FpNormalize_8U_49U_else_and_tmp_6);
  assign nl_acc_6_nl = ({FpAdd_8U_23U_qr_8_lpi_1_dfm_5_7_4_1 , FpAdd_8U_23U_qr_8_lpi_1_dfm_5_3_0_1
      , (FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_22_nl)}) + conv_s2u_8_9({FpNormalize_8U_49U_else_and_tmp_6
      , (FpAdd_8U_23U_if_3_if_mux_70_nl) , 1'b1});
  assign acc_6_nl = nl_acc_6_nl[8:0];
  assign z_out_6 = readslicef_9_8_1((acc_6_nl));
  assign FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_23_nl = ~((fsm_output[1])
      & (FpAdd_8U_23U_int_mant_p1_8_lpi_1_dfm_5[49]));
  assign FpAdd_8U_23U_if_3_if_mux_71_nl = MUX_v_6_2_2(6'b1, (~ IntLeadZero_49U_leading_sign_49_0_rtn_8_sva_2),
      FpNormalize_8U_49U_else_and_tmp_7);
  assign nl_acc_7_nl = ({FpAdd_8U_23U_qr_9_lpi_1_dfm_5_7_4_1 , FpAdd_8U_23U_qr_9_lpi_1_dfm_5_3_0_1
      , (FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_23_nl)}) + conv_s2u_8_9({FpNormalize_8U_49U_else_and_tmp_7
      , (FpAdd_8U_23U_if_3_if_mux_71_nl) , 1'b1});
  assign acc_7_nl = nl_acc_7_nl[8:0];
  assign z_out_7 = readslicef_9_8_1((acc_7_nl));
  assign FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_24_nl = ~((fsm_output[1])
      & (FpAdd_8U_23U_int_mant_p1_9_lpi_1_dfm_5[49]));
  assign FpAdd_8U_23U_if_3_if_mux_72_nl = MUX_v_6_2_2(6'b1, (~ IntLeadZero_49U_leading_sign_49_0_rtn_9_sva_2),
      FpNormalize_8U_49U_else_and_tmp_8);
  assign nl_acc_8_nl = ({FpAdd_8U_23U_qr_10_lpi_1_dfm_5_7_4_1 , FpAdd_8U_23U_qr_10_lpi_1_dfm_5_3_0_1
      , (FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_24_nl)}) + conv_s2u_8_9({FpNormalize_8U_49U_else_and_tmp_8
      , (FpAdd_8U_23U_if_3_if_mux_72_nl) , 1'b1});
  assign acc_8_nl = nl_acc_8_nl[8:0];
  assign z_out_8 = readslicef_9_8_1((acc_8_nl));
  assign FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_25_nl = ~((fsm_output[1])
      & (FpAdd_8U_23U_int_mant_p1_10_lpi_1_dfm_5[49]));
  assign FpAdd_8U_23U_if_3_if_mux_73_nl = MUX_v_6_2_2(6'b1, (~ IntLeadZero_49U_leading_sign_49_0_rtn_10_sva_2),
      FpNormalize_8U_49U_else_and_tmp_9);
  assign nl_acc_9_nl = ({FpAdd_8U_23U_qr_11_lpi_1_dfm_5_7_4_1 , FpAdd_8U_23U_qr_11_lpi_1_dfm_5_3_0_1
      , (FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_25_nl)}) + conv_s2u_8_9({FpNormalize_8U_49U_else_and_tmp_9
      , (FpAdd_8U_23U_if_3_if_mux_73_nl) , 1'b1});
  assign acc_9_nl = nl_acc_9_nl[8:0];
  assign z_out_9 = readslicef_9_8_1((acc_9_nl));
  assign FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_26_nl = ~((fsm_output[1])
      & (FpAdd_8U_23U_int_mant_p1_11_lpi_1_dfm_5[49]));
  assign FpAdd_8U_23U_if_3_if_mux_74_nl = MUX_v_6_2_2(6'b1, (~ IntLeadZero_49U_leading_sign_49_0_rtn_11_sva_2),
      FpNormalize_8U_49U_else_and_tmp_10);
  assign nl_acc_10_nl = ({FpAdd_8U_23U_qr_12_lpi_1_dfm_5_7_4_1 , FpAdd_8U_23U_qr_12_lpi_1_dfm_5_3_0_1
      , (FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_26_nl)}) + conv_s2u_8_9({FpNormalize_8U_49U_else_and_tmp_10
      , (FpAdd_8U_23U_if_3_if_mux_74_nl) , 1'b1});
  assign acc_10_nl = nl_acc_10_nl[8:0];
  assign z_out_10 = readslicef_9_8_1((acc_10_nl));
  assign FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_27_nl = ~((fsm_output[1])
      & (FpAdd_8U_23U_int_mant_p1_12_lpi_1_dfm_5[49]));
  assign FpAdd_8U_23U_if_3_if_mux_75_nl = MUX_v_6_2_2(6'b1, (~ IntLeadZero_49U_leading_sign_49_0_rtn_12_sva_2),
      FpNormalize_8U_49U_else_and_tmp_11);
  assign nl_acc_11_nl = ({FpAdd_8U_23U_qr_13_lpi_1_dfm_5_7_4_1 , FpAdd_8U_23U_qr_13_lpi_1_dfm_5_3_0_1
      , (FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_27_nl)}) + conv_s2u_8_9({FpNormalize_8U_49U_else_and_tmp_11
      , (FpAdd_8U_23U_if_3_if_mux_75_nl) , 1'b1});
  assign acc_11_nl = nl_acc_11_nl[8:0];
  assign z_out_11 = readslicef_9_8_1((acc_11_nl));
  assign FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_28_nl = ~((fsm_output[1])
      & (FpAdd_8U_23U_int_mant_p1_13_lpi_1_dfm_5[49]));
  assign FpAdd_8U_23U_if_3_if_mux_76_nl = MUX_v_6_2_2(6'b1, (~ IntLeadZero_49U_leading_sign_49_0_rtn_13_sva_2),
      FpNormalize_8U_49U_else_and_tmp_12);
  assign nl_acc_12_nl = ({FpAdd_8U_23U_qr_14_lpi_1_dfm_5_7_4_1 , FpAdd_8U_23U_qr_14_lpi_1_dfm_5_3_0_1
      , (FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_28_nl)}) + conv_s2u_8_9({FpNormalize_8U_49U_else_and_tmp_12
      , (FpAdd_8U_23U_if_3_if_mux_76_nl) , 1'b1});
  assign acc_12_nl = nl_acc_12_nl[8:0];
  assign z_out_12 = readslicef_9_8_1((acc_12_nl));
  assign FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_29_nl = ~((fsm_output[1])
      & (FpAdd_8U_23U_int_mant_p1_14_lpi_1_dfm_5[49]));
  assign FpAdd_8U_23U_if_3_if_mux_77_nl = MUX_v_6_2_2(6'b1, (~ IntLeadZero_49U_leading_sign_49_0_rtn_14_sva_2),
      FpNormalize_8U_49U_else_and_tmp_13);
  assign nl_acc_13_nl = ({FpAdd_8U_23U_qr_15_lpi_1_dfm_5_7_4_1 , FpAdd_8U_23U_qr_15_lpi_1_dfm_5_3_0_1
      , (FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_29_nl)}) + conv_s2u_8_9({FpNormalize_8U_49U_else_and_tmp_13
      , (FpAdd_8U_23U_if_3_if_mux_77_nl) , 1'b1});
  assign acc_13_nl = nl_acc_13_nl[8:0];
  assign z_out_13 = readslicef_9_8_1((acc_13_nl));
  assign FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_30_nl = ~((fsm_output[1])
      & (FpAdd_8U_23U_int_mant_p1_15_lpi_1_dfm_5[49]));
  assign FpAdd_8U_23U_if_3_if_mux_78_nl = MUX_v_6_2_2(6'b1, (~ IntLeadZero_49U_leading_sign_49_0_rtn_15_sva_2),
      FpNormalize_8U_49U_else_and_tmp_14);
  assign nl_acc_14_nl = ({FpAdd_8U_23U_qr_16_lpi_1_dfm_5_7_4_1 , FpAdd_8U_23U_qr_16_lpi_1_dfm_5_3_0_1
      , (FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_30_nl)}) + conv_s2u_8_9({FpNormalize_8U_49U_else_and_tmp_14
      , (FpAdd_8U_23U_if_3_if_mux_78_nl) , 1'b1});
  assign acc_14_nl = nl_acc_14_nl[8:0];
  assign z_out_14 = readslicef_9_8_1((acc_14_nl));
  assign FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_31_nl = ~((fsm_output[1])
      & (FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49]));
  assign FpAdd_8U_23U_if_3_if_mux_79_nl = MUX_v_6_2_2(6'b1, (~ IntLeadZero_49U_leading_sign_49_0_rtn_sva_2),
      FpNormalize_8U_49U_else_and_tmp_15);
  assign nl_acc_15_nl = ({FpAdd_8U_23U_qr_lpi_1_dfm_5_7_4_1 , FpAdd_8U_23U_qr_lpi_1_dfm_5_3_0_1
      , (FpAdd_8U_23U_if_3_if_FpAdd_8U_23U_if_3_if_nand_31_nl)}) + conv_s2u_8_9({FpNormalize_8U_49U_else_and_tmp_15
      , (FpAdd_8U_23U_if_3_if_mux_79_nl) , 1'b1});
  assign acc_15_nl = nl_acc_15_nl[8:0];
  assign z_out_15 = readslicef_9_8_1((acc_15_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_32_nl = MUX_v_8_2_2((AluIn_data_sva_501[30:23]),
      ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_9}),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_33_nl = MUX_v_8_2_2(({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_9)}), (~ (AluIn_data_sva_501[30:23])),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp);
  assign nl_acc_16_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_32_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_33_nl)
      , 1'b1});
  assign acc_16_nl = nl_acc_16_nl[8:0];
  assign z_out_16 = readslicef_9_8_1((acc_16_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_34_nl = MUX_v_8_2_2((AluIn_data_sva_501[510:503]),
      ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_9}),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_1);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_35_nl = MUX_v_8_2_2(({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_9)}), (~ (AluIn_data_sva_501[510:503])),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_1);
  assign nl_acc_17_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_34_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_35_nl)
      , 1'b1});
  assign acc_17_nl = nl_acc_17_nl[8:0];
  assign z_out_17 = readslicef_9_8_1((acc_17_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_36_nl = MUX_v_8_2_2((AluIn_data_sva_501[62:55]),
      ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_9}),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_2);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_37_nl = MUX_v_8_2_2(({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_9)}), (~ (AluIn_data_sva_501[62:55])),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_2);
  assign nl_acc_18_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_36_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_37_nl)
      , 1'b1});
  assign acc_18_nl = nl_acc_18_nl[8:0];
  assign z_out_18 = readslicef_9_8_1((acc_18_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_38_nl = MUX_v_8_2_2((AluIn_data_sva_501[478:471]),
      ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_9}),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_3);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_39_nl = MUX_v_8_2_2(({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_9)}), (~ (AluIn_data_sva_501[478:471])),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_3);
  assign nl_acc_19_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_38_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_39_nl)
      , 1'b1});
  assign acc_19_nl = nl_acc_19_nl[8:0];
  assign z_out_19 = readslicef_9_8_1((acc_19_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_40_nl = MUX_v_8_2_2((AluIn_data_sva_501[94:87]),
      ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_9}),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_4);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_41_nl = MUX_v_8_2_2(({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_9)}), (~ (AluIn_data_sva_501[94:87])),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_4);
  assign nl_acc_20_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_40_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_41_nl)
      , 1'b1});
  assign acc_20_nl = nl_acc_20_nl[8:0];
  assign z_out_20 = readslicef_9_8_1((acc_20_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_42_nl = MUX_v_8_2_2((AluIn_data_sva_501[446:439]),
      ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_9}),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_5);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_43_nl = MUX_v_8_2_2(({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_9)}), (~ (AluIn_data_sva_501[446:439])),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_5);
  assign nl_acc_21_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_42_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_43_nl)
      , 1'b1});
  assign acc_21_nl = nl_acc_21_nl[8:0];
  assign z_out_21 = readslicef_9_8_1((acc_21_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_44_nl = MUX_v_8_2_2((AluIn_data_sva_501[126:119]),
      ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_9}),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_6);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_45_nl = MUX_v_8_2_2(({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_9)}), (~ (AluIn_data_sva_501[126:119])),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_6);
  assign nl_acc_22_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_44_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_45_nl)
      , 1'b1});
  assign acc_22_nl = nl_acc_22_nl[8:0];
  assign z_out_22 = readslicef_9_8_1((acc_22_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_46_nl = MUX_v_8_2_2((AluIn_data_sva_501[414:407]),
      ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_9}),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_7);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_47_nl = MUX_v_8_2_2(({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_9)}), (~ (AluIn_data_sva_501[414:407])),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_7);
  assign nl_acc_23_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_46_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_47_nl)
      , 1'b1});
  assign acc_23_nl = nl_acc_23_nl[8:0];
  assign z_out_23 = readslicef_9_8_1((acc_23_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_48_nl = MUX_v_8_2_2((AluIn_data_sva_501[158:151]),
      ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_9}),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_8);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_49_nl = MUX_v_8_2_2(({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_9)}), (~ (AluIn_data_sva_501[158:151])),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_8);
  assign nl_acc_24_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_48_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_49_nl)
      , 1'b1});
  assign acc_24_nl = nl_acc_24_nl[8:0];
  assign z_out_24 = readslicef_9_8_1((acc_24_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_50_nl = MUX_v_8_2_2((AluIn_data_sva_501[382:375]),
      ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_9}),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_9);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_51_nl = MUX_v_8_2_2(({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_9)}), (~ (AluIn_data_sva_501[382:375])),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_9);
  assign nl_acc_25_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_50_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_51_nl)
      , 1'b1});
  assign acc_25_nl = nl_acc_25_nl[8:0];
  assign z_out_25 = readslicef_9_8_1((acc_25_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_52_nl = MUX_v_8_2_2((AluIn_data_sva_501[190:183]),
      ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_9}),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_10);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_53_nl = MUX_v_8_2_2(({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_9)}), (~ (AluIn_data_sva_501[190:183])),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_10);
  assign nl_acc_26_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_52_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_53_nl)
      , 1'b1});
  assign acc_26_nl = nl_acc_26_nl[8:0];
  assign z_out_26 = readslicef_9_8_1((acc_26_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_54_nl = MUX_v_8_2_2((AluIn_data_sva_501[350:343]),
      ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_9}),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_11);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_55_nl = MUX_v_8_2_2(({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_9)}), (~ (AluIn_data_sva_501[350:343])),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_11);
  assign nl_acc_27_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_54_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_55_nl)
      , 1'b1});
  assign acc_27_nl = nl_acc_27_nl[8:0];
  assign z_out_27 = readslicef_9_8_1((acc_27_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_56_nl = MUX_v_8_2_2((AluIn_data_sva_501[222:215]),
      ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_9}),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_12);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_57_nl = MUX_v_8_2_2(({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_9)}), (~ (AluIn_data_sva_501[222:215])),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_12);
  assign nl_acc_28_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_56_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_57_nl)
      , 1'b1});
  assign acc_28_nl = nl_acc_28_nl[8:0];
  assign z_out_28 = readslicef_9_8_1((acc_28_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_58_nl = MUX_v_8_2_2((AluIn_data_sva_501[318:311]),
      ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_9}),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_13);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_59_nl = MUX_v_8_2_2(({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_9)}), (~ (AluIn_data_sva_501[318:311])),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_13);
  assign nl_acc_29_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_58_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_59_nl)
      , 1'b1});
  assign acc_29_nl = nl_acc_29_nl[8:0];
  assign z_out_29 = readslicef_9_8_1((acc_29_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_60_nl = MUX_v_8_2_2((AluIn_data_sva_501[254:247]),
      ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_9}),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_14);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_61_nl = MUX_v_8_2_2(({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_9)}), (~ (AluIn_data_sva_501[254:247])),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_14);
  assign nl_acc_30_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_60_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_61_nl)
      , 1'b1});
  assign acc_30_nl = nl_acc_30_nl[8:0];
  assign z_out_30 = readslicef_9_8_1((acc_30_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_62_nl = MUX_v_8_2_2((AluIn_data_sva_501[286:279]),
      ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_9 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_9}),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_15);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_63_nl = MUX_v_8_2_2(({(~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_9)
      , (~ FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_9)}), (~ (AluIn_data_sva_501[286:279])),
      FpAdd_8U_23U_a_right_shift_qelse_and_tmp_15);
  assign nl_acc_31_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_62_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_63_nl)
      , 1'b1});
  assign acc_31_nl = nl_acc_31_nl[8:0];
  assign z_out_31 = readslicef_9_8_1((acc_31_nl));
  function [0:0] MUX1HOT_s_1_1_2;
    input [0:0] input_0;
    input [0:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction
  function [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction
  function [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction
  function [0:0] MUX1HOT_s_1_5_2;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [4:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction
  function [0:0] MUX1HOT_s_1_7_2;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [6:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    MUX1HOT_s_1_7_2 = result;
  end
  endfunction
  function [9:0] MUX1HOT_v_10_3_2;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [2:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    MUX1HOT_v_10_3_2 = result;
  end
  endfunction
  function [21:0] MUX1HOT_v_22_3_2;
    input [21:0] input_2;
    input [21:0] input_1;
    input [21:0] input_0;
    input [2:0] sel;
    reg [21:0] result;
  begin
    result = input_0 & {22{sel[0]}};
    result = result | ( input_1 & {22{sel[1]}});
    result = result | ( input_2 & {22{sel[2]}});
    MUX1HOT_v_22_3_2 = result;
  end
  endfunction
  function [21:0] MUX1HOT_v_22_4_2;
    input [21:0] input_3;
    input [21:0] input_2;
    input [21:0] input_1;
    input [21:0] input_0;
    input [3:0] sel;
    reg [21:0] result;
  begin
    result = input_0 & {22{sel[0]}};
    result = result | ( input_1 & {22{sel[1]}});
    result = result | ( input_2 & {22{sel[2]}});
    result = result | ( input_3 & {22{sel[3]}});
    MUX1HOT_v_22_4_2 = result;
  end
  endfunction
  function [22:0] MUX1HOT_v_23_3_2;
    input [22:0] input_2;
    input [22:0] input_1;
    input [22:0] input_0;
    input [2:0] sel;
    reg [22:0] result;
  begin
    result = input_0 & {23{sel[0]}};
    result = result | ( input_1 & {23{sel[1]}});
    result = result | ( input_2 & {23{sel[2]}});
    MUX1HOT_v_23_3_2 = result;
  end
  endfunction
  function [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    result = result | ( input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction
  function [29:0] MUX1HOT_v_30_3_2;
    input [29:0] input_2;
    input [29:0] input_1;
    input [29:0] input_0;
    input [2:0] sel;
    reg [29:0] result;
  begin
    result = input_0 & {30{sel[0]}};
    result = result | ( input_1 & {30{sel[1]}});
    result = result | ( input_2 & {30{sel[2]}});
    MUX1HOT_v_30_3_2 = result;
  end
  endfunction
  function [29:0] MUX1HOT_v_30_4_2;
    input [29:0] input_3;
    input [29:0] input_2;
    input [29:0] input_1;
    input [29:0] input_0;
    input [3:0] sel;
    reg [29:0] result;
  begin
    result = input_0 & {30{sel[0]}};
    result = result | ( input_1 & {30{sel[1]}});
    result = result | ( input_2 & {30{sel[2]}});
    result = result | ( input_3 & {30{sel[3]}});
    MUX1HOT_v_30_4_2 = result;
  end
  endfunction
  function [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction
  function [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction
  function [3:0] MUX1HOT_v_4_5_2;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [4:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    result = result | ( input_4 & {4{sel[4]}});
    MUX1HOT_v_4_5_2 = result;
  end
  endfunction
  function [49:0] MUX1HOT_v_50_3_2;
    input [49:0] input_2;
    input [49:0] input_1;
    input [49:0] input_0;
    input [2:0] sel;
    reg [49:0] result;
  begin
    result = input_0 & {50{sel[0]}};
    result = result | ( input_1 & {50{sel[1]}});
    result = result | ( input_2 & {50{sel[2]}});
    MUX1HOT_v_50_3_2 = result;
  end
  endfunction
  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction
  function [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction
  function [21:0] MUX_v_22_2_2;
    input [21:0] input_0;
    input [21:0] input_1;
    input [0:0] sel;
    reg [21:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_22_2_2 = result;
  end
  endfunction
  function [22:0] MUX_v_23_2_2;
    input [22:0] input_0;
    input [22:0] input_1;
    input [0:0] sel;
    reg [22:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_23_2_2 = result;
  end
  endfunction
  function [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction
  function [29:0] MUX_v_30_2_2;
    input [29:0] input_0;
    input [29:0] input_1;
    input [0:0] sel;
    reg [29:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_30_2_2 = result;
  end
  endfunction
  function [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction
  function [48:0] MUX_v_49_2_2;
    input [48:0] input_0;
    input [48:0] input_1;
    input [0:0] sel;
    reg [48:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_49_2_2 = result;
  end
  endfunction
  function [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction
  function [49:0] MUX_v_50_2_2;
    input [49:0] input_0;
    input [49:0] input_1;
    input [0:0] sel;
    reg [49:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_50_2_2 = result;
  end
  endfunction
  function [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction
  function [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction
  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction
  function [0:0] readslicef_24_1_23;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 23;
    readslicef_24_1_23 = tmp[0:0];
  end
  endfunction
  function [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction
  function [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction
  function [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction
  function [7:0] readslicef_9_8_1;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_9_8_1 = tmp[7:0];
  end
  endfunction
  function [1:0] signext_2_1;
    input [0:0] vector;
  begin
    signext_2_1= {{1{vector[0]}}, vector};
  end
  endfunction
  function [32:0] conv_s2s_32_33 ;
    input [31:0] vector ;
  begin
    conv_s2s_32_33 = {vector[31], vector};
  end
  endfunction
  function [8:0] conv_s2u_8_9 ;
    input [7:0] vector ;
  begin
    conv_s2u_8_9 = {vector[7], vector};
  end
  endfunction
  function [32:0] conv_s2u_32_33 ;
    input [31:0] vector ;
  begin
    conv_s2u_32_33 = {vector[31], vector};
  end
  endfunction
  function [8:0] conv_u2s_6_9 ;
    input [5:0] vector ;
  begin
    conv_u2s_6_9 = {{3{1'b0}}, vector};
  end
  endfunction
  function [22:0] conv_u2u_1_23 ;
    input [0:0] vector ;
  begin
    conv_u2u_1_23 = {{22{1'b0}}, vector};
  end
  endfunction
  function [3:0] conv_u2u_3_4 ;
    input [2:0] vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction
  function [5:0] conv_u2u_5_6 ;
    input [4:0] vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction
  function [8:0] conv_u2u_8_9 ;
    input [7:0] vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction
  function [23:0] conv_u2u_23_24 ;
    input [22:0] vector ;
  begin
    conv_u2u_23_24 = {1'b0, vector};
  end
  endfunction
  function [49:0] conv_u2u_49_50 ;
    input [48:0] vector ;
  begin
    conv_u2u_49_50 = {1'b0, vector};
  end
  endfunction
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul_core
// ------------------------------------------------------------------
module SDP_X_X_mul_core (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_in_rsc_slz, chn_mul_in_rsc_sz, chn_mul_in_rsc_z,
      chn_mul_in_rsc_vz, chn_mul_in_rsc_lz, chn_mul_op_rsc_z, chn_mul_op_rsc_vz,
      chn_mul_op_rsc_lz, cfg_mul_op_rsc_triosy_lz, cfg_mul_bypass_rsc_triosy_lz,
      cfg_mul_prelu_rsc_triosy_lz, cfg_mul_src_rsc_triosy_lz, cfg_nan_to_zero, cfg_precision,
      chn_mul_out_rsc_z, chn_mul_out_rsc_vz, chn_mul_out_rsc_lz, chn_mul_in_rsci_oswt,
      chn_mul_in_rsci_oswt_unreg, chn_mul_op_rsci_oswt, chn_mul_op_rsci_oswt_unreg,
      cfg_mul_op_rsci_d, cfg_mul_bypass_rsci_d, cfg_mul_prelu_rsci_d, cfg_mul_src_rsci_d,
      chn_mul_out_rsci_oswt, chn_mul_out_rsci_oswt_unreg, cfg_mul_op_rsc_triosy_obj_oswt,
      cfg_mul_bypass_rsc_triosy_obj_oswt, cfg_mul_prelu_rsc_triosy_obj_oswt, cfg_mul_src_rsc_triosy_obj_oswt,
      cfg_mul_op_rsc_triosy_obj_oswt_unreg_pff
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output chn_mul_in_rsc_slz;
  input chn_mul_in_rsc_sz;
  input [527:0] chn_mul_in_rsc_z;
  input chn_mul_in_rsc_vz;
  output chn_mul_in_rsc_lz;
  input [255:0] chn_mul_op_rsc_z;
  input chn_mul_op_rsc_vz;
  output chn_mul_op_rsc_lz;
  output cfg_mul_op_rsc_triosy_lz;
  output cfg_mul_bypass_rsc_triosy_lz;
  output cfg_mul_prelu_rsc_triosy_lz;
  output cfg_mul_src_rsc_triosy_lz;
  input cfg_nan_to_zero;
  input [1:0] cfg_precision;
  output [799:0] chn_mul_out_rsc_z;
  input chn_mul_out_rsc_vz;
  output chn_mul_out_rsc_lz;
  input chn_mul_in_rsci_oswt;
  output chn_mul_in_rsci_oswt_unreg;
  input chn_mul_op_rsci_oswt;
  output chn_mul_op_rsci_oswt_unreg;
  input [15:0] cfg_mul_op_rsci_d;
  input cfg_mul_bypass_rsci_d;
  input cfg_mul_prelu_rsci_d;
  input cfg_mul_src_rsci_d;
  input chn_mul_out_rsci_oswt;
  output chn_mul_out_rsci_oswt_unreg;
  input cfg_mul_op_rsc_triosy_obj_oswt;
  input cfg_mul_bypass_rsc_triosy_obj_oswt;
  input cfg_mul_prelu_rsc_triosy_obj_oswt;
  input cfg_mul_src_rsc_triosy_obj_oswt;
  output cfg_mul_op_rsc_triosy_obj_oswt_unreg_pff;
// Interconnect Declarations
  wire core_wen;
  reg chn_mul_in_rsci_iswt0;
  wire chn_mul_in_rsci_bawt;
  wire chn_mul_in_rsci_wen_comp;
  reg chn_mul_in_rsci_ld_core_psct;
  wire [527:0] chn_mul_in_rsci_d_mxwt;
  wire core_wten;
  reg chn_mul_op_rsci_iswt0;
  wire chn_mul_op_rsci_bawt;
  wire chn_mul_op_rsci_wen_comp;
  reg chn_mul_op_rsci_ld_core_psct;
  wire [255:0] chn_mul_op_rsci_d_mxwt;
  reg chn_mul_out_rsci_iswt0;
  wire chn_mul_out_rsci_bawt;
  wire chn_mul_out_rsci_wen_comp;
  wire cfg_mul_op_rsc_triosy_obj_bawt;
  wire cfg_mul_bypass_rsc_triosy_obj_bawt;
  wire cfg_mul_prelu_rsc_triosy_obj_bawt;
  wire cfg_mul_src_rsc_triosy_obj_bawt;
  reg chn_mul_out_rsci_d_799;
  reg chn_mul_out_rsci_d_798;
  reg chn_mul_out_rsci_d_797;
  reg chn_mul_out_rsci_d_796;
  reg chn_mul_out_rsci_d_795;
  reg chn_mul_out_rsci_d_794;
  reg chn_mul_out_rsci_d_793;
  reg chn_mul_out_rsci_d_792;
  reg chn_mul_out_rsci_d_791;
  reg chn_mul_out_rsci_d_790;
  reg chn_mul_out_rsci_d_789;
  reg chn_mul_out_rsci_d_788;
  reg chn_mul_out_rsci_d_787;
  reg chn_mul_out_rsci_d_786;
  reg chn_mul_out_rsci_d_785;
  reg chn_mul_out_rsci_d_784;
  reg [17:0] chn_mul_out_rsci_d_783_766;
  reg [1:0] chn_mul_out_rsci_d_765_764;
  reg [1:0] chn_mul_out_rsci_d_763_762;
  reg [3:0] chn_mul_out_rsci_d_761_758;
  reg [9:0] chn_mul_out_rsci_d_757_748;
  reg [2:0] chn_mul_out_rsci_d_747_745;
  reg [9:0] chn_mul_out_rsci_d_744_735;
  reg [17:0] chn_mul_out_rsci_d_734_717;
  reg [1:0] chn_mul_out_rsci_d_716_715;
  reg [1:0] chn_mul_out_rsci_d_714_713;
  reg [3:0] chn_mul_out_rsci_d_712_709;
  reg [9:0] chn_mul_out_rsci_d_708_699;
  reg [2:0] chn_mul_out_rsci_d_698_696;
  reg [9:0] chn_mul_out_rsci_d_695_686;
  reg [17:0] chn_mul_out_rsci_d_685_668;
  reg [1:0] chn_mul_out_rsci_d_667_666;
  reg [1:0] chn_mul_out_rsci_d_665_664;
  reg [3:0] chn_mul_out_rsci_d_663_660;
  reg [9:0] chn_mul_out_rsci_d_659_650;
  reg [2:0] chn_mul_out_rsci_d_649_647;
  reg [9:0] chn_mul_out_rsci_d_646_637;
  reg [17:0] chn_mul_out_rsci_d_636_619;
  reg [1:0] chn_mul_out_rsci_d_618_617;
  reg [1:0] chn_mul_out_rsci_d_616_615;
  reg [3:0] chn_mul_out_rsci_d_614_611;
  reg [9:0] chn_mul_out_rsci_d_610_601;
  reg [2:0] chn_mul_out_rsci_d_600_598;
  reg [9:0] chn_mul_out_rsci_d_597_588;
  reg [17:0] chn_mul_out_rsci_d_587_570;
  reg [1:0] chn_mul_out_rsci_d_569_568;
  reg [1:0] chn_mul_out_rsci_d_567_566;
  reg [3:0] chn_mul_out_rsci_d_565_562;
  reg [9:0] chn_mul_out_rsci_d_561_552;
  reg [2:0] chn_mul_out_rsci_d_551_549;
  reg [9:0] chn_mul_out_rsci_d_548_539;
  reg [17:0] chn_mul_out_rsci_d_538_521;
  reg [1:0] chn_mul_out_rsci_d_520_519;
  reg [1:0] chn_mul_out_rsci_d_518_517;
  reg [3:0] chn_mul_out_rsci_d_516_513;
  reg [9:0] chn_mul_out_rsci_d_512_503;
  reg [2:0] chn_mul_out_rsci_d_502_500;
  reg [9:0] chn_mul_out_rsci_d_499_490;
  reg [17:0] chn_mul_out_rsci_d_489_472;
  reg [1:0] chn_mul_out_rsci_d_471_470;
  reg [1:0] chn_mul_out_rsci_d_469_468;
  reg [3:0] chn_mul_out_rsci_d_467_464;
  reg [9:0] chn_mul_out_rsci_d_463_454;
  reg [2:0] chn_mul_out_rsci_d_453_451;
  reg [9:0] chn_mul_out_rsci_d_450_441;
  reg [17:0] chn_mul_out_rsci_d_440_423;
  reg [1:0] chn_mul_out_rsci_d_422_421;
  reg [1:0] chn_mul_out_rsci_d_420_419;
  reg [3:0] chn_mul_out_rsci_d_418_415;
  reg [9:0] chn_mul_out_rsci_d_414_405;
  reg [2:0] chn_mul_out_rsci_d_404_402;
  reg [9:0] chn_mul_out_rsci_d_401_392;
  reg [17:0] chn_mul_out_rsci_d_391_374;
  reg [1:0] chn_mul_out_rsci_d_373_372;
  reg [1:0] chn_mul_out_rsci_d_371_370;
  reg [3:0] chn_mul_out_rsci_d_369_366;
  reg [9:0] chn_mul_out_rsci_d_365_356;
  reg [2:0] chn_mul_out_rsci_d_355_353;
  reg [9:0] chn_mul_out_rsci_d_352_343;
  reg [17:0] chn_mul_out_rsci_d_342_325;
  reg [1:0] chn_mul_out_rsci_d_324_323;
  reg [1:0] chn_mul_out_rsci_d_322_321;
  reg [3:0] chn_mul_out_rsci_d_320_317;
  reg [9:0] chn_mul_out_rsci_d_316_307;
  reg [2:0] chn_mul_out_rsci_d_306_304;
  reg [9:0] chn_mul_out_rsci_d_303_294;
  reg [17:0] chn_mul_out_rsci_d_293_276;
  reg [1:0] chn_mul_out_rsci_d_275_274;
  reg [1:0] chn_mul_out_rsci_d_273_272;
  reg [3:0] chn_mul_out_rsci_d_271_268;
  reg [9:0] chn_mul_out_rsci_d_267_258;
  reg [2:0] chn_mul_out_rsci_d_257_255;
  reg [9:0] chn_mul_out_rsci_d_254_245;
  reg [17:0] chn_mul_out_rsci_d_244_227;
  reg [1:0] chn_mul_out_rsci_d_226_225;
  reg [1:0] chn_mul_out_rsci_d_224_223;
  reg [3:0] chn_mul_out_rsci_d_222_219;
  reg [9:0] chn_mul_out_rsci_d_218_209;
  reg [2:0] chn_mul_out_rsci_d_208_206;
  reg [9:0] chn_mul_out_rsci_d_205_196;
  reg [17:0] chn_mul_out_rsci_d_195_178;
  reg [1:0] chn_mul_out_rsci_d_177_176;
  reg [1:0] chn_mul_out_rsci_d_175_174;
  reg [3:0] chn_mul_out_rsci_d_173_170;
  reg [9:0] chn_mul_out_rsci_d_169_160;
  reg [2:0] chn_mul_out_rsci_d_159_157;
  reg [9:0] chn_mul_out_rsci_d_156_147;
  reg [17:0] chn_mul_out_rsci_d_146_129;
  reg [1:0] chn_mul_out_rsci_d_128_127;
  reg [1:0] chn_mul_out_rsci_d_126_125;
  reg [3:0] chn_mul_out_rsci_d_124_121;
  reg [9:0] chn_mul_out_rsci_d_120_111;
  reg [2:0] chn_mul_out_rsci_d_110_108;
  reg [9:0] chn_mul_out_rsci_d_107_98;
  reg [17:0] chn_mul_out_rsci_d_97_80;
  reg [1:0] chn_mul_out_rsci_d_79_78;
  reg [1:0] chn_mul_out_rsci_d_77_76;
  reg [3:0] chn_mul_out_rsci_d_75_72;
  reg [9:0] chn_mul_out_rsci_d_71_62;
  reg [2:0] chn_mul_out_rsci_d_61_59;
  reg [9:0] chn_mul_out_rsci_d_58_49;
  reg [17:0] chn_mul_out_rsci_d_48_31;
  reg [1:0] chn_mul_out_rsci_d_30_29;
  reg [1:0] chn_mul_out_rsci_d_28_27;
  reg [3:0] chn_mul_out_rsci_d_26_23;
  reg [9:0] chn_mul_out_rsci_d_22_13;
  reg [2:0] chn_mul_out_rsci_d_12_10;
  reg [9:0] chn_mul_out_rsci_d_9_0;
  wire [1:0] fsm_output;
  wire IsNaN_5U_10U_nor_15_tmp;
  wire IsNaN_5U_10U_nor_14_tmp;
  wire IsNaN_5U_10U_nor_13_tmp;
  wire IsNaN_5U_10U_nor_12_tmp;
  wire IsNaN_5U_10U_nor_11_tmp;
  wire IsNaN_5U_10U_nor_10_tmp;
  wire IsNaN_5U_10U_nor_9_tmp;
  wire IsNaN_5U_10U_nor_8_tmp;
  wire IsNaN_5U_10U_nor_7_tmp;
  wire IsNaN_5U_10U_nor_6_tmp;
  wire IsNaN_5U_10U_nor_5_tmp;
  wire IsNaN_5U_10U_nor_4_tmp;
  wire IsNaN_5U_10U_nor_3_tmp;
  wire IsNaN_5U_10U_nor_2_tmp;
  wire IsNaN_5U_10U_nor_1_tmp;
  wire IsNaN_5U_10U_nor_tmp;
  wire [4:0] else_mux_47_tmp;
  wire [4:0] else_mux_44_tmp;
  wire [4:0] else_mux_41_tmp;
  wire [4:0] else_mux_38_tmp;
  wire [4:0] else_mux_35_tmp;
  wire [4:0] else_mux_32_tmp;
  wire [4:0] else_mux_29_tmp;
  wire [4:0] else_mux_26_tmp;
  wire [4:0] else_mux_23_tmp;
  wire [4:0] else_mux_20_tmp;
  wire [4:0] else_mux_17_tmp;
  wire [4:0] else_mux_14_tmp;
  wire [4:0] else_mux_11_tmp;
  wire [4:0] else_mux_8_tmp;
  wire [4:0] else_mux_5_tmp;
  wire [4:0] else_mux_2_tmp;
  wire [47:0] mul_loop_mul_16_FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire [47:0] mul_loop_mul_15_FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire [47:0] mul_loop_mul_14_FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire [47:0] mul_loop_mul_13_FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire [47:0] mul_loop_mul_12_FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire [47:0] mul_loop_mul_11_FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire [47:0] mul_loop_mul_10_FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire [47:0] mul_loop_mul_9_FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire [47:0] mul_loop_mul_8_FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire [47:0] mul_loop_mul_7_FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire [47:0] mul_loop_mul_6_FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire [47:0] mul_loop_mul_5_FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire [47:0] mul_loop_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire [47:0] mul_loop_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire [47:0] mul_loop_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire [47:0] mul_loop_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_30_tmp;
  wire IsNaN_5U_23U_nor_15_tmp;
  wire FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_28_tmp;
  wire IsNaN_5U_23U_nor_14_tmp;
  wire IsNaN_5U_23U_nor_13_tmp;
  wire FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_24_tmp;
  wire IsNaN_5U_23U_nor_12_tmp;
  wire IsNaN_5U_23U_nor_11_tmp;
  wire IsNaN_5U_23U_nor_10_tmp;
  wire IsNaN_5U_23U_nor_9_tmp;
  wire FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_16_tmp;
  wire IsNaN_5U_23U_nor_8_tmp;
  wire FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_14_tmp;
  wire IsNaN_5U_23U_nor_7_tmp;
  wire IsNaN_5U_23U_nor_6_tmp;
  wire IsNaN_5U_23U_nor_5_tmp;
  wire FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_8_tmp;
  wire IsNaN_5U_23U_nor_4_tmp;
  wire IsNaN_5U_23U_nor_3_tmp;
  wire FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_4_tmp;
  wire IsNaN_5U_23U_nor_2_tmp;
  wire FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_2_tmp;
  wire IsNaN_5U_23U_nor_1_tmp;
  wire FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_tmp;
  wire IsNaN_5U_23U_nor_tmp;
  wire and_dcpl_2;
  wire and_dcpl_3;
  wire and_dcpl_4;
  wire and_dcpl_5;
  wire or_dcpl_4;
  wire and_dcpl_7;
  wire or_tmp_4;
  wire or_tmp_5;
  wire mux_tmp_1;
  wire nand_tmp_1;
  wire or_tmp_8;
  wire nand_tmp_2;
  wire not_tmp_8;
  wire mux_tmp_2;
  wire or_tmp_9;
  wire or_tmp_10;
  wire mux_tmp_5;
  wire mux_tmp_8;
  wire or_tmp_14;
  wire or_tmp_15;
  wire mux_tmp_14;
  wire mux_tmp_18;
  wire or_tmp_21;
  wire or_tmp_22;
  wire mux_tmp_24;
  wire mux_tmp_28;
  wire mux_tmp_33;
  wire or_tmp_29;
  wire or_tmp_30;
  wire mux_tmp_34;
  wire mux_tmp_35;
  wire mux_tmp_36;
  wire mux_tmp_38;
  wire or_tmp_37;
  wire or_tmp_38;
  wire mux_tmp_44;
  wire mux_tmp_48;
  wire or_tmp_44;
  wire or_tmp_45;
  wire mux_tmp_53;
  wire mux_tmp_55;
  wire or_tmp_50;
  wire or_tmp_51;
  wire mux_tmp_60;
  wire mux_tmp_62;
  wire or_tmp_56;
  wire or_tmp_57;
  wire mux_tmp_68;
  wire mux_tmp_72;
  wire or_tmp_63;
  wire or_tmp_64;
  wire mux_tmp_78;
  wire mux_tmp_82;
  wire or_tmp_70;
  wire or_tmp_71;
  wire mux_tmp_87;
  wire mux_tmp_89;
  wire or_tmp_76;
  wire or_tmp_77;
  wire mux_tmp_94;
  wire mux_tmp_96;
  wire or_tmp_82;
  wire or_tmp_83;
  wire mux_tmp_101;
  wire mux_tmp_103;
  wire or_tmp_88;
  wire or_tmp_89;
  wire mux_tmp_109;
  wire mux_tmp_113;
  wire or_tmp_95;
  wire or_tmp_96;
  wire mux_tmp_118;
  wire mux_tmp_120;
  wire or_tmp_101;
  wire or_tmp_102;
  wire mux_tmp_126;
  wire mux_tmp_130;
  wire or_tmp_108;
  wire or_tmp_109;
  wire mux_tmp_136;
  wire mux_tmp_140;
  wire or_tmp_115;
  wire mux_tmp_148;
  wire not_tmp_30;
  wire or_tmp_122;
  wire or_tmp_123;
  wire or_tmp_128;
  wire or_tmp_129;
  wire or_tmp_134;
  wire or_tmp_135;
  wire or_tmp_139;
  wire or_tmp_141;
  wire or_tmp_142;
  wire or_tmp_147;
  wire or_tmp_148;
  wire or_tmp_151;
  wire or_tmp_152;
  wire or_tmp_155;
  wire or_tmp_156;
  wire or_tmp_161;
  wire or_tmp_162;
  wire or_tmp_167;
  wire or_tmp_168;
  wire or_tmp_171;
  wire or_tmp_172;
  wire or_tmp_175;
  wire or_tmp_176;
  wire or_tmp_179;
  wire or_tmp_180;
  wire or_tmp_185;
  wire or_tmp_186;
  wire or_tmp_189;
  wire or_tmp_190;
  wire or_tmp_195;
  wire or_tmp_196;
  wire or_tmp_201;
  wire or_tmp_202;
  wire or_tmp_204;
  wire or_tmp_213;
  wire or_tmp_228;
  wire or_tmp_236;
  wire or_tmp_248;
  wire or_tmp_256;
  wire or_tmp_264;
  wire or_tmp_279;
  wire or_tmp_287;
  wire or_tmp_302;
  wire or_tmp_310;
  wire or_tmp_321;
  wire or_tmp_322;
  wire or_tmp_331;
  wire or_tmp_339;
  wire or_tmp_354;
  wire or_tmp_362;
  wire or_tmp_377;
  wire or_tmp_385;
  wire or_tmp_397;
  wire or_tmp_405;
  wire or_tmp_413;
  wire or_tmp_424;
  wire or_tmp_425;
  wire or_tmp_434;
  wire or_tmp_442;
  wire or_tmp_453;
  wire or_tmp_454;
  wire or_tmp_460;
  wire or_tmp_463;
  wire or_tmp_471;
  wire or_tmp_486;
  wire or_tmp_494;
  wire or_tmp_509;
  wire or_tmp_517;
  wire or_tmp_532;
  wire or_tmp_540;
  wire or_tmp_555;
  wire or_tmp_563;
  wire or_tmp_578;
  wire or_tmp_586;
  wire or_tmp_597;
  wire or_tmp_598;
  wire or_tmp_606;
  wire or_tmp_608;
  wire mux_tmp_399;
  wire mux_tmp_402;
  wire mux_tmp_403;
  wire mux_tmp_406;
  wire mux_tmp_409;
  wire mux_tmp_412;
  wire mux_tmp_415;
  wire mux_tmp_418;
  wire mux_tmp_421;
  wire mux_tmp_424;
  wire mux_tmp_427;
  wire mux_tmp_430;
  wire mux_tmp_433;
  wire mux_tmp_436;
  wire mux_tmp_439;
  wire mux_tmp_442;
  wire mux_tmp_445;
  wire mux_tmp_448;
  wire mux_tmp_451;
  wire mux_tmp_454;
  wire mux_tmp_457;
  wire mux_tmp_460;
  wire mux_tmp_463;
  wire mux_tmp_466;
  wire mux_tmp_469;
  wire mux_tmp_472;
  wire mux_tmp_475;
  wire mux_tmp_478;
  wire mux_tmp_481;
  wire mux_tmp_484;
  wire mux_tmp_487;
  wire mux_tmp_490;
  wire mux_tmp_493;
  wire or_tmp_893;
  wire or_tmp_898;
  wire or_tmp_932;
  wire or_tmp_958;
  wire or_tmp_975;
  wire or_tmp_980;
  wire or_tmp_1012;
  wire or_tmp_1038;
  wire or_tmp_1055;
  wire or_tmp_1060;
  wire or_tmp_1088;
  wire or_tmp_1094;
  wire or_tmp_1120;
  wire or_tmp_1137;
  wire or_tmp_1142;
  wire or_tmp_1177;
  wire or_tmp_1203;
  wire or_tmp_1220;
  wire or_tmp_1225;
  wire or_tmp_1257;
  wire or_tmp_1283;
  wire or_tmp_1300;
  wire or_tmp_1305;
  wire or_tmp_1333;
  wire or_tmp_1339;
  wire or_tmp_1365;
  wire or_tmp_1382;
  wire or_tmp_1387;
  wire or_tmp_1415;
  wire or_tmp_1421;
  wire or_tmp_1447;
  wire or_tmp_1464;
  wire or_tmp_1469;
  wire or_tmp_1501;
  wire or_tmp_1527;
  wire or_tmp_1544;
  wire or_tmp_1549;
  wire or_tmp_1581;
  wire or_tmp_1607;
  wire or_tmp_1624;
  wire or_tmp_1629;
  wire or_tmp_1661;
  wire or_tmp_1687;
  wire or_tmp_1703;
  wire or_tmp_1709;
  wire or_tmp_1736;
  wire mux_tmp_748;
  wire or_tmp_1744;
  wire or_tmp_1765;
  wire or_tmp_1782;
  wire or_tmp_1786;
  wire or_tmp_1822;
  wire or_tmp_1848;
  wire or_tmp_1865;
  wire or_tmp_1869;
  wire or_tmp_1905;
  wire or_tmp_1931;
  wire or_tmp_1947;
  wire or_tmp_1957;
  wire or_tmp_1985;
  wire or_tmp_1991;
  wire or_tmp_2015;
  wire or_tmp_2032;
  wire or_tmp_2036;
  wire or_tmp_2065;
  wire or_tmp_2071;
  wire or_tmp_2097;
  wire or_tmp_2114;
  wire or_tmp_2118;
  wire or_tmp_2151;
  wire or_tmp_2177;
  wire or_tmp_2227;
  wire or_tmp_2254;
  wire and_tmp_72;
  wire or_tmp_2298;
  wire and_tmp_76;
  wire or_tmp_2310;
  wire or_tmp_2319;
  wire or_tmp_2358;
  wire or_tmp_2366;
  wire or_tmp_2376;
  wire or_tmp_2384;
  wire or_tmp_2392;
  wire or_tmp_2400;
  wire or_tmp_2408;
  wire or_tmp_2414;
  wire or_tmp_2424;
  wire or_tmp_2432;
  wire or_tmp_2440;
  wire or_tmp_2448;
  wire or_tmp_2456;
  wire or_tmp_2464;
  wire or_tmp_2472;
  wire or_tmp_2480;
  wire or_tmp_2490;
  wire or_tmp_2492;
  wire and_tmp_86;
  wire or_tmp_2503;
  wire or_tmp_2521;
  wire or_tmp_2523;
  wire and_tmp_90;
  wire or_tmp_2534;
  wire or_tmp_2538;
  wire or_tmp_2544;
  wire or_tmp_2546;
  wire and_tmp_95;
  wire or_tmp_2557;
  wire or_tmp_2588;
  wire or_tmp_2590;
  wire and_tmp_99;
  wire or_tmp_2601;
  wire or_tmp_2604;
  wire or_tmp_2635;
  wire or_tmp_2637;
  wire and_tmp_104;
  wire or_tmp_2648;
  wire or_tmp_2652;
  wire or_tmp_2658;
  wire or_tmp_2660;
  wire and_tmp_109;
  wire or_tmp_2671;
  wire or_tmp_2674;
  wire or_tmp_2711;
  wire or_tmp_2713;
  wire and_tmp_114;
  wire or_tmp_2724;
  wire or_tmp_2728;
  wire or_tmp_2747;
  wire or_tmp_2749;
  wire and_tmp_119;
  wire or_tmp_2760;
  wire or_tmp_2778;
  wire or_tmp_2780;
  wire and_tmp_123;
  wire or_tmp_2791;
  wire or_tmp_2795;
  wire mux_tmp_1422;
  wire not_tmp_845;
  wire mux_tmp_1427;
  wire mux_tmp_1430;
  wire or_tmp_2894;
  wire or_tmp_2905;
  wire or_tmp_2916;
  wire or_tmp_2927;
  wire or_tmp_2938;
  wire or_tmp_2949;
  wire or_tmp_2960;
  wire or_tmp_2971;
  wire or_tmp_2982;
  wire or_tmp_2993;
  wire or_tmp_3004;
  wire or_tmp_3015;
  wire or_tmp_3026;
  wire or_tmp_3037;
  wire or_tmp_3048;
  wire mux_tmp_1504;
  wire mux_tmp_1507;
  wire mux_tmp_1510;
  wire mux_tmp_1513;
  wire mux_tmp_1516;
  wire mux_tmp_1535;
  wire mux_tmp_1538;
  wire and_dcpl_47;
  wire and_dcpl_50;
  wire and_dcpl_52;
  wire or_dcpl_27;
  wire and_dcpl_53;
  wire and_dcpl_56;
  wire and_dcpl_58;
  wire and_dcpl_59;
  wire or_dcpl_31;
  wire and_dcpl_67;
  wire nor_tmp_568;
  wire and_dcpl_72;
  wire and_dcpl_75;
  wire and_dcpl_85;
  wire and_dcpl_87;
  wire or_dcpl_46;
  wire and_dcpl_91;
  wire and_dcpl_95;
  wire and_dcpl_100;
  wire and_dcpl_102;
  wire and_dcpl_104;
  wire and_dcpl_108;
  wire and_dcpl_112;
  wire and_dcpl_116;
  wire and_dcpl_120;
  wire and_dcpl_124;
  wire and_dcpl_128;
  wire and_dcpl_132;
  wire and_dcpl_136;
  wire and_dcpl_140;
  wire and_dcpl_144;
  wire and_dcpl_148;
  wire and_dcpl_152;
  wire and_dcpl_156;
  wire and_dcpl_160;
  wire and_dcpl_164;
  wire and_dcpl_172;
  wire and_dcpl_177;
  wire and_dcpl_182;
  wire and_dcpl_187;
  wire and_dcpl_192;
  wire and_dcpl_197;
  wire and_dcpl_202;
  wire and_dcpl_207;
  wire and_dcpl_212;
  wire and_dcpl_217;
  wire and_dcpl_222;
  wire and_dcpl_227;
  wire and_dcpl_232;
  wire and_dcpl_237;
  wire and_dcpl_242;
  wire and_dcpl_247;
  wire or_dcpl_87;
  wire or_dcpl_92;
  wire or_dcpl_95;
  wire or_dcpl_96;
  wire or_dcpl_100;
  wire or_dcpl_103;
  wire or_dcpl_107;
  wire or_dcpl_110;
  wire or_dcpl_115;
  wire or_dcpl_118;
  wire or_dcpl_122;
  wire or_dcpl_125;
  wire or_dcpl_129;
  wire or_dcpl_132;
  wire or_dcpl_136;
  wire or_dcpl_139;
  wire or_dcpl_143;
  wire or_dcpl_146;
  wire or_dcpl_150;
  wire or_dcpl_153;
  wire or_dcpl_157;
  wire or_dcpl_160;
  wire or_dcpl_165;
  wire or_dcpl_168;
  wire or_dcpl_173;
  wire or_dcpl_176;
  wire or_dcpl_181;
  wire or_dcpl_184;
  wire or_dcpl_188;
  wire or_dcpl_191;
  wire or_dcpl_195;
  wire or_dcpl_198;
  wire or_dcpl_202;
  wire or_dcpl_205;
  wire and_dcpl_254;
  wire and_dcpl_255;
  wire and_dcpl_258;
  wire and_dcpl_259;
  wire or_dcpl_206;
  wire and_dcpl_262;
  wire and_dcpl_263;
  wire or_dcpl_212;
  wire and_dcpl_266;
  wire or_dcpl_216;
  wire or_dcpl_217;
  wire and_dcpl_269;
  wire and_dcpl_270;
  wire and_dcpl_273;
  wire and_dcpl_274;
  wire or_dcpl_218;
  wire and_dcpl_277;
  wire and_dcpl_278;
  wire or_dcpl_224;
  wire and_dcpl_281;
  wire or_dcpl_227;
  wire and_dcpl_284;
  wire and_dcpl_285;
  wire and_dcpl_288;
  wire and_dcpl_289;
  wire or_dcpl_228;
  wire and_dcpl_292;
  wire and_dcpl_293;
  wire or_dcpl_234;
  wire and_dcpl_296;
  wire or_dcpl_237;
  wire and_dcpl_299;
  wire and_dcpl_300;
  wire and_dcpl_303;
  wire and_dcpl_304;
  wire or_dcpl_238;
  wire and_dcpl_307;
  wire and_dcpl_308;
  wire or_dcpl_244;
  wire and_dcpl_311;
  wire or_dcpl_247;
  wire and_dcpl_314;
  wire and_dcpl_315;
  wire and_dcpl_318;
  wire and_dcpl_319;
  wire or_dcpl_248;
  wire and_dcpl_322;
  wire and_dcpl_323;
  wire or_dcpl_254;
  wire and_dcpl_326;
  wire or_dcpl_257;
  wire and_dcpl_329;
  wire and_dcpl_330;
  wire and_dcpl_333;
  wire and_dcpl_334;
  wire or_dcpl_258;
  wire and_dcpl_337;
  wire and_dcpl_338;
  wire or_dcpl_264;
  wire and_dcpl_341;
  wire or_dcpl_267;
  wire and_dcpl_344;
  wire and_dcpl_345;
  wire or_dcpl_268;
  wire and_dcpl_349;
  wire and_dcpl_352;
  wire and_dcpl_353;
  wire or_dcpl_274;
  wire and_dcpl_356;
  wire or_dcpl_277;
  wire and_dcpl_359;
  wire and_dcpl_360;
  wire or_dcpl_278;
  wire and_dcpl_364;
  wire and_dcpl_367;
  wire and_dcpl_368;
  wire or_dcpl_284;
  wire and_dcpl_371;
  wire or_dcpl_287;
  wire and_dcpl_374;
  wire and_dcpl_375;
  wire or_dcpl_288;
  wire and_dcpl_379;
  wire and_dcpl_382;
  wire and_dcpl_383;
  wire or_dcpl_294;
  wire and_dcpl_386;
  wire or_dcpl_297;
  wire and_dcpl_389;
  wire and_dcpl_390;
  wire and_dcpl_393;
  wire and_dcpl_394;
  wire or_dcpl_298;
  wire and_dcpl_397;
  wire and_dcpl_398;
  wire or_dcpl_304;
  wire and_dcpl_401;
  wire or_dcpl_307;
  wire and_dcpl_404;
  wire and_dcpl_405;
  wire and_dcpl_408;
  wire and_dcpl_409;
  wire or_dcpl_308;
  wire and_dcpl_412;
  wire and_dcpl_413;
  wire or_dcpl_314;
  wire and_dcpl_416;
  wire or_dcpl_317;
  wire and_dcpl_419;
  wire and_dcpl_420;
  wire and_dcpl_423;
  wire and_dcpl_424;
  wire or_dcpl_318;
  wire and_dcpl_427;
  wire and_dcpl_428;
  wire or_dcpl_324;
  wire and_dcpl_431;
  wire or_dcpl_327;
  wire and_dcpl_434;
  wire and_dcpl_435;
  wire and_dcpl_438;
  wire and_dcpl_439;
  wire or_dcpl_328;
  wire and_dcpl_442;
  wire and_dcpl_443;
  wire or_dcpl_334;
  wire and_dcpl_446;
  wire or_dcpl_337;
  wire and_dcpl_449;
  wire and_dcpl_450;
  wire and_dcpl_453;
  wire and_dcpl_454;
  wire or_dcpl_338;
  wire and_dcpl_457;
  wire and_dcpl_458;
  wire or_dcpl_344;
  wire and_dcpl_461;
  wire or_dcpl_347;
  wire and_dcpl_464;
  wire and_dcpl_465;
  wire and_dcpl_468;
  wire and_dcpl_469;
  wire or_dcpl_348;
  wire and_dcpl_472;
  wire and_dcpl_473;
  wire or_dcpl_354;
  wire and_dcpl_476;
  wire or_dcpl_357;
  wire and_dcpl_479;
  wire and_dcpl_480;
  wire and_dcpl_483;
  wire and_dcpl_484;
  wire or_dcpl_358;
  wire and_dcpl_487;
  wire and_dcpl_488;
  wire or_dcpl_364;
  wire and_dcpl_491;
  wire or_dcpl_367;
  wire and_dcpl_492;
  wire or_dcpl_369;
  wire or_dcpl_373;
  wire or_dcpl_382;
  wire or_dcpl_385;
  wire and_dcpl_494;
  wire and_dcpl_497;
  wire and_dcpl_500;
  wire and_dcpl_503;
  wire and_dcpl_506;
  wire and_dcpl_509;
  wire and_dcpl_512;
  wire and_dcpl_515;
  wire and_dcpl_518;
  wire and_dcpl_521;
  wire and_dcpl_524;
  wire and_dcpl_527;
  wire and_dcpl_530;
  wire and_dcpl_533;
  wire and_dcpl_536;
  wire and_dcpl_539;
  wire and_dcpl_542;
  wire and_dcpl_546;
  wire and_dcpl_555;
  wire and_dcpl_564;
  wire and_dcpl_573;
  wire and_dcpl_582;
  wire and_dcpl_591;
  wire and_dcpl_600;
  wire and_dcpl_609;
  wire and_dcpl_618;
  wire and_dcpl_627;
  wire and_dcpl_636;
  wire and_dcpl_645;
  wire and_dcpl_654;
  wire and_dcpl_663;
  wire and_dcpl_672;
  wire and_dcpl_681;
  wire and_dcpl_770;
  wire and_dcpl_873;
  wire and_dcpl_879;
  wire and_dcpl_891;
  wire and_dcpl_903;
  wire and_dcpl_915;
  wire and_dcpl_927;
  wire and_dcpl_939;
  wire and_dcpl_951;
  wire and_dcpl_963;
  wire and_dcpl_975;
  wire and_dcpl_987;
  wire and_dcpl_999;
  wire and_dcpl_1011;
  wire and_dcpl_1023;
  wire and_dcpl_1035;
  wire and_dcpl_1047;
  wire and_dcpl_1059;
  wire or_dcpl_665;
  wire or_tmp_3606;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3;
  reg IsZero_8U_23U_land_1_lpi_1_dfm;
  reg IsZero_8U_23U_1_land_1_lpi_1_dfm;
  reg mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_1_sva;
  reg [7:0] FpMul_8U_23U_p_expo_1_sva_1;
  reg FpMantRNE_48U_24U_else_carry_1_sva;
  reg mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3;
  reg IsZero_8U_23U_land_2_lpi_1_dfm;
  reg IsZero_8U_23U_1_land_2_lpi_1_dfm;
  reg mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_2_sva;
  reg [7:0] FpMul_8U_23U_p_expo_2_sva_1;
  reg FpMantRNE_48U_24U_else_carry_2_sva;
  reg mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3;
  reg IsZero_8U_23U_land_3_lpi_1_dfm;
  reg IsZero_8U_23U_1_land_3_lpi_1_dfm;
  reg mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_3_sva;
  reg [7:0] FpMul_8U_23U_p_expo_3_sva_1;
  reg FpMantRNE_48U_24U_else_carry_3_sva;
  reg mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3;
  reg IsZero_8U_23U_land_4_lpi_1_dfm;
  reg IsZero_8U_23U_1_land_4_lpi_1_dfm;
  reg mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_4_sva;
  reg [7:0] FpMul_8U_23U_p_expo_4_sva_1;
  reg FpMantRNE_48U_24U_else_carry_4_sva;
  reg mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs;
  reg IsNaN_8U_23U_land_4_lpi_1_dfm;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3;
  reg IsZero_8U_23U_land_5_lpi_1_dfm;
  reg IsZero_8U_23U_1_land_5_lpi_1_dfm;
  reg mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_5_sva;
  reg [7:0] FpMul_8U_23U_p_expo_5_sva_1;
  reg FpMantRNE_48U_24U_else_carry_5_sva;
  reg mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs;
  reg IsNaN_8U_23U_land_5_lpi_1_dfm;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3;
  reg IsZero_8U_23U_land_6_lpi_1_dfm;
  reg IsZero_8U_23U_1_land_6_lpi_1_dfm;
  reg mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_6_sva;
  reg [7:0] FpMul_8U_23U_p_expo_6_sva_1;
  reg FpMantRNE_48U_24U_else_carry_6_sva;
  reg mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs;
  reg IsNaN_8U_23U_land_6_lpi_1_dfm;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3;
  reg IsZero_8U_23U_land_7_lpi_1_dfm;
  reg IsZero_8U_23U_1_land_7_lpi_1_dfm;
  reg mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_7_sva;
  reg [7:0] FpMul_8U_23U_p_expo_7_sva_1;
  reg FpMantRNE_48U_24U_else_carry_7_sva;
  reg mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs;
  reg IsNaN_8U_23U_land_7_lpi_1_dfm;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3;
  reg IsZero_8U_23U_land_8_lpi_1_dfm;
  reg IsZero_8U_23U_1_land_8_lpi_1_dfm;
  reg mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_8_sva;
  reg [7:0] FpMul_8U_23U_p_expo_8_sva_1;
  reg FpMantRNE_48U_24U_else_carry_8_sva;
  reg mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs;
  reg IsNaN_8U_23U_land_8_lpi_1_dfm;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3;
  reg IsZero_8U_23U_land_9_lpi_1_dfm;
  reg IsZero_8U_23U_1_land_9_lpi_1_dfm;
  reg mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_9_sva;
  reg [7:0] FpMul_8U_23U_p_expo_9_sva_1;
  reg FpMantRNE_48U_24U_else_carry_9_sva;
  reg mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs;
  reg IsNaN_8U_23U_land_9_lpi_1_dfm;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3;
  reg IsZero_8U_23U_land_10_lpi_1_dfm;
  reg IsZero_8U_23U_1_land_10_lpi_1_dfm;
  reg mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_10_sva;
  reg [7:0] FpMul_8U_23U_p_expo_10_sva_1;
  reg FpMantRNE_48U_24U_else_carry_10_sva;
  reg mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs;
  reg IsNaN_8U_23U_land_10_lpi_1_dfm;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3;
  reg IsZero_8U_23U_land_11_lpi_1_dfm;
  reg IsZero_8U_23U_1_land_11_lpi_1_dfm;
  reg mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_11_sva;
  reg [7:0] FpMul_8U_23U_p_expo_11_sva_1;
  reg FpMantRNE_48U_24U_else_carry_11_sva;
  reg mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs;
  reg IsNaN_8U_23U_land_11_lpi_1_dfm;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3;
  reg IsZero_8U_23U_land_12_lpi_1_dfm;
  reg IsZero_8U_23U_1_land_12_lpi_1_dfm;
  reg mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_12_sva;
  reg [7:0] FpMul_8U_23U_p_expo_12_sva_1;
  reg FpMantRNE_48U_24U_else_carry_12_sva;
  reg mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs;
  reg IsNaN_8U_23U_land_12_lpi_1_dfm;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3;
  reg IsZero_8U_23U_land_13_lpi_1_dfm;
  reg IsZero_8U_23U_1_land_13_lpi_1_dfm;
  reg mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_13_sva;
  reg [7:0] FpMul_8U_23U_p_expo_13_sva_1;
  reg FpMantRNE_48U_24U_else_carry_13_sva;
  reg mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs;
  reg IsNaN_8U_23U_land_13_lpi_1_dfm;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3;
  reg IsZero_8U_23U_land_14_lpi_1_dfm;
  reg IsZero_8U_23U_1_land_14_lpi_1_dfm;
  reg mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_14_sva;
  reg [7:0] FpMul_8U_23U_p_expo_14_sva_1;
  reg FpMantRNE_48U_24U_else_carry_14_sva;
  reg mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs;
  reg IsNaN_8U_23U_land_14_lpi_1_dfm;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3;
  reg IsZero_8U_23U_land_15_lpi_1_dfm;
  reg IsZero_8U_23U_1_land_15_lpi_1_dfm;
  reg mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_15_sva;
  reg [7:0] FpMul_8U_23U_p_expo_15_sva_1;
  reg FpMantRNE_48U_24U_else_carry_15_sva;
  reg mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs;
  reg IsNaN_8U_23U_land_15_lpi_1_dfm;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3;
  reg IsZero_8U_23U_land_lpi_1_dfm;
  reg IsZero_8U_23U_1_land_lpi_1_dfm;
  reg mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_sva;
  reg [7:0] FpMul_8U_23U_p_expo_sva_1;
  reg FpMantRNE_48U_24U_else_carry_sva;
  reg mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs;
  reg IsNaN_8U_23U_land_lpi_1_dfm;
  reg main_stage_v_1;
  reg main_stage_v_2;
  reg main_stage_v_3;
  reg main_stage_v_4;
  reg mul_loop_mul_if_land_lpi_1_dfm_7;
  reg mul_loop_mul_if_land_lpi_1_dfm_8;
  reg mul_loop_mul_if_land_lpi_1_dfm_9;
  reg mul_loop_mul_if_land_lpi_1_dfm_10;
  reg mul_loop_mul_if_land_15_lpi_1_dfm_7;
  reg mul_loop_mul_if_land_15_lpi_1_dfm_8;
  reg mul_loop_mul_if_land_15_lpi_1_dfm_9;
  reg mul_loop_mul_if_land_15_lpi_1_dfm_10;
  reg mul_loop_mul_if_land_14_lpi_1_dfm_7;
  reg mul_loop_mul_if_land_14_lpi_1_dfm_8;
  reg mul_loop_mul_if_land_14_lpi_1_dfm_9;
  reg mul_loop_mul_if_land_14_lpi_1_dfm_10;
  reg mul_loop_mul_if_land_13_lpi_1_dfm_7;
  reg mul_loop_mul_if_land_13_lpi_1_dfm_8;
  reg mul_loop_mul_if_land_13_lpi_1_dfm_9;
  reg mul_loop_mul_if_land_13_lpi_1_dfm_10;
  reg mul_loop_mul_if_land_12_lpi_1_dfm_7;
  reg mul_loop_mul_if_land_12_lpi_1_dfm_8;
  reg mul_loop_mul_if_land_12_lpi_1_dfm_9;
  reg mul_loop_mul_if_land_12_lpi_1_dfm_10;
  reg mul_loop_mul_if_land_11_lpi_1_dfm_7;
  reg mul_loop_mul_if_land_11_lpi_1_dfm_8;
  reg mul_loop_mul_if_land_11_lpi_1_dfm_9;
  reg mul_loop_mul_if_land_11_lpi_1_dfm_10;
  reg mul_loop_mul_if_land_10_lpi_1_dfm_7;
  reg mul_loop_mul_if_land_10_lpi_1_dfm_8;
  reg mul_loop_mul_if_land_10_lpi_1_dfm_9;
  reg mul_loop_mul_if_land_10_lpi_1_dfm_10;
  reg mul_loop_mul_if_land_9_lpi_1_dfm_7;
  reg mul_loop_mul_if_land_9_lpi_1_dfm_8;
  reg mul_loop_mul_if_land_9_lpi_1_dfm_9;
  reg mul_loop_mul_if_land_9_lpi_1_dfm_10;
  reg mul_loop_mul_if_land_8_lpi_1_dfm_7;
  reg mul_loop_mul_if_land_8_lpi_1_dfm_8;
  reg mul_loop_mul_if_land_8_lpi_1_dfm_9;
  reg mul_loop_mul_if_land_8_lpi_1_dfm_10;
  reg mul_loop_mul_if_land_7_lpi_1_dfm_7;
  reg mul_loop_mul_if_land_7_lpi_1_dfm_8;
  reg mul_loop_mul_if_land_7_lpi_1_dfm_9;
  reg mul_loop_mul_if_land_7_lpi_1_dfm_10;
  reg mul_loop_mul_if_land_6_lpi_1_dfm_7;
  reg mul_loop_mul_if_land_6_lpi_1_dfm_8;
  reg mul_loop_mul_if_land_6_lpi_1_dfm_9;
  reg mul_loop_mul_if_land_6_lpi_1_dfm_10;
  reg mul_loop_mul_if_land_5_lpi_1_dfm_7;
  reg mul_loop_mul_if_land_5_lpi_1_dfm_8;
  reg mul_loop_mul_if_land_5_lpi_1_dfm_9;
  reg mul_loop_mul_if_land_5_lpi_1_dfm_10;
  reg mul_loop_mul_if_land_4_lpi_1_dfm_7;
  reg mul_loop_mul_if_land_4_lpi_1_dfm_8;
  reg mul_loop_mul_if_land_4_lpi_1_dfm_9;
  reg mul_loop_mul_if_land_4_lpi_1_dfm_10;
  reg mul_loop_mul_if_land_3_lpi_1_dfm_7;
  reg mul_loop_mul_if_land_3_lpi_1_dfm_8;
  reg mul_loop_mul_if_land_3_lpi_1_dfm_9;
  reg mul_loop_mul_if_land_3_lpi_1_dfm_10;
  reg mul_loop_mul_if_land_2_lpi_1_dfm_7;
  reg mul_loop_mul_if_land_2_lpi_1_dfm_8;
  reg mul_loop_mul_if_land_2_lpi_1_dfm_9;
  reg mul_loop_mul_if_land_2_lpi_1_dfm_10;
  reg mul_loop_mul_if_land_1_lpi_1_dfm_7;
  reg mul_loop_mul_if_land_1_lpi_1_dfm_8;
  reg mul_loop_mul_if_land_1_lpi_1_dfm_9;
  reg mul_loop_mul_if_land_1_lpi_1_dfm_10;
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_9;
  reg mul_nan_to_zero_op_sign_lpi_1_dfm_4;
  reg IsNaN_8U_23U_1_land_15_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_15_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_15_lpi_1_dfm_9;
  reg mul_nan_to_zero_op_sign_15_lpi_1_dfm_4;
  reg IsNaN_8U_23U_1_land_14_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_14_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_14_lpi_1_dfm_9;
  reg mul_nan_to_zero_op_sign_14_lpi_1_dfm_4;
  reg IsNaN_8U_23U_1_land_13_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_13_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_13_lpi_1_dfm_9;
  reg mul_nan_to_zero_op_sign_13_lpi_1_dfm_4;
  reg IsNaN_8U_23U_1_land_12_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_12_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_12_lpi_1_dfm_9;
  reg mul_nan_to_zero_op_sign_12_lpi_1_dfm_4;
  reg IsNaN_8U_23U_1_land_11_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_11_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_11_lpi_1_dfm_9;
  reg mul_nan_to_zero_op_sign_11_lpi_1_dfm_4;
  reg IsNaN_8U_23U_1_land_10_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_10_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_10_lpi_1_dfm_9;
  reg mul_nan_to_zero_op_sign_10_lpi_1_dfm_4;
  reg IsNaN_8U_23U_1_land_9_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_9_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_9_lpi_1_dfm_9;
  reg mul_nan_to_zero_op_sign_9_lpi_1_dfm_4;
  reg IsNaN_8U_23U_1_land_8_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_8_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_8_lpi_1_dfm_9;
  reg mul_nan_to_zero_op_sign_8_lpi_1_dfm_4;
  reg IsNaN_8U_23U_1_land_7_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_7_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_7_lpi_1_dfm_9;
  reg mul_nan_to_zero_op_sign_7_lpi_1_dfm_4;
  reg IsNaN_8U_23U_1_land_6_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_6_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_6_lpi_1_dfm_9;
  reg mul_nan_to_zero_op_sign_6_lpi_1_dfm_4;
  reg IsNaN_8U_23U_1_land_5_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_5_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_5_lpi_1_dfm_9;
  reg mul_nan_to_zero_op_sign_5_lpi_1_dfm_4;
  reg IsNaN_8U_23U_1_land_4_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_4_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_4_lpi_1_dfm_9;
  reg mul_nan_to_zero_op_sign_4_lpi_1_dfm_4;
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_9;
  reg mul_nan_to_zero_op_sign_3_lpi_1_dfm_4;
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_9;
  reg mul_nan_to_zero_op_sign_2_lpi_1_dfm_4;
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_9;
  reg mul_nan_to_zero_op_sign_1_lpi_1_dfm_4;
  reg [48:0] MulOut_data_15_sva_8;
  reg [48:0] MulOut_data_15_sva_9;
  reg [48:0] MulOut_data_15_sva_10;
  reg mul_loop_mul_else_land_lpi_1_dfm_7;
  reg mul_loop_mul_else_land_lpi_1_dfm_8;
  reg mul_loop_mul_else_land_lpi_1_dfm_9;
  reg mul_loop_mul_else_land_lpi_1_dfm_10;
  reg [48:0] MulOut_data_14_sva_8;
  reg [48:0] MulOut_data_14_sva_9;
  reg [48:0] MulOut_data_14_sva_10;
  reg mul_loop_mul_else_land_15_lpi_1_dfm_7;
  reg mul_loop_mul_else_land_15_lpi_1_dfm_8;
  reg mul_loop_mul_else_land_15_lpi_1_dfm_9;
  reg mul_loop_mul_else_land_15_lpi_1_dfm_10;
  reg [48:0] MulOut_data_13_sva_8;
  reg [48:0] MulOut_data_13_sva_9;
  reg [48:0] MulOut_data_13_sva_10;
  reg mul_loop_mul_else_land_14_lpi_1_dfm_7;
  reg mul_loop_mul_else_land_14_lpi_1_dfm_8;
  reg mul_loop_mul_else_land_14_lpi_1_dfm_9;
  reg mul_loop_mul_else_land_14_lpi_1_dfm_10;
  reg [48:0] MulOut_data_12_sva_8;
  reg [48:0] MulOut_data_12_sva_9;
  reg [48:0] MulOut_data_12_sva_10;
  reg mul_loop_mul_else_land_13_lpi_1_dfm_7;
  reg mul_loop_mul_else_land_13_lpi_1_dfm_8;
  reg mul_loop_mul_else_land_13_lpi_1_dfm_9;
  reg mul_loop_mul_else_land_13_lpi_1_dfm_10;
  reg [48:0] MulOut_data_11_sva_8;
  reg [48:0] MulOut_data_11_sva_9;
  reg [48:0] MulOut_data_11_sva_10;
  reg mul_loop_mul_else_land_12_lpi_1_dfm_7;
  reg mul_loop_mul_else_land_12_lpi_1_dfm_8;
  reg mul_loop_mul_else_land_12_lpi_1_dfm_9;
  reg mul_loop_mul_else_land_12_lpi_1_dfm_10;
  reg [48:0] MulOut_data_10_sva_8;
  reg [48:0] MulOut_data_10_sva_9;
  reg [48:0] MulOut_data_10_sva_10;
  reg mul_loop_mul_else_land_11_lpi_1_dfm_7;
  reg mul_loop_mul_else_land_11_lpi_1_dfm_8;
  reg mul_loop_mul_else_land_11_lpi_1_dfm_9;
  reg mul_loop_mul_else_land_11_lpi_1_dfm_10;
  reg [48:0] MulOut_data_9_sva_8;
  reg [48:0] MulOut_data_9_sva_9;
  reg [48:0] MulOut_data_9_sva_10;
  reg mul_loop_mul_else_land_10_lpi_1_dfm_7;
  reg mul_loop_mul_else_land_10_lpi_1_dfm_8;
  reg mul_loop_mul_else_land_10_lpi_1_dfm_9;
  reg mul_loop_mul_else_land_10_lpi_1_dfm_10;
  reg [48:0] MulOut_data_8_sva_8;
  reg [48:0] MulOut_data_8_sva_9;
  reg [48:0] MulOut_data_8_sva_10;
  reg mul_loop_mul_else_land_9_lpi_1_dfm_7;
  reg mul_loop_mul_else_land_9_lpi_1_dfm_8;
  reg mul_loop_mul_else_land_9_lpi_1_dfm_9;
  reg mul_loop_mul_else_land_9_lpi_1_dfm_10;
  reg [48:0] MulOut_data_7_sva_8;
  reg [48:0] MulOut_data_7_sva_9;
  reg [48:0] MulOut_data_7_sva_10;
  reg mul_loop_mul_else_land_8_lpi_1_dfm_7;
  reg mul_loop_mul_else_land_8_lpi_1_dfm_8;
  reg mul_loop_mul_else_land_8_lpi_1_dfm_9;
  reg mul_loop_mul_else_land_8_lpi_1_dfm_10;
  reg [48:0] MulOut_data_6_sva_8;
  reg [48:0] MulOut_data_6_sva_9;
  reg [48:0] MulOut_data_6_sva_10;
  reg mul_loop_mul_else_land_7_lpi_1_dfm_7;
  reg mul_loop_mul_else_land_7_lpi_1_dfm_8;
  reg mul_loop_mul_else_land_7_lpi_1_dfm_9;
  reg mul_loop_mul_else_land_7_lpi_1_dfm_10;
  reg [48:0] MulOut_data_5_sva_8;
  reg [48:0] MulOut_data_5_sva_9;
  reg [48:0] MulOut_data_5_sva_10;
  reg mul_loop_mul_else_land_6_lpi_1_dfm_7;
  reg mul_loop_mul_else_land_6_lpi_1_dfm_8;
  reg mul_loop_mul_else_land_6_lpi_1_dfm_9;
  reg mul_loop_mul_else_land_6_lpi_1_dfm_10;
  reg [48:0] MulOut_data_4_sva_8;
  reg [48:0] MulOut_data_4_sva_9;
  reg [48:0] MulOut_data_4_sva_10;
  reg mul_loop_mul_else_land_5_lpi_1_dfm_7;
  reg mul_loop_mul_else_land_5_lpi_1_dfm_8;
  reg mul_loop_mul_else_land_5_lpi_1_dfm_9;
  reg mul_loop_mul_else_land_5_lpi_1_dfm_10;
  reg [48:0] MulOut_data_3_sva_8;
  reg [48:0] MulOut_data_3_sva_9;
  reg [48:0] MulOut_data_3_sva_10;
  reg mul_loop_mul_else_land_4_lpi_1_dfm_7;
  reg mul_loop_mul_else_land_4_lpi_1_dfm_8;
  reg mul_loop_mul_else_land_4_lpi_1_dfm_9;
  reg mul_loop_mul_else_land_4_lpi_1_dfm_10;
  reg [48:0] MulOut_data_2_sva_8;
  reg [48:0] MulOut_data_2_sva_9;
  reg [48:0] MulOut_data_2_sva_10;
  reg mul_loop_mul_else_land_3_lpi_1_dfm_7;
  reg mul_loop_mul_else_land_3_lpi_1_dfm_8;
  reg mul_loop_mul_else_land_3_lpi_1_dfm_9;
  reg mul_loop_mul_else_land_3_lpi_1_dfm_10;
  reg [48:0] MulOut_data_1_sva_8;
  reg [48:0] MulOut_data_1_sva_9;
  reg [48:0] MulOut_data_1_sva_10;
  reg mul_loop_mul_else_land_2_lpi_1_dfm_7;
  reg mul_loop_mul_else_land_2_lpi_1_dfm_8;
  reg mul_loop_mul_else_land_2_lpi_1_dfm_9;
  reg mul_loop_mul_else_land_2_lpi_1_dfm_10;
  reg [48:0] MulOut_data_0_sva_8;
  reg [48:0] MulOut_data_0_sva_9;
  reg [48:0] MulOut_data_0_sva_10;
  reg mul_loop_mul_else_land_1_lpi_1_dfm_7;
  reg mul_loop_mul_else_land_1_lpi_1_dfm_8;
  reg mul_loop_mul_else_land_1_lpi_1_dfm_9;
  reg mul_loop_mul_else_land_1_lpi_1_dfm_10;
  reg [15:0] cfg_mul_op_1_sva_1;
  reg cfg_mul_src_1_sva_1;
  reg [527:0] MulIn_data_sva_533;
  reg [527:0] MulIn_data_sva_534;
  reg [527:0] MulIn_data_sva_535;
  reg [527:0] MulIn_data_sva_536;
  reg io_read_cfg_mul_bypass_rsc_svs_5;
  reg io_read_cfg_mul_bypass_rsc_svs_6;
  reg io_read_cfg_mul_bypass_rsc_svs_7;
  reg io_read_cfg_mul_bypass_rsc_svs_8;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_10;
  reg IsZero_8U_23U_land_1_lpi_1_dfm_7;
  reg IsZero_8U_23U_land_1_lpi_1_dfm_5;
  reg IsZero_8U_23U_land_1_lpi_1_dfm_8;
  reg IsZero_8U_23U_1_land_1_lpi_1_dfm_6;
  reg IsZero_8U_23U_1_land_1_lpi_1_dfm_7;
  reg FpMul_8U_23U_lor_18_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_18_lpi_1_dfm_7;
  reg mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg FpMantRNE_48U_24U_else_carry_1_sva_2;
  reg mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs_2;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_10;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_10;
  reg IsZero_8U_23U_land_2_lpi_1_dfm_7;
  reg IsZero_8U_23U_land_2_lpi_1_dfm_5;
  reg IsZero_8U_23U_land_2_lpi_1_dfm_8;
  reg IsZero_8U_23U_1_land_2_lpi_1_dfm_6;
  reg IsZero_8U_23U_1_land_2_lpi_1_dfm_7;
  reg FpMul_8U_23U_lor_19_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_19_lpi_1_dfm_7;
  reg mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg FpMantRNE_48U_24U_else_carry_2_sva_2;
  reg mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs_2;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_10;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_10;
  reg IsZero_8U_23U_land_3_lpi_1_dfm_7;
  reg IsZero_8U_23U_land_3_lpi_1_dfm_5;
  reg IsZero_8U_23U_land_3_lpi_1_dfm_8;
  reg IsZero_8U_23U_1_land_3_lpi_1_dfm_6;
  reg IsZero_8U_23U_1_land_3_lpi_1_dfm_7;
  reg FpMul_8U_23U_lor_20_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_20_lpi_1_dfm_7;
  reg mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg FpMantRNE_48U_24U_else_carry_3_sva_2;
  reg mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs_2;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_10;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_10;
  reg IsZero_8U_23U_land_4_lpi_1_dfm_7;
  reg IsZero_8U_23U_land_4_lpi_1_dfm_5;
  reg IsZero_8U_23U_land_4_lpi_1_dfm_8;
  reg IsZero_8U_23U_1_land_4_lpi_1_dfm_4;
  reg IsZero_8U_23U_1_land_4_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_21_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_21_lpi_1_dfm_7;
  reg mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg FpMantRNE_48U_24U_else_carry_4_sva_2;
  reg mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs_2;
  reg IsNaN_8U_23U_land_4_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_4_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_4_lpi_1_dfm_10;
  reg IsNaN_8U_23U_land_4_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_10;
  reg IsZero_8U_23U_land_5_lpi_1_dfm_7;
  reg IsZero_8U_23U_land_5_lpi_1_dfm_5;
  reg IsZero_8U_23U_land_5_lpi_1_dfm_8;
  reg IsZero_8U_23U_1_land_5_lpi_1_dfm_6;
  reg IsZero_8U_23U_1_land_5_lpi_1_dfm_7;
  reg FpMul_8U_23U_lor_22_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_22_lpi_1_dfm_7;
  reg mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg FpMantRNE_48U_24U_else_carry_5_sva_2;
  reg mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs_2;
  reg IsNaN_8U_23U_land_5_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_5_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_5_lpi_1_dfm_10;
  reg IsNaN_8U_23U_land_5_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_10;
  reg IsZero_8U_23U_land_6_lpi_1_dfm_7;
  reg IsZero_8U_23U_land_6_lpi_1_dfm_5;
  reg IsZero_8U_23U_land_6_lpi_1_dfm_8;
  reg IsZero_8U_23U_1_land_6_lpi_1_dfm_4;
  reg IsZero_8U_23U_1_land_6_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_23_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_23_lpi_1_dfm_7;
  reg mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg FpMantRNE_48U_24U_else_carry_6_sva_2;
  reg mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs_2;
  reg IsNaN_8U_23U_land_6_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_6_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_6_lpi_1_dfm_10;
  reg IsNaN_8U_23U_land_6_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_10;
  reg IsZero_8U_23U_land_7_lpi_1_dfm_7;
  reg IsZero_8U_23U_land_7_lpi_1_dfm_5;
  reg IsZero_8U_23U_land_7_lpi_1_dfm_8;
  reg IsZero_8U_23U_1_land_7_lpi_1_dfm_4;
  reg IsZero_8U_23U_1_land_7_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_24_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_24_lpi_1_dfm_7;
  reg mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg FpMantRNE_48U_24U_else_carry_7_sva_2;
  reg mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs_2;
  reg IsNaN_8U_23U_land_7_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_7_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_7_lpi_1_dfm_10;
  reg IsNaN_8U_23U_land_7_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_10;
  reg IsZero_8U_23U_land_8_lpi_1_dfm_7;
  reg IsZero_8U_23U_land_8_lpi_1_dfm_5;
  reg IsZero_8U_23U_land_8_lpi_1_dfm_8;
  reg IsZero_8U_23U_1_land_8_lpi_1_dfm_6;
  reg IsZero_8U_23U_1_land_8_lpi_1_dfm_7;
  reg FpMul_8U_23U_lor_25_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_25_lpi_1_dfm_7;
  reg mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg FpMantRNE_48U_24U_else_carry_8_sva_2;
  reg mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs_2;
  reg IsNaN_8U_23U_land_8_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_8_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_8_lpi_1_dfm_10;
  reg IsNaN_8U_23U_land_8_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_10;
  reg IsZero_8U_23U_land_9_lpi_1_dfm_7;
  reg IsZero_8U_23U_land_9_lpi_1_dfm_5;
  reg IsZero_8U_23U_land_9_lpi_1_dfm_8;
  reg IsZero_8U_23U_1_land_9_lpi_1_dfm_6;
  reg IsZero_8U_23U_1_land_9_lpi_1_dfm_7;
  reg FpMul_8U_23U_lor_26_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_26_lpi_1_dfm_7;
  reg mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg FpMantRNE_48U_24U_else_carry_9_sva_2;
  reg mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs_2;
  reg IsNaN_8U_23U_land_9_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_9_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_9_lpi_1_dfm_10;
  reg IsNaN_8U_23U_land_9_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_10;
  reg IsZero_8U_23U_land_10_lpi_1_dfm_7;
  reg IsZero_8U_23U_land_10_lpi_1_dfm_5;
  reg IsZero_8U_23U_land_10_lpi_1_dfm_8;
  reg IsZero_8U_23U_1_land_10_lpi_1_dfm_4;
  reg IsZero_8U_23U_1_land_10_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_27_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_27_lpi_1_dfm_7;
  reg mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg FpMantRNE_48U_24U_else_carry_10_sva_2;
  reg mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs_2;
  reg IsNaN_8U_23U_land_10_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_10_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_10_lpi_1_dfm_10;
  reg IsNaN_8U_23U_land_10_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_10;
  reg IsZero_8U_23U_land_11_lpi_1_dfm_7;
  reg IsZero_8U_23U_land_11_lpi_1_dfm_5;
  reg IsZero_8U_23U_land_11_lpi_1_dfm_8;
  reg IsZero_8U_23U_1_land_11_lpi_1_dfm_4;
  reg IsZero_8U_23U_1_land_11_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_28_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_28_lpi_1_dfm_7;
  reg mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg FpMantRNE_48U_24U_else_carry_11_sva_2;
  reg mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs_2;
  reg IsNaN_8U_23U_land_11_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_11_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_11_lpi_1_dfm_10;
  reg IsNaN_8U_23U_land_11_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_10;
  reg IsZero_8U_23U_land_12_lpi_1_dfm_7;
  reg IsZero_8U_23U_land_12_lpi_1_dfm_5;
  reg IsZero_8U_23U_land_12_lpi_1_dfm_8;
  reg IsZero_8U_23U_1_land_12_lpi_1_dfm_4;
  reg IsZero_8U_23U_1_land_12_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_29_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_29_lpi_1_dfm_7;
  reg mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg FpMantRNE_48U_24U_else_carry_12_sva_2;
  reg mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs_2;
  reg IsNaN_8U_23U_land_12_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_12_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_12_lpi_1_dfm_10;
  reg IsNaN_8U_23U_land_12_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_10;
  reg IsZero_8U_23U_land_13_lpi_1_dfm_7;
  reg IsZero_8U_23U_land_13_lpi_1_dfm_5;
  reg IsZero_8U_23U_land_13_lpi_1_dfm_8;
  reg IsZero_8U_23U_1_land_13_lpi_1_dfm_6;
  reg IsZero_8U_23U_1_land_13_lpi_1_dfm_7;
  reg FpMul_8U_23U_lor_30_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_30_lpi_1_dfm_7;
  reg mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg FpMantRNE_48U_24U_else_carry_13_sva_2;
  reg mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs_2;
  reg IsNaN_8U_23U_land_13_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_13_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_13_lpi_1_dfm_10;
  reg IsNaN_8U_23U_land_13_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_10;
  reg IsZero_8U_23U_land_14_lpi_1_dfm_7;
  reg IsZero_8U_23U_land_14_lpi_1_dfm_5;
  reg IsZero_8U_23U_land_14_lpi_1_dfm_8;
  reg IsZero_8U_23U_1_land_14_lpi_1_dfm_4;
  reg IsZero_8U_23U_1_land_14_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_31_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_31_lpi_1_dfm_7;
  reg mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg FpMantRNE_48U_24U_else_carry_14_sva_2;
  reg mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs_2;
  reg IsNaN_8U_23U_land_14_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_14_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_14_lpi_1_dfm_10;
  reg IsNaN_8U_23U_land_14_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_10;
  reg IsZero_8U_23U_land_15_lpi_1_dfm_7;
  reg IsZero_8U_23U_land_15_lpi_1_dfm_5;
  reg IsZero_8U_23U_land_15_lpi_1_dfm_8;
  reg IsZero_8U_23U_1_land_15_lpi_1_dfm_6;
  reg IsZero_8U_23U_1_land_15_lpi_1_dfm_7;
  reg FpMul_8U_23U_lor_32_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_32_lpi_1_dfm_7;
  reg mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg FpMantRNE_48U_24U_else_carry_15_sva_2;
  reg mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs_2;
  reg IsNaN_8U_23U_land_15_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_15_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_15_lpi_1_dfm_10;
  reg IsNaN_8U_23U_land_15_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_10;
  reg IsZero_8U_23U_land_lpi_1_dfm_7;
  reg IsZero_8U_23U_land_lpi_1_dfm_5;
  reg IsZero_8U_23U_land_lpi_1_dfm_8;
  reg IsZero_8U_23U_1_land_lpi_1_dfm_6;
  reg IsZero_8U_23U_1_land_lpi_1_dfm_7;
  reg FpMul_8U_23U_lor_1_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_1_lpi_1_dfm_7;
  reg mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg FpMantRNE_48U_24U_else_carry_sva_2;
  reg mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs_2;
  reg IsNaN_8U_23U_land_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_lpi_1_dfm_10;
  reg IsNaN_8U_23U_land_lpi_1_dfm_11;
  reg cfg_mul_src_1_sva_st;
  reg mul_loop_mul_if_land_1_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_3_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_18_lpi_1_dfm_st;
  reg mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st;
  reg mul_loop_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_2;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_2;
  reg FpMul_8U_23U_FpMul_8U_23U_and_itm;
  reg FpMul_8U_23U_FpMul_8U_23U_and_itm_2;
  reg [22:0] mul_loop_mul_1_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2;
  reg [22:0] mul_loop_mul_1_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3;
  reg FpMul_8U_23U_mux_12_itm;
  reg FpMul_8U_23U_mux_12_itm_3;
  reg FpMul_8U_23U_mux_12_itm_4;
  reg mul_loop_mul_if_land_2_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_4_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_19_lpi_1_dfm_st;
  reg mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st;
  reg mul_loop_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_2;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_2;
  reg FpMul_8U_23U_FpMul_8U_23U_and_64_itm;
  reg FpMul_8U_23U_FpMul_8U_23U_and_64_itm_2;
  reg [22:0] mul_loop_mul_2_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2;
  reg [22:0] mul_loop_mul_2_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3;
  reg FpMul_8U_23U_mux_28_itm;
  reg FpMul_8U_23U_mux_28_itm_3;
  reg FpMul_8U_23U_mux_28_itm_4;
  reg mul_loop_mul_if_land_3_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_5_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_20_lpi_1_dfm_st;
  reg mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st;
  reg mul_loop_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_2;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_2;
  reg FpMul_8U_23U_FpMul_8U_23U_and_65_itm;
  reg FpMul_8U_23U_FpMul_8U_23U_and_65_itm_2;
  reg [22:0] mul_loop_mul_3_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2;
  reg [22:0] mul_loop_mul_3_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3;
  reg FpMul_8U_23U_mux_44_itm;
  reg FpMul_8U_23U_mux_44_itm_3;
  reg FpMul_8U_23U_mux_44_itm_4;
  reg mul_loop_mul_if_land_4_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_6_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_21_lpi_1_dfm_st;
  reg mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st;
  reg mul_loop_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_4_sva_st_2;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_2;
  reg FpMul_8U_23U_FpMul_8U_23U_and_66_itm;
  reg FpMul_8U_23U_FpMul_8U_23U_and_66_itm_2;
  reg [22:0] mul_loop_mul_4_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2;
  reg [22:0] mul_loop_mul_4_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3;
  reg FpMul_8U_23U_mux_60_itm;
  reg FpMul_8U_23U_mux_60_itm_3;
  reg FpMul_8U_23U_mux_60_itm_4;
  reg mul_loop_mul_if_land_5_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_7_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_22_lpi_1_dfm_st;
  reg mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st;
  reg mul_loop_mul_5_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_5_sva_st_2;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_4_itm;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_4_itm_2;
  reg FpMul_8U_23U_FpMul_8U_23U_and_67_itm;
  reg FpMul_8U_23U_FpMul_8U_23U_and_67_itm_2;
  reg [22:0] mul_loop_mul_5_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2;
  reg [22:0] mul_loop_mul_5_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3;
  reg FpMul_8U_23U_mux_76_itm;
  reg FpMul_8U_23U_mux_76_itm_3;
  reg FpMul_8U_23U_mux_76_itm_4;
  reg mul_loop_mul_if_land_6_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_8_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_23_lpi_1_dfm_st;
  reg mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st;
  reg mul_loop_mul_6_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_6_sva_st_2;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_5_itm;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_5_itm_2;
  reg FpMul_8U_23U_FpMul_8U_23U_and_68_itm;
  reg FpMul_8U_23U_FpMul_8U_23U_and_68_itm_2;
  reg [22:0] mul_loop_mul_6_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2;
  reg [22:0] mul_loop_mul_6_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3;
  reg FpMul_8U_23U_mux_92_itm;
  reg FpMul_8U_23U_mux_92_itm_3;
  reg FpMul_8U_23U_mux_92_itm_4;
  reg mul_loop_mul_if_land_7_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_9_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_24_lpi_1_dfm_st;
  reg mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st;
  reg mul_loop_mul_7_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_7_sva_st_2;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_6_itm;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_6_itm_2;
  reg FpMul_8U_23U_FpMul_8U_23U_and_69_itm;
  reg FpMul_8U_23U_FpMul_8U_23U_and_69_itm_2;
  reg [22:0] mul_loop_mul_7_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2;
  reg [22:0] mul_loop_mul_7_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3;
  reg FpMul_8U_23U_mux_108_itm;
  reg FpMul_8U_23U_mux_108_itm_3;
  reg FpMul_8U_23U_mux_108_itm_4;
  reg mul_loop_mul_if_land_8_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_10_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_25_lpi_1_dfm_st;
  reg mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st;
  reg mul_loop_mul_8_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_8_sva_st_2;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_7_itm;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_7_itm_2;
  reg FpMul_8U_23U_FpMul_8U_23U_and_70_itm;
  reg FpMul_8U_23U_FpMul_8U_23U_and_70_itm_2;
  reg [22:0] mul_loop_mul_8_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2;
  reg [22:0] mul_loop_mul_8_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3;
  reg FpMul_8U_23U_mux_124_itm;
  reg FpMul_8U_23U_mux_124_itm_3;
  reg FpMul_8U_23U_mux_124_itm_4;
  reg mul_loop_mul_if_land_9_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_11_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_26_lpi_1_dfm_st;
  reg mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st;
  reg mul_loop_mul_9_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_9_sva_st_2;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_8_itm;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_8_itm_2;
  reg FpMul_8U_23U_FpMul_8U_23U_and_71_itm;
  reg FpMul_8U_23U_FpMul_8U_23U_and_71_itm_2;
  reg [22:0] mul_loop_mul_9_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2;
  reg [22:0] mul_loop_mul_9_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3;
  reg FpMul_8U_23U_mux_140_itm;
  reg FpMul_8U_23U_mux_140_itm_3;
  reg FpMul_8U_23U_mux_140_itm_4;
  reg mul_loop_mul_if_land_10_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_12_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_27_lpi_1_dfm_st;
  reg mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st;
  reg mul_loop_mul_10_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_10_sva_st_2;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_9_itm;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_9_itm_2;
  reg FpMul_8U_23U_FpMul_8U_23U_and_72_itm;
  reg FpMul_8U_23U_FpMul_8U_23U_and_72_itm_2;
  reg [22:0] mul_loop_mul_10_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2;
  reg [22:0] mul_loop_mul_10_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3;
  reg FpMul_8U_23U_mux_156_itm;
  reg FpMul_8U_23U_mux_156_itm_3;
  reg FpMul_8U_23U_mux_156_itm_4;
  reg mul_loop_mul_if_land_11_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_13_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_28_lpi_1_dfm_st;
  reg mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st;
  reg mul_loop_mul_11_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_11_sva_st_2;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_10_itm;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_10_itm_2;
  reg FpMul_8U_23U_FpMul_8U_23U_and_73_itm;
  reg FpMul_8U_23U_FpMul_8U_23U_and_73_itm_2;
  reg [22:0] mul_loop_mul_11_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2;
  reg [22:0] mul_loop_mul_11_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3;
  reg FpMul_8U_23U_mux_172_itm;
  reg FpMul_8U_23U_mux_172_itm_3;
  reg FpMul_8U_23U_mux_172_itm_4;
  reg mul_loop_mul_if_land_12_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_14_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_29_lpi_1_dfm_st;
  reg mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st;
  reg mul_loop_mul_12_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_12_sva_st_2;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_11_itm;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_11_itm_2;
  reg FpMul_8U_23U_FpMul_8U_23U_and_74_itm;
  reg FpMul_8U_23U_FpMul_8U_23U_and_74_itm_2;
  reg [22:0] mul_loop_mul_12_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2;
  reg [22:0] mul_loop_mul_12_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3;
  reg FpMul_8U_23U_mux_188_itm;
  reg FpMul_8U_23U_mux_188_itm_3;
  reg FpMul_8U_23U_mux_188_itm_4;
  reg mul_loop_mul_if_land_13_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_15_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_30_lpi_1_dfm_st;
  reg mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st;
  reg mul_loop_mul_13_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_13_sva_st_2;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_12_itm;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_12_itm_2;
  reg FpMul_8U_23U_FpMul_8U_23U_and_75_itm;
  reg FpMul_8U_23U_FpMul_8U_23U_and_75_itm_2;
  reg [22:0] mul_loop_mul_13_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2;
  reg [22:0] mul_loop_mul_13_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3;
  reg FpMul_8U_23U_mux_204_itm;
  reg FpMul_8U_23U_mux_204_itm_3;
  reg FpMul_8U_23U_mux_204_itm_4;
  reg mul_loop_mul_if_land_14_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_16_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_31_lpi_1_dfm_st;
  reg mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st;
  reg mul_loop_mul_14_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_14_sva_st_2;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_13_itm;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_13_itm_2;
  reg FpMul_8U_23U_FpMul_8U_23U_and_76_itm;
  reg FpMul_8U_23U_FpMul_8U_23U_and_76_itm_2;
  reg [22:0] mul_loop_mul_14_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2;
  reg [22:0] mul_loop_mul_14_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3;
  reg FpMul_8U_23U_mux_220_itm;
  reg FpMul_8U_23U_mux_220_itm_3;
  reg FpMul_8U_23U_mux_220_itm_4;
  reg mul_loop_mul_if_land_15_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_17_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_32_lpi_1_dfm_st;
  reg mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st;
  reg mul_loop_mul_15_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_15_sva_st_2;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_14_itm;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_14_itm_2;
  reg FpMul_8U_23U_FpMul_8U_23U_and_77_itm;
  reg FpMul_8U_23U_FpMul_8U_23U_and_77_itm_2;
  reg [22:0] mul_loop_mul_15_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2;
  reg [22:0] mul_loop_mul_15_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3;
  reg FpMul_8U_23U_mux_236_itm;
  reg FpMul_8U_23U_mux_236_itm_3;
  reg FpMul_8U_23U_mux_236_itm_4;
  reg mul_loop_mul_if_land_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_lpi_1_dfm_st;
  reg FpMul_8U_23U_lor_1_lpi_1_dfm_st;
  reg mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st;
  reg mul_loop_mul_16_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_2;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_15_itm;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_15_itm_2;
  reg FpMul_8U_23U_FpMul_8U_23U_and_78_itm;
  reg FpMul_8U_23U_FpMul_8U_23U_and_78_itm_2;
  reg [22:0] mul_loop_mul_16_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2;
  reg [22:0] mul_loop_mul_16_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3;
  reg FpMul_8U_23U_mux_252_itm;
  reg FpMul_8U_23U_mux_252_itm_3;
  reg FpMul_8U_23U_mux_252_itm_4;
  reg io_read_cfg_mul_bypass_rsc_svs_st_1;
  reg cfg_mul_src_1_sva_st_1;
  reg io_read_cfg_mul_bypass_rsc_svs_st_5;
  reg io_read_cfg_mul_bypass_rsc_svs_st_6;
  reg io_read_cfg_mul_bypass_rsc_svs_st_7;
  reg mul_loop_mul_if_land_1_lpi_1_dfm_st_5;
  reg mul_loop_mul_if_land_1_lpi_1_dfm_st_6;
  reg mul_loop_mul_if_land_1_lpi_1_dfm_st_7;
  reg FpMul_8U_23U_lor_18_lpi_1_dfm_st_3;
  reg mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  reg mul_loop_mul_if_land_1_lpi_1_dfm_st_8;
  reg FpMul_8U_23U_lor_18_lpi_1_dfm_st_4;
  reg mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  reg mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs_st_2;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_st_6;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_st_7;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_st_8;
  reg mul_loop_mul_if_land_2_lpi_1_dfm_st_5;
  reg mul_loop_mul_if_land_2_lpi_1_dfm_st_6;
  reg mul_loop_mul_if_land_2_lpi_1_dfm_st_7;
  reg FpMul_8U_23U_lor_19_lpi_1_dfm_st_3;
  reg mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  reg mul_loop_mul_if_land_2_lpi_1_dfm_st_8;
  reg FpMul_8U_23U_lor_19_lpi_1_dfm_st_4;
  reg mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  reg mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs_st_2;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_st_6;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_st_7;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_st_8;
  reg mul_loop_mul_if_land_3_lpi_1_dfm_st_5;
  reg mul_loop_mul_if_land_3_lpi_1_dfm_st_6;
  reg mul_loop_mul_if_land_3_lpi_1_dfm_st_7;
  reg FpMul_8U_23U_lor_20_lpi_1_dfm_st_3;
  reg mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  reg mul_loop_mul_if_land_3_lpi_1_dfm_st_8;
  reg FpMul_8U_23U_lor_20_lpi_1_dfm_st_4;
  reg mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  reg mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs_st_2;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_st_6;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_st_7;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_st_8;
  reg mul_loop_mul_if_land_4_lpi_1_dfm_st_5;
  reg mul_loop_mul_if_land_4_lpi_1_dfm_st_6;
  reg mul_loop_mul_if_land_4_lpi_1_dfm_st_7;
  reg FpMul_8U_23U_lor_21_lpi_1_dfm_st_3;
  reg mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  reg mul_loop_mul_if_land_4_lpi_1_dfm_st_8;
  reg FpMul_8U_23U_lor_21_lpi_1_dfm_st_4;
  reg mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  reg mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs_st_2;
  reg IsNaN_8U_23U_land_4_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_land_4_lpi_1_dfm_st_6;
  reg IsNaN_8U_23U_land_4_lpi_1_dfm_st_7;
  reg IsNaN_8U_23U_land_4_lpi_1_dfm_st_8;
  reg mul_loop_mul_if_land_5_lpi_1_dfm_st_5;
  reg mul_loop_mul_if_land_5_lpi_1_dfm_st_6;
  reg mul_loop_mul_if_land_5_lpi_1_dfm_st_7;
  reg FpMul_8U_23U_lor_22_lpi_1_dfm_st_3;
  reg mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  reg mul_loop_mul_if_land_5_lpi_1_dfm_st_8;
  reg FpMul_8U_23U_lor_22_lpi_1_dfm_st_4;
  reg mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  reg mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs_st_2;
  reg IsNaN_8U_23U_land_5_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_land_5_lpi_1_dfm_st_6;
  reg IsNaN_8U_23U_land_5_lpi_1_dfm_st_7;
  reg IsNaN_8U_23U_land_5_lpi_1_dfm_st_8;
  reg mul_loop_mul_if_land_6_lpi_1_dfm_st_5;
  reg mul_loop_mul_if_land_6_lpi_1_dfm_st_6;
  reg mul_loop_mul_if_land_6_lpi_1_dfm_st_7;
  reg FpMul_8U_23U_lor_23_lpi_1_dfm_st_3;
  reg mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  reg mul_loop_mul_if_land_6_lpi_1_dfm_st_8;
  reg FpMul_8U_23U_lor_23_lpi_1_dfm_st_4;
  reg mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  reg mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs_st_2;
  reg IsNaN_8U_23U_land_6_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_land_6_lpi_1_dfm_st_6;
  reg IsNaN_8U_23U_land_6_lpi_1_dfm_st_7;
  reg IsNaN_8U_23U_land_6_lpi_1_dfm_st_8;
  reg mul_loop_mul_if_land_7_lpi_1_dfm_st_5;
  reg mul_loop_mul_if_land_7_lpi_1_dfm_st_6;
  reg mul_loop_mul_if_land_7_lpi_1_dfm_st_7;
  reg FpMul_8U_23U_lor_24_lpi_1_dfm_st_3;
  reg mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  reg mul_loop_mul_if_land_7_lpi_1_dfm_st_8;
  reg FpMul_8U_23U_lor_24_lpi_1_dfm_st_4;
  reg mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  reg mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs_st_2;
  reg IsNaN_8U_23U_land_7_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_land_7_lpi_1_dfm_st_6;
  reg IsNaN_8U_23U_land_7_lpi_1_dfm_st_7;
  reg IsNaN_8U_23U_land_7_lpi_1_dfm_st_8;
  reg mul_loop_mul_if_land_8_lpi_1_dfm_st_5;
  reg mul_loop_mul_if_land_8_lpi_1_dfm_st_6;
  reg mul_loop_mul_if_land_8_lpi_1_dfm_st_7;
  reg FpMul_8U_23U_lor_25_lpi_1_dfm_st_3;
  reg mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  reg mul_loop_mul_if_land_8_lpi_1_dfm_st_8;
  reg FpMul_8U_23U_lor_25_lpi_1_dfm_st_4;
  reg mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  reg mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs_st_2;
  reg IsNaN_8U_23U_land_8_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_land_8_lpi_1_dfm_st_6;
  reg IsNaN_8U_23U_land_8_lpi_1_dfm_st_7;
  reg IsNaN_8U_23U_land_8_lpi_1_dfm_st_8;
  reg mul_loop_mul_if_land_9_lpi_1_dfm_st_5;
  reg mul_loop_mul_if_land_9_lpi_1_dfm_st_6;
  reg mul_loop_mul_if_land_9_lpi_1_dfm_st_7;
  reg FpMul_8U_23U_lor_26_lpi_1_dfm_st_3;
  reg mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  reg mul_loop_mul_if_land_9_lpi_1_dfm_st_8;
  reg FpMul_8U_23U_lor_26_lpi_1_dfm_st_4;
  reg mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  reg mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs_st_2;
  reg IsNaN_8U_23U_land_9_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_land_9_lpi_1_dfm_st_6;
  reg IsNaN_8U_23U_land_9_lpi_1_dfm_st_7;
  reg IsNaN_8U_23U_land_9_lpi_1_dfm_st_8;
  reg mul_loop_mul_if_land_10_lpi_1_dfm_st_5;
  reg mul_loop_mul_if_land_10_lpi_1_dfm_st_6;
  reg mul_loop_mul_if_land_10_lpi_1_dfm_st_7;
  reg FpMul_8U_23U_lor_27_lpi_1_dfm_st_3;
  reg mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  reg mul_loop_mul_if_land_10_lpi_1_dfm_st_8;
  reg FpMul_8U_23U_lor_27_lpi_1_dfm_st_4;
  reg mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  reg mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs_st_2;
  reg IsNaN_8U_23U_land_10_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_land_10_lpi_1_dfm_st_6;
  reg IsNaN_8U_23U_land_10_lpi_1_dfm_st_7;
  reg IsNaN_8U_23U_land_10_lpi_1_dfm_st_8;
  reg mul_loop_mul_if_land_11_lpi_1_dfm_st_5;
  reg mul_loop_mul_if_land_11_lpi_1_dfm_st_6;
  reg mul_loop_mul_if_land_11_lpi_1_dfm_st_7;
  reg FpMul_8U_23U_lor_28_lpi_1_dfm_st_3;
  reg mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  reg mul_loop_mul_if_land_11_lpi_1_dfm_st_8;
  reg FpMul_8U_23U_lor_28_lpi_1_dfm_st_4;
  reg mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  reg mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs_st_2;
  reg IsNaN_8U_23U_land_11_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_land_11_lpi_1_dfm_st_6;
  reg IsNaN_8U_23U_land_11_lpi_1_dfm_st_7;
  reg IsNaN_8U_23U_land_11_lpi_1_dfm_st_8;
  reg mul_loop_mul_if_land_12_lpi_1_dfm_st_5;
  reg mul_loop_mul_if_land_12_lpi_1_dfm_st_6;
  reg mul_loop_mul_if_land_12_lpi_1_dfm_st_7;
  reg FpMul_8U_23U_lor_29_lpi_1_dfm_st_3;
  reg mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  reg mul_loop_mul_if_land_12_lpi_1_dfm_st_8;
  reg FpMul_8U_23U_lor_29_lpi_1_dfm_st_4;
  reg mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  reg mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs_st_2;
  reg IsNaN_8U_23U_land_12_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_land_12_lpi_1_dfm_st_6;
  reg IsNaN_8U_23U_land_12_lpi_1_dfm_st_7;
  reg IsNaN_8U_23U_land_12_lpi_1_dfm_st_8;
  reg mul_loop_mul_if_land_13_lpi_1_dfm_st_5;
  reg mul_loop_mul_if_land_13_lpi_1_dfm_st_6;
  reg mul_loop_mul_if_land_13_lpi_1_dfm_st_7;
  reg FpMul_8U_23U_lor_30_lpi_1_dfm_st_3;
  reg mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  reg mul_loop_mul_if_land_13_lpi_1_dfm_st_8;
  reg FpMul_8U_23U_lor_30_lpi_1_dfm_st_4;
  reg mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  reg mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs_st_2;
  reg IsNaN_8U_23U_land_13_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_land_13_lpi_1_dfm_st_6;
  reg IsNaN_8U_23U_land_13_lpi_1_dfm_st_7;
  reg IsNaN_8U_23U_land_13_lpi_1_dfm_st_8;
  reg mul_loop_mul_if_land_14_lpi_1_dfm_st_5;
  reg mul_loop_mul_if_land_14_lpi_1_dfm_st_6;
  reg mul_loop_mul_if_land_14_lpi_1_dfm_st_7;
  reg FpMul_8U_23U_lor_31_lpi_1_dfm_st_3;
  reg mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  reg mul_loop_mul_if_land_14_lpi_1_dfm_st_8;
  reg FpMul_8U_23U_lor_31_lpi_1_dfm_st_4;
  reg mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  reg mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs_st_2;
  reg IsNaN_8U_23U_land_14_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_land_14_lpi_1_dfm_st_6;
  reg IsNaN_8U_23U_land_14_lpi_1_dfm_st_7;
  reg IsNaN_8U_23U_land_14_lpi_1_dfm_st_8;
  reg mul_loop_mul_if_land_15_lpi_1_dfm_st_5;
  reg mul_loop_mul_if_land_15_lpi_1_dfm_st_6;
  reg mul_loop_mul_if_land_15_lpi_1_dfm_st_7;
  reg FpMul_8U_23U_lor_32_lpi_1_dfm_st_3;
  reg mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  reg mul_loop_mul_if_land_15_lpi_1_dfm_st_8;
  reg FpMul_8U_23U_lor_32_lpi_1_dfm_st_4;
  reg mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  reg mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs_st_2;
  reg IsNaN_8U_23U_land_15_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_land_15_lpi_1_dfm_st_6;
  reg IsNaN_8U_23U_land_15_lpi_1_dfm_st_7;
  reg IsNaN_8U_23U_land_15_lpi_1_dfm_st_8;
  reg mul_loop_mul_if_land_lpi_1_dfm_st_5;
  reg mul_loop_mul_if_land_lpi_1_dfm_st_6;
  reg mul_loop_mul_if_land_lpi_1_dfm_st_7;
  reg FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
  reg mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  reg mul_loop_mul_if_land_lpi_1_dfm_st_8;
  reg FpMul_8U_23U_lor_1_lpi_1_dfm_st_4;
  reg mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  reg mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs_st_2;
  reg IsNaN_8U_23U_land_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_land_lpi_1_dfm_st_6;
  reg IsNaN_8U_23U_land_lpi_1_dfm_st_7;
  reg IsNaN_8U_23U_land_lpi_1_dfm_st_8;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_9_0;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_3_2;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_1_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_9_0;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_3_2;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_1_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_9_0;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_3_2;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_1_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_9_0;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_3_2;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_1_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_9_0;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_3_2;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_1_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_9_0;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_3_2;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_1_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_9_0;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_3_2;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_1_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_9_0;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_3_2;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_1_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_9_0;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_3_2;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_1_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_9_0;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_3_2;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_1_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_9_0;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_3_2;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_1_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_9_0;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_3_2;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_1_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_9_0;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_3_2;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_1_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_9_0;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_3_2;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_1_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_9_0;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_3_2;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_1_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_22_13;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_12_10;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_9_0;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_3_2;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_1_0;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_9_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_9_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_9_9_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_7_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_7_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_8_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_8_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_9_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_9_1_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_9_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_9_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_9_9_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_7_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_7_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_8_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_8_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_9_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_9_1_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_9_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_9_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_9_9_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_7_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_7_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_8_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_8_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_9_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_9_1_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_9_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_9_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_9_9_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_7_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_7_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_8_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_8_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_9_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_9_1_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_9_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_9_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_9_9_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_7_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_7_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_8_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_8_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_9_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_9_1_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_9_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_9_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_9_9_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_7_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_7_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_8_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_8_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_9_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_9_1_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_9_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_9_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_9_9_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_7_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_7_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_8_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_8_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_9_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_9_1_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_9_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_9_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_9_9_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_7_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_7_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_8_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_8_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_9_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_9_1_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_9_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_9_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_9_9_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_7_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_7_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_8_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_8_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_9_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_9_1_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_9_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_9_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_9_9_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_7_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_7_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_8_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_8_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_9_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_9_1_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_9_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_9_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_9_9_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_7_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_7_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_8_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_8_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_9_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_9_1_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_9_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_9_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_9_9_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_7_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_7_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_8_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_8_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_9_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_9_1_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_9_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_9_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_9_9_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_7_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_7_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_8_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_8_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_9_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_9_1_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_9_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_9_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_9_9_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_7_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_7_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_8_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_8_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_9_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_9_1_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_9_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_9_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_9_9_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_7_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_7_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_8_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_8_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_9_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_9_1_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_9_0_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_9_22_13_1;
  reg [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_9_12_10_1;
  reg [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_9_9_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_7_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_7_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_8_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_8_1_0_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_9_3_2_1;
  reg [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_9_1_0_1;
  wire and_1647_cse;
  wire main_stage_en_1;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_sva;
  wire [4:0] else_MulOp_data_15_14_10_lpi_1_dfm_mx0;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_15_sva;
  wire [4:0] else_MulOp_data_14_14_10_lpi_1_dfm_mx0;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_14_sva;
  wire [4:0] else_MulOp_data_13_14_10_lpi_1_dfm_mx0;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_13_sva;
  wire [4:0] else_MulOp_data_12_14_10_lpi_1_dfm_mx0;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_12_sva;
  wire [4:0] else_MulOp_data_11_14_10_lpi_1_dfm_mx0;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_11_sva;
  wire [4:0] else_MulOp_data_10_14_10_lpi_1_dfm_mx0;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_10_sva;
  wire [4:0] else_MulOp_data_9_14_10_lpi_1_dfm_mx0;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_9_sva;
  wire [4:0] else_MulOp_data_8_14_10_lpi_1_dfm_mx0;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_8_sva;
  wire [4:0] else_MulOp_data_7_14_10_lpi_1_dfm_mx0;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_7_sva;
  wire [4:0] else_MulOp_data_6_14_10_lpi_1_dfm_mx0;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_6_sva;
  wire [4:0] else_MulOp_data_5_14_10_lpi_1_dfm_mx0;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_5_sva;
  wire [4:0] else_MulOp_data_4_14_10_lpi_1_dfm_mx0;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_4_sva;
  wire [4:0] else_MulOp_data_3_14_10_lpi_1_dfm_mx0;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_3_sva;
  wire [4:0] else_MulOp_data_2_14_10_lpi_1_dfm_mx0;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_2_sva;
  wire [4:0] else_MulOp_data_1_14_10_lpi_1_dfm_mx0;
  wire IsZero_5U_23U_IsZero_5U_23U_nor_cse_1_sva;
  wire [4:0] else_MulOp_data_0_14_10_lpi_1_dfm_mx0;
  wire or_17_ssc;
  wire and_116_ssc;
  wire and_1_m1c;
  wire nor_m1c;
  wire or_1_ssc;
  wire and_51_ssc;
  wire or_2_ssc;
  wire and_55_ssc;
  wire or_3_ssc;
  wire and_59_ssc;
  wire or_4_ssc;
  wire and_63_ssc;
  wire or_5_ssc;
  wire and_67_ssc;
  wire or_6_ssc;
  wire and_71_ssc;
  wire or_7_ssc;
  wire and_75_ssc;
  wire or_8_ssc;
  wire and_79_ssc;
  wire or_9_ssc;
  wire and_83_ssc;
  wire or_10_ssc;
  wire and_87_ssc;
  wire or_11_ssc;
  wire and_91_ssc;
  wire or_12_ssc;
  wire and_95_ssc;
  wire or_13_ssc;
  wire and_99_ssc;
  wire or_14_ssc;
  wire and_103_ssc;
  wire or_15_ssc;
  wire and_107_ssc;
  wire else_unequal_tmp;
  wire FpMul_8U_23U_is_inf_lpi_1_dfm_2;
  wire FpMul_8U_23U_is_inf_15_lpi_1_dfm_2;
  wire FpMul_8U_23U_is_inf_14_lpi_1_dfm_2;
  wire FpMul_8U_23U_is_inf_13_lpi_1_dfm_2;
  wire FpMul_8U_23U_is_inf_12_lpi_1_dfm_2;
  wire FpMul_8U_23U_is_inf_11_lpi_1_dfm_2;
  wire FpMul_8U_23U_is_inf_10_lpi_1_dfm_2;
  wire FpMul_8U_23U_is_inf_9_lpi_1_dfm_2;
  wire FpMul_8U_23U_is_inf_8_lpi_1_dfm_2;
  wire FpMul_8U_23U_is_inf_7_lpi_1_dfm_2;
  wire FpMul_8U_23U_is_inf_6_lpi_1_dfm_2;
  wire FpMul_8U_23U_is_inf_5_lpi_1_dfm_2;
  wire FpMul_8U_23U_is_inf_4_lpi_1_dfm_2;
  wire FpMul_8U_23U_is_inf_3_lpi_1_dfm_2;
  wire FpMul_8U_23U_is_inf_2_lpi_1_dfm_2;
  wire FpMul_8U_23U_is_inf_1_lpi_1_dfm_2;
  wire IsDenorm_5U_23U_land_lpi_1_dfm;
  wire IsInf_5U_23U_land_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_15_cse;
  wire IsDenorm_5U_23U_land_15_lpi_1_dfm;
  wire IsInf_5U_23U_land_15_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_14_cse;
  wire IsZero_8U_23U_1_land_14_lpi_1_dfm_mx0w0;
  wire IsDenorm_5U_23U_land_14_lpi_1_dfm;
  wire IsInf_5U_23U_land_14_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_13_cse;
  wire IsDenorm_5U_23U_land_13_lpi_1_dfm;
  wire IsInf_5U_23U_land_13_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_12_cse;
  wire IsZero_8U_23U_1_land_12_lpi_1_dfm_mx0w0;
  wire IsDenorm_5U_23U_land_12_lpi_1_dfm;
  wire IsInf_5U_23U_land_12_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_11_cse;
  wire IsZero_8U_23U_1_land_11_lpi_1_dfm_mx0w0;
  wire IsDenorm_5U_23U_land_11_lpi_1_dfm;
  wire IsInf_5U_23U_land_11_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_10_cse;
  wire IsZero_8U_23U_1_land_10_lpi_1_dfm_mx0w0;
  wire IsDenorm_5U_23U_land_10_lpi_1_dfm;
  wire IsInf_5U_23U_land_10_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_9_cse;
  wire IsDenorm_5U_23U_land_9_lpi_1_dfm;
  wire IsInf_5U_23U_land_9_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_8_cse;
  wire IsDenorm_5U_23U_land_8_lpi_1_dfm;
  wire IsInf_5U_23U_land_8_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_7_cse;
  wire IsZero_8U_23U_1_land_7_lpi_1_dfm_mx0w0;
  wire IsDenorm_5U_23U_land_7_lpi_1_dfm;
  wire IsInf_5U_23U_land_7_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_6_cse;
  wire IsZero_8U_23U_1_land_6_lpi_1_dfm_mx0w0;
  wire IsDenorm_5U_23U_land_6_lpi_1_dfm;
  wire IsInf_5U_23U_land_6_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_5_cse;
  wire IsDenorm_5U_23U_land_5_lpi_1_dfm;
  wire IsInf_5U_23U_land_5_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_4_cse;
  wire IsZero_8U_23U_1_land_4_lpi_1_dfm_mx0w0;
  wire IsDenorm_5U_23U_land_4_lpi_1_dfm;
  wire IsInf_5U_23U_land_4_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_3_cse;
  wire IsDenorm_5U_23U_land_3_lpi_1_dfm;
  wire IsInf_5U_23U_land_3_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_2_cse;
  wire IsDenorm_5U_23U_land_2_lpi_1_dfm;
  wire IsInf_5U_23U_land_2_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_1_cse;
  wire IsDenorm_5U_23U_land_1_lpi_1_dfm;
  wire IsInf_5U_23U_land_1_lpi_1_dfm;
  wire IsNaN_5U_23U_IsNaN_5U_23U_nand_cse;
  wire FpMantRNE_48U_24U_else_carry_sva_mx0w0;
  wire FpMantRNE_48U_24U_else_carry_15_sva_mx0w0;
  wire FpMantRNE_48U_24U_else_carry_14_sva_mx0w0;
  wire FpMantRNE_48U_24U_else_carry_13_sva_mx0w0;
  wire FpMantRNE_48U_24U_else_carry_12_sva_mx0w0;
  wire FpMantRNE_48U_24U_else_carry_11_sva_mx0w0;
  wire FpMantRNE_48U_24U_else_carry_10_sva_mx0w0;
  wire FpMantRNE_48U_24U_else_carry_9_sva_mx0w0;
  wire FpMantRNE_48U_24U_else_carry_8_sva_mx0w0;
  wire FpMantRNE_48U_24U_else_carry_7_sva_mx0w0;
  wire FpMantRNE_48U_24U_else_carry_6_sva_mx0w0;
  wire FpMantRNE_48U_24U_else_carry_5_sva_mx0w0;
  wire FpMantRNE_48U_24U_else_carry_4_sva_mx0w0;
  wire FpMantRNE_48U_24U_else_carry_3_sva_mx0w0;
  wire FpMantRNE_48U_24U_else_carry_2_sva_mx0w0;
  wire FpMantRNE_48U_24U_else_carry_1_sva_mx0w0;
  wire mul_nan_to_zero_land_lpi_1_dfm;
  wire mul_nan_to_zero_land_15_lpi_1_dfm;
  wire mul_nan_to_zero_land_14_lpi_1_dfm;
  wire mul_nan_to_zero_land_13_lpi_1_dfm;
  wire mul_nan_to_zero_land_12_lpi_1_dfm;
  wire mul_nan_to_zero_land_11_lpi_1_dfm;
  wire mul_nan_to_zero_land_10_lpi_1_dfm;
  wire mul_nan_to_zero_land_9_lpi_1_dfm;
  wire mul_nan_to_zero_land_8_lpi_1_dfm;
  wire mul_nan_to_zero_land_7_lpi_1_dfm;
  wire mul_nan_to_zero_land_6_lpi_1_dfm;
  wire mul_nan_to_zero_land_5_lpi_1_dfm;
  wire mul_nan_to_zero_land_4_lpi_1_dfm;
  wire mul_nan_to_zero_land_3_lpi_1_dfm;
  wire mul_nan_to_zero_land_2_lpi_1_dfm;
  wire mul_nan_to_zero_land_1_lpi_1_dfm;
  wire [3:0] FpMul_8U_23U_o_expo_7_4_lpi_1_dfm;
  wire [3:0] FpMul_8U_23U_o_expo_3_0_lpi_1_dfm_mx1;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_lpi_1_dfm_1;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_15;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1;
  wire [3:0] FpMul_8U_23U_o_expo_7_4_15_lpi_1_dfm;
  wire [3:0] FpMul_8U_23U_o_expo_3_0_15_lpi_1_dfm_mx1;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_15_lpi_1_dfm_1;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_14;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_15_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_15_sva_1;
  wire [3:0] FpMul_8U_23U_o_expo_7_4_14_lpi_1_dfm;
  wire [3:0] FpMul_8U_23U_o_expo_3_0_14_lpi_1_dfm_mx1;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_14_lpi_1_dfm_1;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_13;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_14_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_14_sva_1;
  wire [3:0] FpMul_8U_23U_o_expo_7_4_13_lpi_1_dfm;
  wire [3:0] FpMul_8U_23U_o_expo_3_0_13_lpi_1_dfm_mx1;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_13_lpi_1_dfm_1;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_12;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_13_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_13_sva_1;
  wire [3:0] FpMul_8U_23U_o_expo_7_4_12_lpi_1_dfm;
  wire [3:0] FpMul_8U_23U_o_expo_3_0_12_lpi_1_dfm_mx1;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_12_lpi_1_dfm_1;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_11;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_12_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_12_sva_1;
  wire [3:0] FpMul_8U_23U_o_expo_7_4_11_lpi_1_dfm;
  wire [3:0] FpMul_8U_23U_o_expo_3_0_11_lpi_1_dfm_mx1;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_11_lpi_1_dfm_1;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_10;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_11_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_11_sva_1;
  wire [3:0] FpMul_8U_23U_o_expo_7_4_10_lpi_1_dfm;
  wire [3:0] FpMul_8U_23U_o_expo_3_0_10_lpi_1_dfm_mx1;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_10_lpi_1_dfm_1;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_9;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_10_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_10_sva_1;
  wire [3:0] FpMul_8U_23U_o_expo_7_4_9_lpi_1_dfm;
  wire [3:0] FpMul_8U_23U_o_expo_3_0_9_lpi_1_dfm_mx1;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_9_lpi_1_dfm_1;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_8;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_9_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_9_sva_1;
  wire [3:0] FpMul_8U_23U_o_expo_7_4_8_lpi_1_dfm;
  wire [3:0] FpMul_8U_23U_o_expo_3_0_8_lpi_1_dfm_mx1;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_8_lpi_1_dfm_1;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_7;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_8_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_8_sva_1;
  wire [3:0] FpMul_8U_23U_o_expo_7_4_7_lpi_1_dfm;
  wire [3:0] FpMul_8U_23U_o_expo_3_0_7_lpi_1_dfm_mx1;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_7_lpi_1_dfm_1;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_6;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_7_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_7_sva_1;
  wire [3:0] FpMul_8U_23U_o_expo_7_4_6_lpi_1_dfm;
  wire [3:0] FpMul_8U_23U_o_expo_3_0_6_lpi_1_dfm_mx1;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_6_lpi_1_dfm_1;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_5;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_6_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_6_sva_1;
  wire [3:0] FpMul_8U_23U_o_expo_7_4_5_lpi_1_dfm;
  wire [3:0] FpMul_8U_23U_o_expo_3_0_5_lpi_1_dfm_mx1;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_5_lpi_1_dfm_1;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_4;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_5_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_5_sva_1;
  wire [3:0] FpMul_8U_23U_o_expo_7_4_4_lpi_1_dfm;
  wire [3:0] FpMul_8U_23U_o_expo_3_0_4_lpi_1_dfm_mx1;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_4_lpi_1_dfm_1;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_3;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_4_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_4_sva_1;
  wire [3:0] FpMul_8U_23U_o_expo_7_4_3_lpi_1_dfm;
  wire [3:0] FpMul_8U_23U_o_expo_3_0_3_lpi_1_dfm_mx1;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_lpi_1_dfm_1;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_2;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1;
  wire [3:0] FpMul_8U_23U_o_expo_7_4_2_lpi_1_dfm;
  wire [3:0] FpMul_8U_23U_o_expo_3_0_2_lpi_1_dfm_mx1;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_lpi_1_dfm_1;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_1;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1;
  wire [3:0] FpMul_8U_23U_o_expo_7_4_1_lpi_1_dfm;
  wire [3:0] FpMul_8U_23U_o_expo_3_0_1_lpi_1_dfm_mx1;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_lpi_1_dfm_1;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_15_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_15_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_14_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_14_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_13_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_13_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_12_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_12_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_11_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_11_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_10_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_10_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_9_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_9_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_8_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_8_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_7_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_7_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_6_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_6_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_5_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_5_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_4_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_4_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_3_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_3_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_2_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_2_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_1_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_1_lpi_1_dfm;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0;
  wire [9:0] mul_nan_to_zero_op_mant_lpi_1_dfm;
  wire [9:0] mul_nan_to_zero_op_mant_15_lpi_1_dfm;
  wire [9:0] mul_nan_to_zero_op_mant_14_lpi_1_dfm;
  wire [9:0] mul_nan_to_zero_op_mant_13_lpi_1_dfm;
  wire [9:0] mul_nan_to_zero_op_mant_12_lpi_1_dfm;
  wire [9:0] mul_nan_to_zero_op_mant_11_lpi_1_dfm;
  wire [9:0] mul_nan_to_zero_op_mant_10_lpi_1_dfm;
  wire [9:0] mul_nan_to_zero_op_mant_9_lpi_1_dfm;
  wire [9:0] mul_nan_to_zero_op_mant_8_lpi_1_dfm;
  wire [9:0] mul_nan_to_zero_op_mant_7_lpi_1_dfm;
  wire [9:0] mul_nan_to_zero_op_mant_6_lpi_1_dfm;
  wire [9:0] mul_nan_to_zero_op_mant_5_lpi_1_dfm;
  wire [9:0] mul_nan_to_zero_op_mant_4_lpi_1_dfm;
  wire [9:0] mul_nan_to_zero_op_mant_3_lpi_1_dfm;
  wire [9:0] mul_nan_to_zero_op_mant_2_lpi_1_dfm;
  wire [9:0] mul_nan_to_zero_op_mant_1_lpi_1_dfm;
  wire [47:0] FpMul_8U_23U_p_mant_p1_sva_mx1;
  wire [47:0] FpMul_8U_23U_p_mant_p1_15_sva_mx1;
  wire [47:0] FpMul_8U_23U_p_mant_p1_14_sva_mx1;
  wire [47:0] FpMul_8U_23U_p_mant_p1_13_sva_mx1;
  wire [47:0] FpMul_8U_23U_p_mant_p1_12_sva_mx1;
  wire [47:0] FpMul_8U_23U_p_mant_p1_11_sva_mx1;
  wire [47:0] FpMul_8U_23U_p_mant_p1_10_sva_mx1;
  wire [47:0] FpMul_8U_23U_p_mant_p1_9_sva_mx1;
  wire [47:0] FpMul_8U_23U_p_mant_p1_8_sva_mx1;
  wire [47:0] FpMul_8U_23U_p_mant_p1_7_sva_mx1;
  wire [47:0] FpMul_8U_23U_p_mant_p1_6_sva_mx1;
  wire [47:0] FpMul_8U_23U_p_mant_p1_5_sva_mx1;
  wire [47:0] FpMul_8U_23U_p_mant_p1_4_sva_mx1;
  wire [47:0] FpMul_8U_23U_p_mant_p1_3_sva_mx1;
  wire [47:0] FpMul_8U_23U_p_mant_p1_2_sva_mx1;
  wire [47:0] FpMul_8U_23U_p_mant_p1_1_sva_mx1;
  wire [4:0] mul_nan_to_zero_op_expo_lpi_1_dfm;
  wire [4:0] mul_nan_to_zero_op_expo_15_lpi_1_dfm;
  wire [4:0] mul_nan_to_zero_op_expo_14_lpi_1_dfm;
  wire [4:0] mul_nan_to_zero_op_expo_13_lpi_1_dfm;
  wire [4:0] mul_nan_to_zero_op_expo_12_lpi_1_dfm;
  wire [4:0] mul_nan_to_zero_op_expo_11_lpi_1_dfm;
  wire [4:0] mul_nan_to_zero_op_expo_10_lpi_1_dfm;
  wire [4:0] mul_nan_to_zero_op_expo_9_lpi_1_dfm;
  wire [4:0] mul_nan_to_zero_op_expo_8_lpi_1_dfm;
  wire [4:0] mul_nan_to_zero_op_expo_7_lpi_1_dfm;
  wire [4:0] mul_nan_to_zero_op_expo_6_lpi_1_dfm;
  wire [4:0] mul_nan_to_zero_op_expo_5_lpi_1_dfm;
  wire [4:0] mul_nan_to_zero_op_expo_4_lpi_1_dfm;
  wire [4:0] mul_nan_to_zero_op_expo_3_lpi_1_dfm;
  wire [4:0] mul_nan_to_zero_op_expo_2_lpi_1_dfm;
  wire [4:0] mul_nan_to_zero_op_expo_1_lpi_1_dfm;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_22_13_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_22_13_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_22_13_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_22_13_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_22_13_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_22_13_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_22_13_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_22_13_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_22_13_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_22_13_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_22_13_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_22_13_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_22_13_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_22_13_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_22_13_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_22_13_mx1;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_12_10_mx0w0;
  wire [2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_12_10_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_9_0_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_9_0_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_9_0_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_9_0_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_9_0_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_9_0_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_9_0_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_9_0_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_9_0_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_9_0_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_9_0_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_9_0_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_9_0_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_9_0_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_9_0_mx1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_9_0_mx1;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_3_2_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_3_2_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_3_2_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_3_2_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_3_2_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_3_2_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_3_2_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_3_2_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_3_2_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_3_2_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_3_2_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_3_2_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_3_2_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_3_2_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_3_2_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_3_2_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_1_0_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_1_0_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_1_0_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_1_0_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_1_0_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_1_0_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_1_0_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_1_0_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_1_0_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_1_0_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_1_0_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_1_0_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_1_0_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_1_0_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_1_0_mx0w0;
  wire [1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_1_0_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w0;
  wire and_2496_cse;
  wire and_2497_cse;
  wire or_4733_cse;
  wire chn_mul_out_and_cse;
  wire and_2488_cse;
  wire and_2489_cse;
  wire and_2481_cse;
  wire and_2482_cse;
  wire or_4729_cse;
  wire and_2473_cse;
  wire and_2474_cse;
  wire and_2466_cse;
  wire and_2467_cse;
  wire or_4725_cse;
  wire and_2458_cse;
  wire and_2459_cse;
  wire and_2451_cse;
  wire and_2452_cse;
  wire or_4721_cse;
  wire and_2443_cse;
  wire and_2444_cse;
  wire and_2436_cse;
  wire and_2437_cse;
  wire or_4717_cse;
  wire and_2428_cse;
  wire and_2429_cse;
  wire and_2421_cse;
  wire and_2422_cse;
  wire or_4713_cse;
  wire and_2413_cse;
  wire and_2414_cse;
  wire and_2406_cse;
  wire and_2407_cse;
  wire or_4709_cse;
  wire and_2398_cse;
  wire and_2399_cse;
  wire and_2391_cse;
  wire and_2392_cse;
  wire or_4705_cse;
  wire and_2383_cse;
  wire and_2384_cse;
  wire and_2376_cse;
  wire and_2377_cse;
  wire or_4701_cse;
  wire and_2368_cse;
  wire and_2369_cse;
  wire and_2361_cse;
  wire and_2362_cse;
  wire or_4697_cse;
  wire and_2353_cse;
  wire and_2354_cse;
  wire and_2346_cse;
  wire and_2347_cse;
  wire or_4693_cse;
  wire and_2338_cse;
  wire and_2339_cse;
  wire and_2331_cse;
  wire and_2332_cse;
  wire or_4689_cse;
  wire and_2323_cse;
  wire and_2324_cse;
  wire and_2316_cse;
  wire and_2317_cse;
  wire or_4685_cse;
  wire and_2308_cse;
  wire and_2309_cse;
  wire and_2301_cse;
  wire and_2302_cse;
  wire or_4681_cse;
  wire and_2293_cse;
  wire and_2294_cse;
  wire and_2286_cse;
  wire and_2287_cse;
  wire or_4677_cse;
  wire and_2278_cse;
  wire and_2279_cse;
  wire and_2271_cse;
  wire and_2272_cse;
  wire or_4673_cse;
  wire and_2263_cse;
  wire and_2264_cse;
  reg reg_cfg_mul_src_rsc_triosy_obj_ld_core_psct_cse;
  wire or_90_cse;
  wire cfg_mul_op_and_cse;
  wire or_309_cse;
  wire nor_53_cse;
  wire nor_129_cse;
  wire nor_1490_cse;
  wire nor_145_cse;
  wire nor_161_cse;
  wire nor_193_cse;
  wire nor_209_cse;
  wire nor_225_cse;
  wire nor_241_cse;
  wire nor_257_cse;
  wire nor_273_cse;
  wire nor_283_cse;
  wire nor_336_cse;
  wire nor_332_cse;
  wire nor_352_cse;
  wire nor_368_cse;
  reg reg_chn_mul_out_rsci_ld_core_psct_cse;
  wire nor_872_cse;
  wire nor_133_cse;
  wire FpMul_8U_23U_p_expo_and_cse;
  wire FpMantRNE_48U_24U_else_and_cse;
  wire nor_149_cse;
  wire FpMul_8U_23U_p_expo_and_1_cse;
  wire FpMantRNE_48U_24U_else_and_2_cse;
  wire nor_165_cse;
  wire FpMantRNE_48U_24U_else_carry_and_2_cse;
  wire FpMul_8U_23U_p_expo_and_2_cse;
  wire nor_181_cse;
  wire FpMul_8U_23U_p_expo_and_3_cse;
  wire FpMantRNE_48U_24U_else_and_6_cse;
  wire nor_197_cse;
  wire FpMul_8U_23U_p_expo_and_4_cse;
  wire FpMantRNE_48U_24U_else_and_8_cse;
  wire FpMul_8U_23U_p_expo_and_5_cse;
  wire FpMantRNE_48U_24U_else_and_10_cse;
  wire nor_229_cse;
  wire FpMantRNE_48U_24U_else_carry_and_6_cse;
  wire FpMul_8U_23U_p_expo_and_6_cse;
  wire nor_245_cse;
  wire FpMul_8U_23U_p_expo_and_7_cse;
  wire FpMantRNE_48U_24U_else_and_14_cse;
  wire nor_261_cse;
  wire FpMul_8U_23U_p_expo_and_8_cse;
  wire FpMantRNE_48U_24U_else_and_16_cse;
  wire FpMul_8U_23U_p_expo_and_9_cse;
  wire FpMantRNE_48U_24U_else_and_18_cse;
  wire FpMul_8U_23U_p_expo_and_10_cse;
  wire FpMantRNE_48U_24U_else_and_20_cse;
  wire nor_309_cse;
  wire FpMul_8U_23U_p_expo_and_11_cse;
  wire FpMantRNE_48U_24U_else_and_22_cse;
  wire nor_325_cse;
  wire FpMul_8U_23U_p_expo_and_12_cse;
  wire FpMantRNE_48U_24U_else_and_24_cse;
  wire nor_340_cse;
  wire FpMul_8U_23U_p_expo_and_13_cse;
  wire FpMantRNE_48U_24U_else_and_26_cse;
  wire nor_356_cse;
  wire FpMul_8U_23U_p_expo_and_14_cse;
  wire FpMantRNE_48U_24U_else_and_28_cse;
  wire FpMantRNE_48U_24U_else_carry_and_15_cse;
  wire nor_372_cse;
  wire FpMul_8U_23U_p_expo_and_15_cse;
  wire or_2577_cse;
  wire IsZero_8U_23U_aelse_and_cse;
  wire or_2608_cse;
  wire or_2575_cse;
  wire FpMul_8U_23U_else_2_if_and_cse;
  wire or_2631_cse;
  wire or_2664_cse;
  wire or_2675_cse;
  wire or_414_cse;
  wire IsZero_8U_23U_1_aelse_and_cse;
  wire or_2698_cse;
  wire or_2711_cse;
  wire or_2722_cse;
  wire or_2745_cse;
  wire or_517_cse;
  wire or_2774_cse;
  wire or_2787_cse;
  wire or_2798_cse;
  wire or_616_cse;
  wire or_2823_cse;
  wire or_2834_cse;
  wire or_2865_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_3_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_6_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_9_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_12_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_15_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_18_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_21_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_24_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_27_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_30_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_33_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_36_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_39_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_42_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_45_cse;
  wire mul_loop_mul_if_aelse_and_cse;
  wire and_2130_cse;
  wire and_384_cse;
  wire nor_749_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_3_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_6_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_9_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_12_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_15_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_18_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_21_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_24_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_27_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_30_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_33_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_36_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_39_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_42_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_45_cse;
  wire IsZero_8U_23U_aelse_and_16_cse;
  wire IsZero_8U_23U_aelse_and_17_cse;
  wire IsZero_8U_23U_aelse_and_18_cse;
  wire IsZero_8U_23U_aelse_and_19_cse;
  wire IsZero_8U_23U_aelse_and_20_cse;
  wire IsZero_8U_23U_aelse_and_21_cse;
  wire IsZero_8U_23U_aelse_and_22_cse;
  wire IsZero_8U_23U_aelse_and_23_cse;
  wire IsZero_8U_23U_aelse_and_24_cse;
  wire IsZero_8U_23U_aelse_and_25_cse;
  wire IsZero_8U_23U_aelse_and_26_cse;
  wire IsZero_8U_23U_aelse_and_27_cse;
  wire IsZero_8U_23U_aelse_and_28_cse;
  wire IsZero_8U_23U_aelse_and_29_cse;
  wire IsZero_8U_23U_aelse_and_30_cse;
  wire IsZero_8U_23U_aelse_and_31_cse;
  wire or_2885_cse;
  wire or_662_cse;
  wire or_639_cse;
  wire or_593_cse;
  wire or_570_cse;
  wire or_2742_cse;
  wire or_461_cse;
  wire or_438_cse;
  wire or_386_cse;
  wire or_363_cse;
  wire or_2628_cse;
  wire or_312_cse;
  wire nor_44_cse;
  wire nor_42_cse;
  wire nor_40_cse;
  wire nor_39_cse;
  wire nor_37_cse;
  wire nor_36_cse;
  wire nor_35_cse;
  wire nor_34_cse;
  wire nor_32_cse;
  wire nor_30_cse;
  wire nor_29_cse;
  wire nor_28_cse;
  wire nor_26_cse;
  wire nor_25_cse;
  wire nor_23_cse;
  wire nor_21_cse;
  wire or_1253_cse;
  wire or_2342_cse;
  wire or_2386_cse;
  wire or_1898_cse;
  wire or_1981_cse;
  wire or_4649_cse;
  wire or_2576_cse;
  wire nor_50_cse;
  wire or_4383_cse;
  wire or_2607_cse;
  wire nor_55_cse;
  wire or_4384_cse;
  wire or_2630_cse;
  wire nor_59_cse;
  wire or_4385_cse;
  wire nor_177_cse;
  wire nor_64_cse;
  wire nor_69_cse;
  wire or_4387_cse;
  wire nor_73_cse;
  wire nor_78_cse;
  wire or_4389_cse;
  wire or_2721_cse;
  wire nor_83_cse;
  wire or_4390_cse;
  wire nor_87_cse;
  wire or_4391_cse;
  wire or_2767_cse;
  wire nor_91_cse;
  wire nor_289_cse;
  wire nor_95_cse;
  wire or_1819_cse;
  wire nor_305_cse;
  wire nor_100_cse;
  wire nor_321_cse;
  wire or_2797_cse;
  wire nor_105_cse;
  wire nor_110_cse;
  wire or_4398_cse;
  wire or_2833_cse;
  wire nor_115_cse;
  wire or_4399_cse;
  wire or_2864_cse;
  wire nor_120_cse;
  wire or_4400_cse;
  wire nor_1383_cse;
  wire nor_1351_cse;
  wire nor_1317_cse;
  wire nor_1287_cse;
  wire nor_1255_cse;
  wire nor_1221_cse;
  wire nor_213_cse;
  wire nor_1187_cse;
  wire nor_1155_cse;
  wire nor_1123_cse;
  wire nor_1090_cse;
  wire nor_277_cse;
  wire nor_1103_cse;
  wire nor_1070_cse;
  wire nor_1059_cse;
  wire nor_1037_cse;
  wire nor_1026_cse;
  wire nor_1004_cse;
  wire nor_993_cse;
  wire nor_972_cse;
  wire nor_935_cse;
  wire nor_920_cse;
  wire nor_898_cse;
  wire nor_885_cse;
  wire or_378_cse;
  wire or_430_cse;
  wire or_453_cse;
  wire or_533_cse;
  wire or_562_cse;
  wire or_585_cse;
  wire or_631_cse;
  wire or_70_cse;
  wire or_75_cse;
  wire or_76_cse;
  wire or_77_cse;
  wire or_78_cse;
  wire or_79_cse;
  wire or_80_cse;
  wire or_81_cse;
  wire or_82_cse;
  wire or_83_cse;
  wire or_84_cse;
  wire or_85_cse;
  wire or_86_cse;
  wire or_87_cse;
  wire or_88_cse;
  wire or_89_cse;
  wire not_tmp_1326;
  wire not_tmp_1344;
  wire not_tmp_1362;
  wire not_tmp_1380;
  wire not_tmp_1398;
  wire not_tmp_1416;
  wire not_tmp_1434;
  wire not_tmp_1452;
  wire not_tmp_1470;
  wire not_tmp_1488;
  wire not_tmp_1506;
  wire not_tmp_1524;
  wire not_tmp_1542;
  wire not_tmp_1578;
  wire not_tmp_1596;
  wire and_1108_rgt;
  wire and_1111_rgt;
  wire and_1112_rgt;
  wire and_1117_rgt;
  wire and_1120_rgt;
  wire and_1121_rgt;
  wire and_1126_rgt;
  wire and_1129_rgt;
  wire and_1130_rgt;
  wire and_1135_rgt;
  wire and_1138_rgt;
  wire and_1139_rgt;
  wire and_1144_rgt;
  wire and_1147_rgt;
  wire and_1148_rgt;
  wire and_1153_rgt;
  wire and_1156_rgt;
  wire and_1157_rgt;
  wire and_1162_rgt;
  wire and_1165_rgt;
  wire and_1166_rgt;
  wire and_1171_rgt;
  wire and_1174_rgt;
  wire and_1175_rgt;
  wire and_1180_rgt;
  wire and_1183_rgt;
  wire and_1184_rgt;
  wire and_1189_rgt;
  wire and_1192_rgt;
  wire and_1193_rgt;
  wire and_1198_rgt;
  wire and_1201_rgt;
  wire and_1202_rgt;
  wire and_1207_rgt;
  wire and_1210_rgt;
  wire and_1211_rgt;
  wire and_1216_rgt;
  wire and_1219_rgt;
  wire and_1220_rgt;
  wire and_1225_rgt;
  wire and_1228_rgt;
  wire and_1229_rgt;
  wire and_1234_rgt;
  wire and_1237_rgt;
  wire and_1238_rgt;
  wire and_1243_rgt;
  wire and_1246_rgt;
  wire and_1247_rgt;
  wire and_1252_rgt;
  wire and_1257_rgt;
  wire and_1262_rgt;
  wire and_1267_rgt;
  wire and_1272_rgt;
  wire and_1277_rgt;
  wire and_1282_rgt;
  wire and_1287_rgt;
  wire and_1292_rgt;
  wire and_1297_rgt;
  wire and_1302_rgt;
  wire and_1307_rgt;
  wire and_1312_rgt;
  wire and_1317_rgt;
  wire and_1322_rgt;
  wire and_1327_rgt;
  wire [7:0] FpMul_8U_23U_p_expo_mux1h_1_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_1_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_1_2_itm;
  wire [7:0] FpMul_8U_23U_p_expo_mux1h_3_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_2_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_2_2_itm;
  wire [7:0] FpMul_8U_23U_p_expo_mux1h_5_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_3_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_3_2_itm;
  wire [7:0] FpMul_8U_23U_p_expo_mux1h_7_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_4_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_4_2_itm;
  wire [7:0] FpMul_8U_23U_p_expo_mux1h_9_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_5_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_5_2_itm;
  wire [7:0] FpMul_8U_23U_p_expo_mux1h_11_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_6_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_6_2_itm;
  wire [7:0] FpMul_8U_23U_p_expo_mux1h_13_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_7_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_7_2_itm;
  wire [7:0] FpMul_8U_23U_p_expo_mux1h_15_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_8_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_8_2_itm;
  wire [7:0] FpMul_8U_23U_p_expo_mux1h_17_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_9_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_9_2_itm;
  wire [7:0] FpMul_8U_23U_p_expo_mux1h_19_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_10_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_10_2_itm;
  wire [7:0] FpMul_8U_23U_p_expo_mux1h_21_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_11_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_11_2_itm;
  wire [7:0] FpMul_8U_23U_p_expo_mux1h_23_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_12_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_12_2_itm;
  wire [7:0] FpMul_8U_23U_p_expo_mux1h_25_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_13_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_13_2_itm;
  wire [7:0] FpMul_8U_23U_p_expo_mux1h_27_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_14_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_14_2_itm;
  wire [7:0] FpMul_8U_23U_p_expo_mux1h_29_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_15_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_15_2_itm;
  wire [7:0] FpMul_8U_23U_p_expo_mux1h_31_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_itm;
  reg [3:0] reg_FpMul_8U_23U_p_expo_2_itm_1;
  wire mux_156_itm;
  wire mux_157_itm;
  wire mux_158_itm;
  wire mux_159_itm;
  wire mux_160_itm;
  wire mux_161_itm;
  wire mux_162_itm;
  wire mux_163_itm;
  wire mux_164_itm;
  wire mux_165_itm;
  wire mux_166_itm;
  wire mux_167_itm;
  wire mux_168_itm;
  wire mux_169_itm;
  wire mux_170_itm;
  wire mux_171_itm;
  wire mux_187_itm;
  wire mux_202_itm;
  wire mux_216_itm;
  wire mux_230_itm;
  wire mux_245_itm;
  wire mux_259_itm;
  wire mux_273_itm;
  wire mux_288_itm;
  wire mux_303_itm;
  wire mux_318_itm;
  wire mux_332_itm;
  wire mux_346_itm;
  wire mux_360_itm;
  wire mux_374_itm;
  wire mux_388_itm;
  wire mux_403_itm;
  wire mux_522_itm;
  wire mux_523_itm;
  wire mux_546_itm;
  wire mux_547_itm;
  wire mux_570_itm;
  wire mux_571_itm;
  wire mux_596_itm;
  wire mux_597_itm;
  wire mux_620_itm;
  wire mux_621_itm;
  wire mux_644_itm;
  wire mux_645_itm;
  wire mux_668_itm;
  wire mux_669_itm;
  wire mux_692_itm;
  wire mux_693_itm;
  wire mux_716_itm;
  wire mux_717_itm;
  wire mux_740_itm;
  wire mux_741_itm;
  wire mux_767_itm;
  wire mux_793_itm;
  wire mux_794_itm;
  wire mux_820_itm;
  wire mux_821_itm;
  wire mux_845_itm;
  wire mux_846_itm;
  wire mux_870_itm;
  wire mux_871_itm;
  wire mux_895_itm;
  wire mux_896_itm;
  wire chn_mul_in_rsci_ld_core_psct_mx0c0;
  wire chn_mul_op_rsci_ld_core_psct_mx0c1;
  wire mul_loop_mul_1_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
  wire mul_loop_mul_2_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
  wire mul_loop_mul_3_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
  wire mul_loop_mul_4_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
  wire mul_loop_mul_5_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
  wire mul_loop_mul_6_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
  wire mul_loop_mul_7_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
  wire mul_loop_mul_8_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
  wire mul_loop_mul_9_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
  wire mul_loop_mul_10_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
  wire mul_loop_mul_11_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
  wire mul_loop_mul_12_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
  wire mul_loop_mul_13_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
  wire mul_loop_mul_14_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
  wire mul_loop_mul_15_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
  wire mul_loop_mul_16_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
  wire main_stage_v_1_mx0c1;
  wire cfg_mul_src_1_sva_st_1_mx0c1;
  wire main_stage_v_2_mx0c1;
  wire FpMul_8U_23U_lor_6_lpi_1_dfm_mx0w0;
  wire FpMul_8U_23U_lor_8_lpi_1_dfm_mx0w0;
  wire FpMul_8U_23U_lor_9_lpi_1_dfm_mx0w0;
  wire FpMul_8U_23U_lor_12_lpi_1_dfm_mx0w0;
  wire FpMul_8U_23U_lor_13_lpi_1_dfm_mx0w0;
  wire FpMul_8U_23U_lor_14_lpi_1_dfm_mx0w0;
  wire FpMul_8U_23U_lor_16_lpi_1_dfm_mx0w0;
  wire main_stage_v_3_mx0c1;
  wire main_stage_v_4_mx0c1;
  wire [7:0] FpMul_8U_23U_p_expo_1_sva_1_mx0w0;
  wire [8:0] nl_FpMul_8U_23U_p_expo_1_sva_1_mx0w0;
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_mx0w0;
  wire mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs_mx0w0;
  wire FpMul_8U_23U_FpMul_8U_23U_and_itm_mx0w0;
  wire [7:0] FpMul_8U_23U_p_expo_2_sva_1_mx0w0;
  wire [8:0] nl_FpMul_8U_23U_p_expo_2_sva_1_mx0w0;
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_mx0w0;
  wire mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs_mx0w0;
  wire FpMul_8U_23U_FpMul_8U_23U_and_64_itm_mx0w0;
  wire [7:0] FpMul_8U_23U_p_expo_3_sva_1_mx0w0;
  wire [8:0] nl_FpMul_8U_23U_p_expo_3_sva_1_mx0w0;
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_mx0w0;
  wire mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs_mx0w0;
  wire FpMul_8U_23U_FpMul_8U_23U_and_65_itm_mx0w0;
  wire [7:0] FpMul_8U_23U_p_expo_4_sva_1_mx0w0;
  wire [8:0] nl_FpMul_8U_23U_p_expo_4_sva_1_mx0w0;
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_mx0w0;
  wire mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs_mx0w0;
  wire FpMul_8U_23U_FpMul_8U_23U_and_66_itm_mx0w0;
  wire [7:0] FpMul_8U_23U_p_expo_5_sva_1_mx0w0;
  wire [8:0] nl_FpMul_8U_23U_p_expo_5_sva_1_mx0w0;
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_4_itm_mx0w0;
  wire mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs_mx0w0;
  wire FpMul_8U_23U_FpMul_8U_23U_and_67_itm_mx0w0;
  wire [7:0] FpMul_8U_23U_p_expo_6_sva_1_mx0w0;
  wire [8:0] nl_FpMul_8U_23U_p_expo_6_sva_1_mx0w0;
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_5_itm_mx0w0;
  wire mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs_mx0w0;
  wire FpMul_8U_23U_FpMul_8U_23U_and_68_itm_mx0w0;
  wire [7:0] FpMul_8U_23U_p_expo_7_sva_1_mx0w0;
  wire [8:0] nl_FpMul_8U_23U_p_expo_7_sva_1_mx0w0;
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_6_itm_mx0w0;
  wire mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs_mx0w0;
  wire FpMul_8U_23U_FpMul_8U_23U_and_69_itm_mx0w0;
  wire [7:0] FpMul_8U_23U_p_expo_8_sva_1_mx0w0;
  wire [8:0] nl_FpMul_8U_23U_p_expo_8_sva_1_mx0w0;
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_7_itm_mx0w0;
  wire mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs_mx0w0;
  wire FpMul_8U_23U_FpMul_8U_23U_and_70_itm_mx0w0;
  wire [7:0] FpMul_8U_23U_p_expo_9_sva_1_mx0w0;
  wire [8:0] nl_FpMul_8U_23U_p_expo_9_sva_1_mx0w0;
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_8_itm_mx0w0;
  wire mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs_mx0w0;
  wire FpMul_8U_23U_FpMul_8U_23U_and_71_itm_mx0w0;
  wire [7:0] FpMul_8U_23U_p_expo_10_sva_1_mx0w0;
  wire [8:0] nl_FpMul_8U_23U_p_expo_10_sva_1_mx0w0;
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_9_itm_mx0w0;
  wire mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs_mx0w0;
  wire FpMul_8U_23U_FpMul_8U_23U_and_72_itm_mx0w0;
  wire [7:0] FpMul_8U_23U_p_expo_11_sva_1_mx0w0;
  wire [8:0] nl_FpMul_8U_23U_p_expo_11_sva_1_mx0w0;
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_10_itm_mx0w0;
  wire mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs_mx0w0;
  wire FpMul_8U_23U_FpMul_8U_23U_and_73_itm_mx0w0;
  wire [7:0] FpMul_8U_23U_p_expo_12_sva_1_mx0w0;
  wire [8:0] nl_FpMul_8U_23U_p_expo_12_sva_1_mx0w0;
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_11_itm_mx0w0;
  wire mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs_mx0w0;
  wire FpMul_8U_23U_FpMul_8U_23U_and_74_itm_mx0w0;
  wire [7:0] FpMul_8U_23U_p_expo_13_sva_1_mx0w0;
  wire [8:0] nl_FpMul_8U_23U_p_expo_13_sva_1_mx0w0;
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_12_itm_mx0w0;
  wire mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs_mx0w0;
  wire FpMul_8U_23U_FpMul_8U_23U_and_75_itm_mx0w0;
  wire [7:0] FpMul_8U_23U_p_expo_14_sva_1_mx0w0;
  wire [8:0] nl_FpMul_8U_23U_p_expo_14_sva_1_mx0w0;
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_13_itm_mx0w0;
  wire mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs_mx0w0;
  wire FpMul_8U_23U_FpMul_8U_23U_and_76_itm_mx0w0;
  wire [7:0] FpMul_8U_23U_p_expo_15_sva_1_mx0w0;
  wire [8:0] nl_FpMul_8U_23U_p_expo_15_sva_1_mx0w0;
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_14_itm_mx0w0;
  wire mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs_mx0w0;
  wire FpMul_8U_23U_FpMul_8U_23U_and_77_itm_mx0w0;
  wire [7:0] FpMul_8U_23U_p_expo_sva_1_mx0w0;
  wire [8:0] nl_FpMul_8U_23U_p_expo_sva_1_mx0w0;
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_15_itm_mx0w0;
  wire mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs_mx0w0;
  wire FpMul_8U_23U_FpMul_8U_23U_and_78_itm_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_65_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_64_mx0w1;
  wire IsZero_8U_23U_1_land_1_lpi_1_dfm_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_68_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_67_mx0w1;
  wire IsZero_8U_23U_1_land_2_lpi_1_dfm_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_71_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_70_mx0w1;
  wire IsZero_8U_23U_1_land_3_lpi_1_dfm_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_74_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_73_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_77_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_76_mx0w1;
  wire IsZero_8U_23U_1_land_5_lpi_1_dfm_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_80_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_79_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_83_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_82_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_86_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_85_mx0w1;
  wire IsZero_8U_23U_1_land_8_lpi_1_dfm_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_89_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_88_mx0w1;
  wire IsZero_8U_23U_1_land_9_lpi_1_dfm_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_92_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_91_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_95_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_94_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_98_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_97_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_101_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_100_mx0w1;
  wire IsZero_8U_23U_1_land_13_lpi_1_dfm_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_104_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_103_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_107_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_106_mx0w1;
  wire IsZero_8U_23U_1_land_15_lpi_1_dfm_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_110_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_109_mx0w1;
  wire IsZero_8U_23U_1_land_lpi_1_dfm_mx0w0;
  wire IsZero_8U_23U_land_1_lpi_1_dfm_mx0w0;
  wire IsZero_8U_23U_land_2_lpi_1_dfm_mx0w0;
  wire IsZero_8U_23U_land_3_lpi_1_dfm_mx0w0;
  wire IsZero_8U_23U_land_4_lpi_1_dfm_mx0w0;
  wire IsZero_8U_23U_land_5_lpi_1_dfm_mx0w0;
  wire IsZero_8U_23U_land_6_lpi_1_dfm_mx0w0;
  wire IsZero_8U_23U_land_7_lpi_1_dfm_mx0w0;
  wire IsZero_8U_23U_land_8_lpi_1_dfm_mx0w0;
  wire IsZero_8U_23U_land_9_lpi_1_dfm_mx0w0;
  wire IsZero_8U_23U_land_10_lpi_1_dfm_mx0w0;
  wire IsZero_8U_23U_land_11_lpi_1_dfm_mx0w0;
  wire IsZero_8U_23U_land_12_lpi_1_dfm_mx0w0;
  wire IsZero_8U_23U_land_13_lpi_1_dfm_mx0w0;
  wire IsZero_8U_23U_land_14_lpi_1_dfm_mx0w0;
  wire IsZero_8U_23U_land_15_lpi_1_dfm_mx0w0;
  wire IsZero_8U_23U_land_lpi_1_dfm_mx0w0;
  wire FpMul_8U_23U_else_5_mux_60_mx0w1;
  wire FpMul_8U_23U_else_5_mux_56_mx0w1;
  wire FpMul_8U_23U_else_5_mux_52_mx0w1;
  wire FpMul_8U_23U_else_5_mux_48_mx0w1;
  wire FpMul_8U_23U_else_5_mux_44_mx0w1;
  wire FpMul_8U_23U_else_5_mux_40_mx0w1;
  wire FpMul_8U_23U_lor_27_lpi_1_dfm_mx0w0;
  wire FpMul_8U_23U_else_5_mux_36_mx0w1;
  wire FpMul_8U_23U_lor_26_lpi_1_dfm_mx0w0;
  wire FpMul_8U_23U_else_5_mux_32_mx0w1;
  wire FpMul_8U_23U_else_5_mux_28_mx0w1;
  wire FpMul_8U_23U_else_5_mux_24_mx0w1;
  wire FpMul_8U_23U_else_5_mux_20_mx0w1;
  wire FpMul_8U_23U_lor_22_lpi_1_dfm_mx0w0;
  wire FpMul_8U_23U_else_5_mux_16_mx0w1;
  wire FpMul_8U_23U_else_5_mux_12_mx0w1;
  wire FpMul_8U_23U_else_5_mux_8_mx0w1;
  wire FpMul_8U_23U_else_5_mux_4_mx0w1;
  wire FpMul_8U_23U_else_5_mux_mx0w1;
  wire FpMul_8U_23U_mux_12_itm_mx0c1;
  wire FpMul_8U_23U_mux_28_itm_mx0c1;
  wire FpMul_8U_23U_mux_44_itm_mx0c1;
  wire FpMul_8U_23U_mux_60_itm_mx0c1;
  wire FpMul_8U_23U_mux_76_itm_mx0c1;
  wire FpMul_8U_23U_mux_92_itm_mx0c1;
  wire FpMul_8U_23U_mux_108_itm_mx0c1;
  wire FpMul_8U_23U_mux_124_itm_mx0c1;
  wire FpMul_8U_23U_mux_140_itm_mx0c1;
  wire FpMul_8U_23U_mux_156_itm_mx0c1;
  wire FpMul_8U_23U_mux_172_itm_mx0c1;
  wire FpMul_8U_23U_mux_188_itm_mx0c1;
  wire FpMul_8U_23U_mux_204_itm_mx0c1;
  wire FpMul_8U_23U_mux_220_itm_mx0c1;
  wire FpMul_8U_23U_mux_236_itm_mx0c1;
  wire FpMul_8U_23U_mux_252_itm_mx0c1;
  wire IsNaN_8U_23U_land_1_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_land_2_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_land_3_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_land_4_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_land_5_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_land_6_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_land_7_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_land_8_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_land_9_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_land_10_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_land_11_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_land_12_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_land_13_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_land_14_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_land_15_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_land_lpi_1_dfm_mx0w0;
  wire [9:0] else_MulOp_data_0_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_MulOp_data_1_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_MulOp_data_2_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_MulOp_data_3_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_MulOp_data_4_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_MulOp_data_5_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_MulOp_data_6_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_MulOp_data_7_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_MulOp_data_8_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_MulOp_data_9_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_MulOp_data_10_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_MulOp_data_11_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_MulOp_data_12_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_MulOp_data_13_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_MulOp_data_14_9_0_lpi_1_dfm_mx0;
  wire [9:0] else_MulOp_data_15_9_0_lpi_1_dfm_mx0;
  wire [7:0] FpMul_8U_23U_p_expo_1_lpi_1_dfm_1_mx0;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_1_lpi_1_dfm;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_1_sva;
  wire [23:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_1_sva;
  wire FpMul_8U_23U_lor_33_lpi_1_dfm;
  wire [7:0] FpMul_8U_23U_p_expo_2_lpi_1_dfm_1_mx0;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_2_lpi_1_dfm;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_2_sva;
  wire [23:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_2_sva;
  wire FpMul_8U_23U_lor_34_lpi_1_dfm;
  wire [7:0] FpMul_8U_23U_p_expo_3_lpi_1_dfm_1_mx0;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_3_lpi_1_dfm;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_3_sva;
  wire [23:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_3_sva;
  wire FpMul_8U_23U_lor_35_lpi_1_dfm;
  wire [7:0] FpMul_8U_23U_p_expo_4_lpi_1_dfm_1_mx0;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_4_lpi_1_dfm;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_4_sva;
  wire [23:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_4_sva;
  wire FpMul_8U_23U_lor_36_lpi_1_dfm;
  wire [7:0] FpMul_8U_23U_p_expo_5_lpi_1_dfm_1_mx0;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_5_lpi_1_dfm;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_5_sva;
  wire [23:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_5_sva;
  wire FpMul_8U_23U_lor_37_lpi_1_dfm;
  wire [7:0] FpMul_8U_23U_p_expo_6_lpi_1_dfm_1_mx0;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_6_lpi_1_dfm;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_6_sva;
  wire [23:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_6_sva;
  wire FpMul_8U_23U_lor_38_lpi_1_dfm;
  wire [7:0] FpMul_8U_23U_p_expo_7_lpi_1_dfm_1_mx0;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_7_lpi_1_dfm;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_7_sva;
  wire [23:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_7_sva;
  wire FpMul_8U_23U_lor_39_lpi_1_dfm;
  wire [7:0] FpMul_8U_23U_p_expo_8_lpi_1_dfm_1_mx0;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_8_lpi_1_dfm;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_8_sva;
  wire [23:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_8_sva;
  wire FpMul_8U_23U_lor_40_lpi_1_dfm;
  wire [7:0] FpMul_8U_23U_p_expo_9_lpi_1_dfm_1_mx0;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_9_lpi_1_dfm;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_9_sva;
  wire [23:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_9_sva;
  wire FpMul_8U_23U_lor_41_lpi_1_dfm;
  wire [7:0] FpMul_8U_23U_p_expo_10_lpi_1_dfm_1_mx0;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_10_lpi_1_dfm;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_10_sva;
  wire [23:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_10_sva;
  wire FpMul_8U_23U_lor_42_lpi_1_dfm;
  wire [7:0] FpMul_8U_23U_p_expo_11_lpi_1_dfm_1_mx0;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_11_lpi_1_dfm;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_11_sva;
  wire [23:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_11_sva;
  wire FpMul_8U_23U_lor_43_lpi_1_dfm;
  wire [7:0] FpMul_8U_23U_p_expo_12_lpi_1_dfm_1_mx0;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_12_lpi_1_dfm;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_12_sva;
  wire [23:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_12_sva;
  wire FpMul_8U_23U_lor_44_lpi_1_dfm;
  wire [7:0] FpMul_8U_23U_p_expo_13_lpi_1_dfm_1_mx0;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_13_lpi_1_dfm;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_13_sva;
  wire [23:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_13_sva;
  wire FpMul_8U_23U_lor_45_lpi_1_dfm;
  wire [7:0] FpMul_8U_23U_p_expo_14_lpi_1_dfm_1_mx0;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_14_lpi_1_dfm;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_14_sva;
  wire [23:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_14_sva;
  wire FpMul_8U_23U_lor_46_lpi_1_dfm;
  wire [7:0] FpMul_8U_23U_p_expo_15_lpi_1_dfm_1_mx0;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_15_lpi_1_dfm;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_15_sva;
  wire [23:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_15_sva;
  wire FpMul_8U_23U_lor_47_lpi_1_dfm;
  wire [7:0] FpMul_8U_23U_p_expo_lpi_1_dfm_1_mx0;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_lpi_1_dfm;
  wire [22:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_sva;
  wire [23:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_sva;
  wire FpMul_8U_23U_lor_2_lpi_1_dfm;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_sva_1;
  wire [4:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_sva_1;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_sva_2;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_1_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_1_sva;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_ssc;
  wire IsNaN_5U_23U_land_1_lpi_1_dfm;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_sva_1;
  wire [4:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_sva_1;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_sva_2;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_2_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_2_sva;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_ssc;
  wire IsNaN_5U_23U_land_2_lpi_1_dfm;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_sva_1;
  wire [4:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_sva_1;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_sva_2;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_3_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_3_sva;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_ssc;
  wire IsNaN_5U_23U_land_3_lpi_1_dfm;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_sva_1;
  wire [4:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_sva_1;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_sva_2;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_4_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_4_sva;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_ssc;
  wire IsNaN_5U_23U_land_4_lpi_1_dfm;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_sva_1;
  wire [4:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_sva_1;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_sva_2;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_5_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_5_sva;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_ssc;
  wire IsNaN_5U_23U_land_5_lpi_1_dfm;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_sva_1;
  wire [4:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_sva_1;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_sva_2;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_6_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_6_sva;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_ssc;
  wire IsNaN_5U_23U_land_6_lpi_1_dfm;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_sva_1;
  wire [4:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_sva_1;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_sva_2;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_7_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_7_sva;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_ssc;
  wire IsNaN_5U_23U_land_7_lpi_1_dfm;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_sva_1;
  wire [4:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_sva_1;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_sva_2;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_8_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_8_sva;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_ssc;
  wire IsNaN_5U_23U_land_8_lpi_1_dfm;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_sva_1;
  wire [4:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_sva_1;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_sva_2;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_9_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_9_sva;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_16_ssc;
  wire IsNaN_5U_23U_land_9_lpi_1_dfm;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_sva_1;
  wire [4:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_sva_1;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_sva_2;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_10_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_10_sva;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_18_ssc;
  wire IsNaN_5U_23U_land_10_lpi_1_dfm;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_sva_1;
  wire [4:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_sva_1;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_sva_2;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_11_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_11_sva;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_20_ssc;
  wire IsNaN_5U_23U_land_11_lpi_1_dfm;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_sva_1;
  wire [4:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_sva_1;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_sva_2;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_12_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_12_sva;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_22_ssc;
  wire IsNaN_5U_23U_land_12_lpi_1_dfm;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_sva_1;
  wire [4:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_sva_1;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_sva_2;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_13_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_13_sva;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_24_ssc;
  wire IsNaN_5U_23U_land_13_lpi_1_dfm;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_sva_1;
  wire [4:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_sva_1;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_sva_2;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_14_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_14_sva;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_26_ssc;
  wire IsNaN_5U_23U_land_14_lpi_1_dfm;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_sva_1;
  wire [4:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_sva_1;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_sva_2;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_15_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_15_sva;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_28_ssc;
  wire IsNaN_5U_23U_land_15_lpi_1_dfm;
  wire [3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_sva_1;
  wire [4:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_sva_1;
  wire [22:0] FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_sva_2;
  wire [5:0] FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_sva;
  wire [6:0] nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_sva;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_30_ssc;
  wire IsNaN_5U_23U_land_lpi_1_dfm;
  wire else_MulOp_data_0_15_lpi_1_dfm_mx0;
  wire else_MulOp_data_1_15_lpi_1_dfm_mx0;
  wire else_MulOp_data_2_15_lpi_1_dfm_mx0;
  wire else_MulOp_data_3_15_lpi_1_dfm_mx0;
  wire else_MulOp_data_4_15_lpi_1_dfm_mx0;
  wire else_MulOp_data_5_15_lpi_1_dfm_mx0;
  wire else_MulOp_data_6_15_lpi_1_dfm_mx0;
  wire else_MulOp_data_7_15_lpi_1_dfm_mx0;
  wire else_MulOp_data_8_15_lpi_1_dfm_mx0;
  wire else_MulOp_data_9_15_lpi_1_dfm_mx0;
  wire else_MulOp_data_10_15_lpi_1_dfm_mx0;
  wire else_MulOp_data_11_15_lpi_1_dfm_mx0;
  wire else_MulOp_data_12_15_lpi_1_dfm_mx0;
  wire else_MulOp_data_13_15_lpi_1_dfm_mx0;
  wire else_MulOp_data_14_15_lpi_1_dfm_mx0;
  wire else_MulOp_data_15_15_lpi_1_dfm_mx0;
  wire asn_1163;
  wire asn_1165;
  wire asn_1173;
  wire asn_1175;
  wire asn_1183;
  wire asn_1185;
  wire asn_1193;
  wire asn_1195;
  wire asn_1203;
  wire asn_1205;
  wire asn_1213;
  wire asn_1215;
  wire asn_1223;
  wire asn_1225;
  wire asn_1233;
  wire asn_1235;
  wire asn_1243;
  wire asn_1245;
  wire asn_1253;
  wire asn_1255;
  wire asn_1263;
  wire asn_1265;
  wire asn_1273;
  wire asn_1275;
  wire asn_1283;
  wire asn_1285;
  wire asn_1293;
  wire asn_1295;
  wire asn_1303;
  wire asn_1305;
  wire asn_1313;
  wire asn_1315;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_exs_261_0;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_exs_267_0;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_exs_273_0;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_exs_279_0;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_exs_285_0;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_exs_291_0;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_exs_297_0;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_exs_303_0;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_exs_309_0;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_exs_315_0;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_exs_321_0;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_exs_327_0;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_exs_333_0;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_exs_339_0;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_exs_345_0;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_exs_351_0;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_16;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_17;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_18;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_19;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_20;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_21;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_22;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_23;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_24;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_25;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_26;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_27;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_28;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_29;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_30;
  wire [4:0] libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_31;
  wire IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_31_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_48_cse;
  reg reg_FpMul_8U_23U_lor_3_lpi_1_dfm_4_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_51_cse;
  wire FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_54_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_57_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_60_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_63_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_66_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_69_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_72_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_75_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_78_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_81_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_84_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_87_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_90_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_93_cse;
  wire mul_loop_mul_if_aelse_and_32_cse;
  wire MulIn_data_and_cse;
  wire IsZero_8U_23U_aelse_and_32_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_48_cse;
  wire IsZero_8U_23U_aelse_and_33_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_51_cse;
  wire IsZero_8U_23U_aelse_and_34_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_54_cse;
  wire IsZero_8U_23U_aelse_and_35_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_57_cse;
  wire IsZero_8U_23U_aelse_and_36_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_60_cse;
  wire IsZero_8U_23U_aelse_and_37_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_63_cse;
  wire IsZero_8U_23U_aelse_and_38_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_66_cse;
  wire IsZero_8U_23U_aelse_and_39_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_69_cse;
  wire IsZero_8U_23U_aelse_and_40_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_72_cse;
  wire IsZero_8U_23U_aelse_and_41_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_75_cse;
  wire IsZero_8U_23U_aelse_and_42_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_78_cse;
  wire IsZero_8U_23U_aelse_and_43_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_81_cse;
  wire IsZero_8U_23U_aelse_and_44_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_84_cse;
  wire IsZero_8U_23U_aelse_and_45_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_87_cse;
  wire IsZero_8U_23U_aelse_and_46_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_90_cse;
  wire IsZero_8U_23U_aelse_and_47_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_93_cse;
  wire mul_loop_mul_if_aelse_and_48_cse;
  wire MulIn_data_and_1_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_96_cse;
  wire MulIn_data_and_2_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_96_cse;
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_31_cse;
  wire IsNaN_8U_23U_aelse_and_48_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_98_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_99_cse;
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_29_cse;
  wire IsNaN_8U_23U_aelse_and_50_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_100_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_102_cse;
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_27_cse;
  wire IsNaN_8U_23U_aelse_and_52_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_102_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_105_cse;
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_25_cse;
  wire IsNaN_8U_23U_aelse_and_54_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_104_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_108_cse;
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_23_cse;
  wire IsNaN_8U_23U_aelse_and_56_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_106_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_111_cse;
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_21_cse;
  wire IsNaN_8U_23U_aelse_and_58_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_108_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_114_cse;
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_19_cse;
  wire IsNaN_8U_23U_aelse_and_60_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_110_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_117_cse;
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_17_cse;
  wire IsNaN_8U_23U_aelse_and_62_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_112_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_120_cse;
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_15_cse;
  wire IsNaN_8U_23U_aelse_and_64_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_114_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_123_cse;
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_13_cse;
  wire IsNaN_8U_23U_aelse_and_66_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_116_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_126_cse;
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_11_cse;
  wire IsNaN_8U_23U_aelse_and_68_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_118_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_129_cse;
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_9_cse;
  wire IsNaN_8U_23U_aelse_and_70_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_120_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_132_cse;
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_7_cse;
  wire IsNaN_8U_23U_aelse_and_72_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_122_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_135_cse;
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_5_cse;
  wire IsNaN_8U_23U_aelse_and_74_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_124_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_138_cse;
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_3_cse;
  wire IsNaN_8U_23U_aelse_and_76_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_126_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_141_cse;
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_1_cse;
  wire IsNaN_8U_23U_aelse_and_78_cse;
  wire mul_loop_mul_if_aelse_and_64_cse;
  wire or_cse;
  wire or_4962_cse;
  wire or_4959_cse;
  wire or_4956_cse;
  wire or_4953_cse;
  wire and_2876_cse;
  wire or_4947_cse;
  wire or_4944_cse;
  wire or_4941_cse;
  wire and_2868_cse;
  wire or_4934_cse;
  wire or_4931_cse;
  wire or_4927_cse;
  wire or_4924_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_128_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_131_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_134_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_137_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_140_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_143_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_146_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_149_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_152_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_155_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_158_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_161_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_164_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_167_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_170_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_173_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_144_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_147_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_150_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_153_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_156_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_159_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_162_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_165_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_168_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_171_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_174_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_177_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_180_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_183_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_186_cse;
  wire FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_189_cse;
  wire FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_16_cse;
  wire FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_17_cse;
  wire FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_18_cse;
  wire FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_19_cse;
  wire FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_20_cse;
  wire FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_21_cse;
  wire FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_22_cse;
  wire FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_23_cse;
  wire FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_24_cse;
  wire FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_25_cse;
  wire FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_26_cse;
  wire FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_27_cse;
  wire FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_28_cse;
  wire FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_29_cse;
  wire FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_30_cse;
  wire FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_31_cse;
  wire MulIn_data_and_3_cse;
  wire IsZero_8U_23U_aelse_and_48_cse;
  wire IsZero_8U_23U_aelse_and_49_cse;
  wire IsZero_8U_23U_aelse_and_50_cse;
  wire IsZero_8U_23U_aelse_and_51_cse;
  wire IsZero_8U_23U_aelse_and_52_cse;
  wire IsZero_8U_23U_aelse_and_53_cse;
  wire IsZero_8U_23U_aelse_and_54_cse;
  wire IsZero_8U_23U_aelse_and_55_cse;
  wire IsZero_8U_23U_aelse_and_56_cse;
  wire IsZero_8U_23U_aelse_and_57_cse;
  wire IsZero_8U_23U_aelse_and_58_cse;
  wire IsZero_8U_23U_aelse_and_59_cse;
  wire IsZero_8U_23U_aelse_and_60_cse;
  wire IsZero_8U_23U_aelse_and_61_cse;
  wire IsZero_8U_23U_aelse_and_62_cse;
  wire IsZero_8U_23U_aelse_and_63_cse;
  wire mul_loop_mul_if_aelse_and_16_cse;
  reg reg_FpMul_8U_23U_lor_4_lpi_1_dfm_4_cse;
  reg reg_FpMul_8U_23U_lor_5_lpi_1_dfm_4_cse;
  reg reg_FpMul_8U_23U_lor_6_lpi_1_dfm_4_cse;
  reg reg_FpMul_8U_23U_lor_7_lpi_1_dfm_4_cse;
  reg reg_FpMul_8U_23U_lor_8_lpi_1_dfm_4_cse;
  reg reg_FpMul_8U_23U_lor_9_lpi_1_dfm_4_cse;
  reg reg_FpMul_8U_23U_lor_10_lpi_1_dfm_4_cse;
  reg reg_FpMul_8U_23U_lor_11_lpi_1_dfm_4_cse;
  reg reg_FpMul_8U_23U_lor_12_lpi_1_dfm_4_cse;
  reg reg_FpMul_8U_23U_lor_13_lpi_1_dfm_4_cse;
  reg reg_FpMul_8U_23U_lor_14_lpi_1_dfm_4_cse;
  reg reg_FpMul_8U_23U_lor_15_lpi_1_dfm_4_cse;
  reg reg_FpMul_8U_23U_lor_16_lpi_1_dfm_4_cse;
  reg reg_FpMul_8U_23U_lor_17_lpi_1_dfm_4_cse;
  reg reg_FpMul_8U_23U_lor_lpi_1_dfm_4_cse;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_cse;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_1_cse;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_2_cse;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_3_cse;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_4_cse;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_5_cse;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_6_cse;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_7_cse;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_8_cse;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_9_cse;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_10_cse;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_11_cse;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_12_cse;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_13_cse;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_14_cse;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_15_cse;
  wire nor_821_cse;
  wire mux_1690_cse;
  wire mux_1695_cse;
  wire mux_1700_cse;
  wire mux_1705_cse;
  wire mux_1710_cse;
  wire mux_1715_cse;
  wire mux_1720_cse;
  wire mux_1725_cse;
  wire mux_1730_cse;
  wire mux_1735_cse;
  wire mux_1741_cse;
  wire mux_1747_cse;
  wire mux_1752_cse;
  wire mux_1758_cse;
  wire mux_1764_cse;
  wire mux_1769_cse;
  wire nor_1477_cse;
  wire nor_1413_cse;
  wire mux_1680_itm;
  wire mux_1681_itm;
  wire mux_1682_itm;
  wire mux_1683_itm;
  wire mux_1684_itm;
  wire mux_1685_itm;
  wire mux_1686_itm;
  wire mux_1687_itm;
  wire mux_1688_itm;
  wire mul_loop_mul_1_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire mul_loop_mul_2_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire mul_loop_mul_3_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire mul_loop_mul_4_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire mul_loop_mul_5_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire mul_loop_mul_6_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire mul_loop_mul_7_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire mul_loop_mul_8_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire mul_loop_mul_9_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire mul_loop_mul_10_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire mul_loop_mul_11_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire mul_loop_mul_12_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire mul_loop_mul_13_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire mul_loop_mul_14_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire mul_loop_mul_15_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire mul_loop_mul_16_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire mul_loop_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire mul_loop_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire mul_loop_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire mul_loop_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire mul_loop_mul_5_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire mul_loop_mul_6_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire mul_loop_mul_7_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire mul_loop_mul_8_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire mul_loop_mul_9_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire mul_loop_mul_10_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire mul_loop_mul_11_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire mul_loop_mul_12_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire mul_loop_mul_13_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire mul_loop_mul_14_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire mul_loop_mul_15_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire mul_loop_mul_16_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire mul_loop_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  wire mul_loop_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  wire mul_loop_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  wire mul_loop_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  wire mul_loop_mul_5_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  wire mul_loop_mul_6_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  wire mul_loop_mul_7_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  wire mul_loop_mul_8_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  wire mul_loop_mul_9_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  wire mul_loop_mul_10_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  wire mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  wire mul_loop_mul_12_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  wire mul_loop_mul_13_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  wire mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  wire mul_loop_mul_15_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  wire mul_loop_mul_16_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  wire[0:0] iExpoWidth_oExpoWidth_prb;
  wire[0:0] iMantWidth_oMantWidth_prb;
  wire[0:0] iMantWidth_oMantWidth_prb_1;
  wire[0:0] iExpoWidth_oExpoWidth_prb_1;
  wire[0:0] iMantWidth_oMantWidth_prb_2;
  wire[0:0] iExpoWidth_oExpoWidth_prb_2;
  wire[0:0] iMantWidth_oMantWidth_prb_3;
  wire[0:0] iMantWidth_oMantWidth_prb_4;
  wire[0:0] iExpoWidth_oExpoWidth_prb_3;
  wire[0:0] iMantWidth_oMantWidth_prb_5;
  wire[0:0] iExpoWidth_oExpoWidth_prb_4;
  wire[0:0] iMantWidth_oMantWidth_prb_6;
  wire[0:0] iMantWidth_oMantWidth_prb_7;
  wire[0:0] iExpoWidth_oExpoWidth_prb_5;
  wire[0:0] iMantWidth_oMantWidth_prb_8;
  wire[0:0] iExpoWidth_oExpoWidth_prb_6;
  wire[0:0] iMantWidth_oMantWidth_prb_9;
  wire[0:0] iMantWidth_oMantWidth_prb_10;
  wire[0:0] iExpoWidth_oExpoWidth_prb_7;
  wire[0:0] iMantWidth_oMantWidth_prb_11;
  wire[0:0] iExpoWidth_oExpoWidth_prb_8;
  wire[0:0] iMantWidth_oMantWidth_prb_12;
  wire[0:0] iMantWidth_oMantWidth_prb_13;
  wire[0:0] iExpoWidth_oExpoWidth_prb_9;
  wire[0:0] iMantWidth_oMantWidth_prb_14;
  wire[0:0] iExpoWidth_oExpoWidth_prb_10;
  wire[0:0] iMantWidth_oMantWidth_prb_15;
  wire[0:0] iMantWidth_oMantWidth_prb_16;
  wire[0:0] iExpoWidth_oExpoWidth_prb_11;
  wire[0:0] iMantWidth_oMantWidth_prb_17;
  wire[0:0] iExpoWidth_oExpoWidth_prb_12;
  wire[0:0] iMantWidth_oMantWidth_prb_18;
  wire[0:0] iMantWidth_oMantWidth_prb_19;
  wire[0:0] iExpoWidth_oExpoWidth_prb_13;
  wire[0:0] iMantWidth_oMantWidth_prb_20;
  wire[0:0] iExpoWidth_oExpoWidth_prb_14;
  wire[0:0] iMantWidth_oMantWidth_prb_21;
  wire[0:0] iMantWidth_oMantWidth_prb_22;
  wire[0:0] iExpoWidth_oExpoWidth_prb_15;
  wire[0:0] iMantWidth_oMantWidth_prb_23;
  wire[0:0] iExpoWidth_oExpoWidth_prb_16;
  wire[0:0] iMantWidth_oMantWidth_prb_24;
  wire[0:0] iMantWidth_oMantWidth_prb_25;
  wire[0:0] iExpoWidth_oExpoWidth_prb_17;
  wire[0:0] iMantWidth_oMantWidth_prb_26;
  wire[0:0] iExpoWidth_oExpoWidth_prb_18;
  wire[0:0] iMantWidth_oMantWidth_prb_27;
  wire[0:0] iMantWidth_oMantWidth_prb_28;
  wire[0:0] iExpoWidth_oExpoWidth_prb_19;
  wire[0:0] iMantWidth_oMantWidth_prb_29;
  wire[0:0] iExpoWidth_oExpoWidth_prb_20;
  wire[0:0] iMantWidth_oMantWidth_prb_30;
  wire[0:0] iMantWidth_oMantWidth_prb_31;
  wire[0:0] iExpoWidth_oExpoWidth_prb_21;
  wire[0:0] iMantWidth_oMantWidth_prb_32;
  wire[0:0] iExpoWidth_oExpoWidth_prb_22;
  wire[0:0] iMantWidth_oMantWidth_prb_33;
  wire[0:0] iMantWidth_oMantWidth_prb_34;
  wire[0:0] iExpoWidth_oExpoWidth_prb_23;
  wire[0:0] iMantWidth_oMantWidth_prb_35;
  wire[0:0] iExpoWidth_oExpoWidth_prb_24;
  wire[0:0] iMantWidth_oMantWidth_prb_36;
  wire[0:0] iMantWidth_oMantWidth_prb_37;
  wire[0:0] iExpoWidth_oExpoWidth_prb_25;
  wire[0:0] iMantWidth_oMantWidth_prb_38;
  wire[0:0] iExpoWidth_oExpoWidth_prb_26;
  wire[0:0] iMantWidth_oMantWidth_prb_39;
  wire[0:0] iMantWidth_oMantWidth_prb_40;
  wire[0:0] iExpoWidth_oExpoWidth_prb_27;
  wire[0:0] iMantWidth_oMantWidth_prb_41;
  wire[0:0] iExpoWidth_oExpoWidth_prb_28;
  wire[0:0] iMantWidth_oMantWidth_prb_42;
  wire[0:0] iMantWidth_oMantWidth_prb_43;
  wire[0:0] iExpoWidth_oExpoWidth_prb_29;
  wire[0:0] iMantWidth_oMantWidth_prb_44;
  wire[0:0] iExpoWidth_oExpoWidth_prb_30;
  wire[0:0] iMantWidth_oMantWidth_prb_45;
  wire[0:0] iMantWidth_oMantWidth_prb_46;
  wire[0:0] iExpoWidth_oExpoWidth_prb_31;
  wire[0:0] iMantWidth_oMantWidth_prb_47;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_33_nl;
  wire[9:0] FpMul_8U_23U_nor_32_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_33_nl;
  wire[2:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_32_nl;
  wire[2:0] FpMul_8U_23U_nor_31_nl;
  wire[2:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_32_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_16_nl;
  wire[9:0] FpMul_8U_23U_nor_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_34_nl;
  wire[3:0] FpMul_8U_23U_FpMul_8U_23U_and_95_nl;
  wire[3:0] SetToInf_8U_23U_mux_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_64_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_97_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_96_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_96_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_112_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_35_nl;
  wire[9:0] FpMul_8U_23U_nor_34_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_35_nl;
  wire[2:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_34_nl;
  wire[2:0] FpMul_8U_23U_nor_33_nl;
  wire[2:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_36_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_17_nl;
  wire[9:0] FpMul_8U_23U_nor_16_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_37_nl;
  wire[3:0] FpMul_8U_23U_FpMul_8U_23U_and_98_nl;
  wire[3:0] SetToInf_8U_23U_mux_2_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_66_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_100_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_97_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_99_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_113_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_37_nl;
  wire[9:0] FpMul_8U_23U_nor_36_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_38_nl;
  wire[2:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_36_nl;
  wire[2:0] FpMul_8U_23U_nor_35_nl;
  wire[2:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_39_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_18_nl;
  wire[9:0] FpMul_8U_23U_nor_17_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_40_nl;
  wire[3:0] FpMul_8U_23U_FpMul_8U_23U_and_101_nl;
  wire[3:0] SetToInf_8U_23U_mux_4_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_68_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_103_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_98_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_102_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_114_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_39_nl;
  wire[9:0] FpMul_8U_23U_nor_38_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_41_nl;
  wire[2:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_38_nl;
  wire[2:0] FpMul_8U_23U_nor_37_nl;
  wire[2:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_42_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_19_nl;
  wire[9:0] FpMul_8U_23U_nor_18_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_43_nl;
  wire[3:0] FpMul_8U_23U_FpMul_8U_23U_and_104_nl;
  wire[3:0] SetToInf_8U_23U_mux_6_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_70_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_106_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_99_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_105_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_115_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_41_nl;
  wire[9:0] FpMul_8U_23U_nor_40_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_44_nl;
  wire[2:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_40_nl;
  wire[2:0] FpMul_8U_23U_nor_39_nl;
  wire[2:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_45_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_20_nl;
  wire[9:0] FpMul_8U_23U_nor_19_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_46_nl;
  wire[3:0] FpMul_8U_23U_FpMul_8U_23U_and_107_nl;
  wire[3:0] SetToInf_8U_23U_mux_8_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_72_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_109_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_100_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_108_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_116_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_43_nl;
  wire[9:0] FpMul_8U_23U_nor_42_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_47_nl;
  wire[2:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_42_nl;
  wire[2:0] FpMul_8U_23U_nor_41_nl;
  wire[2:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_48_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_21_nl;
  wire[9:0] FpMul_8U_23U_nor_20_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_49_nl;
  wire[3:0] FpMul_8U_23U_FpMul_8U_23U_and_110_nl;
  wire[3:0] SetToInf_8U_23U_mux_10_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_74_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_112_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_101_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_111_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_117_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_45_nl;
  wire[9:0] FpMul_8U_23U_nor_44_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_50_nl;
  wire[2:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_44_nl;
  wire[2:0] FpMul_8U_23U_nor_43_nl;
  wire[2:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_51_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_22_nl;
  wire[9:0] FpMul_8U_23U_nor_21_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_52_nl;
  wire[3:0] FpMul_8U_23U_FpMul_8U_23U_and_113_nl;
  wire[3:0] SetToInf_8U_23U_mux_12_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_76_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_115_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_102_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_114_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_118_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_47_nl;
  wire[9:0] FpMul_8U_23U_nor_46_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_53_nl;
  wire[2:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_46_nl;
  wire[2:0] FpMul_8U_23U_nor_45_nl;
  wire[2:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_54_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_23_nl;
  wire[9:0] FpMul_8U_23U_nor_22_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_55_nl;
  wire[3:0] FpMul_8U_23U_FpMul_8U_23U_and_116_nl;
  wire[3:0] SetToInf_8U_23U_mux_14_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_78_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_118_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_103_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_117_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_119_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_49_nl;
  wire[9:0] FpMul_8U_23U_nor_48_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_56_nl;
  wire[2:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_48_nl;
  wire[2:0] FpMul_8U_23U_nor_47_nl;
  wire[2:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_57_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_24_nl;
  wire[9:0] FpMul_8U_23U_nor_23_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_16_nl;
  wire[3:0] FpMul_8U_23U_FpMul_8U_23U_and_119_nl;
  wire[3:0] SetToInf_8U_23U_mux_16_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_80_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_121_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_104_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_120_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_120_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_51_nl;
  wire[9:0] FpMul_8U_23U_nor_50_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_58_nl;
  wire[2:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_50_nl;
  wire[2:0] FpMul_8U_23U_nor_49_nl;
  wire[2:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_59_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_25_nl;
  wire[9:0] FpMul_8U_23U_nor_24_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_18_nl;
  wire[3:0] FpMul_8U_23U_FpMul_8U_23U_and_122_nl;
  wire[3:0] SetToInf_8U_23U_mux_18_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_82_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_124_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_105_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_123_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_121_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_53_nl;
  wire[9:0] FpMul_8U_23U_nor_52_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_60_nl;
  wire[2:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_52_nl;
  wire[2:0] FpMul_8U_23U_nor_51_nl;
  wire[2:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_61_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_26_nl;
  wire[9:0] FpMul_8U_23U_nor_25_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_20_nl;
  wire[3:0] FpMul_8U_23U_FpMul_8U_23U_and_125_nl;
  wire[3:0] SetToInf_8U_23U_mux_20_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_84_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_127_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_106_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_126_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_122_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_55_nl;
  wire[9:0] FpMul_8U_23U_nor_54_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_62_nl;
  wire[2:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_54_nl;
  wire[2:0] FpMul_8U_23U_nor_53_nl;
  wire[2:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_63_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_27_nl;
  wire[9:0] FpMul_8U_23U_nor_26_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_22_nl;
  wire[3:0] FpMul_8U_23U_FpMul_8U_23U_and_128_nl;
  wire[3:0] SetToInf_8U_23U_mux_22_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_86_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_130_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_107_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_129_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_123_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_57_nl;
  wire[9:0] FpMul_8U_23U_nor_56_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_64_nl;
  wire[2:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_56_nl;
  wire[2:0] FpMul_8U_23U_nor_55_nl;
  wire[2:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_65_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_28_nl;
  wire[9:0] FpMul_8U_23U_nor_27_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_24_nl;
  wire[3:0] FpMul_8U_23U_FpMul_8U_23U_and_131_nl;
  wire[3:0] SetToInf_8U_23U_mux_24_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_88_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_133_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_108_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_132_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_124_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_59_nl;
  wire[9:0] FpMul_8U_23U_nor_58_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_66_nl;
  wire[2:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_58_nl;
  wire[2:0] FpMul_8U_23U_nor_57_nl;
  wire[2:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_67_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_29_nl;
  wire[9:0] FpMul_8U_23U_nor_28_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_26_nl;
  wire[3:0] FpMul_8U_23U_FpMul_8U_23U_and_134_nl;
  wire[3:0] SetToInf_8U_23U_mux_26_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_90_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_136_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_109_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_135_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_125_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_61_nl;
  wire[9:0] FpMul_8U_23U_nor_60_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_68_nl;
  wire[2:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_60_nl;
  wire[2:0] FpMul_8U_23U_nor_59_nl;
  wire[2:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_69_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_30_nl;
  wire[9:0] FpMul_8U_23U_nor_29_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_28_nl;
  wire[3:0] FpMul_8U_23U_FpMul_8U_23U_and_137_nl;
  wire[3:0] SetToInf_8U_23U_mux_28_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_92_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_139_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_110_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_138_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_126_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_63_nl;
  wire[9:0] FpMul_8U_23U_nor_62_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_70_nl;
  wire[2:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_62_nl;
  wire[2:0] FpMul_8U_23U_nor_61_nl;
  wire[2:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_71_nl;
  wire[9:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_31_nl;
  wire[9:0] FpMul_8U_23U_nor_30_nl;
  wire[9:0] FpMantWidthDec_8U_47U_23U_0U_0U_mux_30_nl;
  wire[3:0] FpMul_8U_23U_FpMul_8U_23U_and_140_nl;
  wire[3:0] SetToInf_8U_23U_mux_30_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_94_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_142_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_111_nl;
  wire[1:0] FpMul_8U_23U_FpMul_8U_23U_and_141_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_127_nl;
  wire[0:0] mux_19_nl;
  wire[0:0] mux_18_nl;
  wire[0:0] mux_16_nl;
  wire[0:0] mux_17_nl;
  wire[0:0] mux_29_nl;
  wire[0:0] mux_28_nl;
  wire[0:0] mux_26_nl;
  wire[0:0] mux_27_nl;
  wire[0:0] mux_39_nl;
  wire[0:0] mux_38_nl;
  wire[0:0] mux_36_nl;
  wire[0:0] mux_37_nl;
  wire[0:0] mux_49_nl;
  wire[0:0] mux_48_nl;
  wire[0:0] mux_46_nl;
  wire[0:0] mux_47_nl;
  wire[0:0] mux_59_nl;
  wire[0:0] mux_58_nl;
  wire[0:0] mux_56_nl;
  wire[0:0] mux_57_nl;
  wire[0:0] mux_66_nl;
  wire[0:0] mux_65_nl;
  wire[0:0] mux_63_nl;
  wire[0:0] mux_64_nl;
  wire[0:0] mux_73_nl;
  wire[0:0] mux_72_nl;
  wire[0:0] mux_70_nl;
  wire[0:0] mux_71_nl;
  wire[0:0] mux_83_nl;
  wire[0:0] mux_82_nl;
  wire[0:0] mux_80_nl;
  wire[0:0] mux_81_nl;
  wire[0:0] mux_93_nl;
  wire[0:0] mux_92_nl;
  wire[0:0] mux_90_nl;
  wire[0:0] mux_91_nl;
  wire[0:0] mux_100_nl;
  wire[0:0] mux_99_nl;
  wire[0:0] mux_97_nl;
  wire[0:0] mux_98_nl;
  wire[0:0] mux_107_nl;
  wire[0:0] mux_106_nl;
  wire[0:0] mux_104_nl;
  wire[0:0] mux_105_nl;
  wire[0:0] mux_114_nl;
  wire[0:0] mux_113_nl;
  wire[0:0] mux_111_nl;
  wire[0:0] mux_112_nl;
  wire[0:0] mux_124_nl;
  wire[0:0] mux_123_nl;
  wire[0:0] mux_121_nl;
  wire[0:0] mux_122_nl;
  wire[0:0] mux_131_nl;
  wire[0:0] mux_130_nl;
  wire[0:0] mux_128_nl;
  wire[0:0] mux_129_nl;
  wire[0:0] mux_141_nl;
  wire[0:0] mux_140_nl;
  wire[0:0] mux_138_nl;
  wire[0:0] mux_139_nl;
  wire[0:0] mux_151_nl;
  wire[0:0] mux_150_nl;
  wire[0:0] mux_148_nl;
  wire[0:0] mux_149_nl;
  wire[0:0] mux_154_nl;
  wire[0:0] mux_153_nl;
  wire[0:0] mux_152_nl;
  wire[0:0] nand_26_nl;
  wire[0:0] mux_172_nl;
  wire[0:0] mux_175_nl;
  wire[0:0] mux_174_nl;
  wire[0:0] and_2249_nl;
  wire[0:0] mux_173_nl;
  wire[0:0] nor_1492_nl;
  wire[0:0] nor_1493_nl;
  wire[0:0] mux_176_nl;
  wire[0:0] mux_183_nl;
  wire[0:0] mux_182_nl;
  wire[0:0] mux_180_nl;
  wire[0:0] mux_179_nl;
  wire[0:0] mux_178_nl;
  wire[0:0] mux_181_nl;
  wire[0:0] or_308_nl;
  wire[0:0] mux_186_nl;
  wire[0:0] nor_1489_nl;
  wire[0:0] mux_185_nl;
  wire[0:0] mux_190_nl;
  wire[0:0] mux_189_nl;
  wire[0:0] and_2248_nl;
  wire[0:0] mux_188_nl;
  wire[0:0] nor_1481_nl;
  wire[0:0] nor_1482_nl;
  wire[0:0] nor_1483_nl;
  wire[0:0] mux_197_nl;
  wire[0:0] mux_196_nl;
  wire[0:0] mux_194_nl;
  wire[0:0] mux_193_nl;
  wire[0:0] mux_192_nl;
  wire[0:0] mux_195_nl;
  wire[0:0] or_331_nl;
  wire[0:0] mux_201_nl;
  wire[0:0] mux_198_nl;
  wire[0:0] or_335_nl;
  wire[0:0] mux_200_nl;
  wire[0:0] or_342_nl;
  wire[0:0] mux_205_nl;
  wire[0:0] mux_204_nl;
  wire[0:0] and_2247_nl;
  wire[0:0] mux_203_nl;
  wire[0:0] nor_1478_nl;
  wire[0:0] nor_1479_nl;
  wire[0:0] mux_212_nl;
  wire[0:0] mux_211_nl;
  wire[0:0] mux_209_nl;
  wire[0:0] mux_208_nl;
  wire[0:0] mux_207_nl;
  wire[0:0] mux_210_nl;
  wire[0:0] or_359_nl;
  wire[0:0] mux_215_nl;
  wire[0:0] nor_1475_nl;
  wire[0:0] mux_214_nl;
  wire[0:0] nor_1476_nl;
  wire[0:0] mux_219_nl;
  wire[0:0] mux_218_nl;
  wire[0:0] and_2246_nl;
  wire[0:0] mux_217_nl;
  wire[0:0] nor_1471_nl;
  wire[0:0] nor_1472_nl;
  wire[0:0] nor_1473_nl;
  wire[0:0] mux_226_nl;
  wire[0:0] mux_225_nl;
  wire[0:0] mux_223_nl;
  wire[0:0] mux_222_nl;
  wire[0:0] mux_221_nl;
  wire[0:0] mux_224_nl;
  wire[0:0] or_382_nl;
  wire[0:0] mux_229_nl;
  wire[0:0] nor_1469_nl;
  wire[0:0] mux_228_nl;
  wire[0:0] nor_1470_nl;
  wire[0:0] mux_233_nl;
  wire[0:0] mux_232_nl;
  wire[0:0] and_2245_nl;
  wire[0:0] mux_231_nl;
  wire[0:0] nor_1465_nl;
  wire[0:0] nor_1466_nl;
  wire[0:0] nor_1467_nl;
  wire[0:0] mux_240_nl;
  wire[0:0] mux_239_nl;
  wire[0:0] mux_237_nl;
  wire[0:0] mux_236_nl;
  wire[0:0] mux_235_nl;
  wire[0:0] mux_238_nl;
  wire[0:0] or_405_nl;
  wire[0:0] mux_244_nl;
  wire[0:0] mux_241_nl;
  wire[0:0] or_409_nl;
  wire[0:0] mux_243_nl;
  wire[0:0] or_417_nl;
  wire[0:0] mux_248_nl;
  wire[0:0] mux_247_nl;
  wire[0:0] and_2244_nl;
  wire[0:0] mux_246_nl;
  wire[0:0] nor_1461_nl;
  wire[0:0] nor_1462_nl;
  wire[0:0] nor_1463_nl;
  wire[0:0] mux_255_nl;
  wire[0:0] mux_254_nl;
  wire[0:0] mux_252_nl;
  wire[0:0] mux_251_nl;
  wire[0:0] mux_250_nl;
  wire[0:0] mux_253_nl;
  wire[0:0] or_434_nl;
  wire[0:0] mux_258_nl;
  wire[0:0] nor_1459_nl;
  wire[0:0] mux_257_nl;
  wire[0:0] nor_1460_nl;
  wire[0:0] mux_262_nl;
  wire[0:0] mux_261_nl;
  wire[0:0] and_2243_nl;
  wire[0:0] mux_260_nl;
  wire[0:0] nor_1455_nl;
  wire[0:0] nor_1456_nl;
  wire[0:0] nor_1457_nl;
  wire[0:0] mux_269_nl;
  wire[0:0] mux_268_nl;
  wire[0:0] mux_266_nl;
  wire[0:0] mux_265_nl;
  wire[0:0] mux_264_nl;
  wire[0:0] mux_267_nl;
  wire[0:0] or_457_nl;
  wire[0:0] mux_272_nl;
  wire[0:0] nor_1453_nl;
  wire[0:0] mux_271_nl;
  wire[0:0] nor_1454_nl;
  wire[0:0] mux_276_nl;
  wire[0:0] mux_275_nl;
  wire[0:0] and_2242_nl;
  wire[0:0] mux_274_nl;
  wire[0:0] nor_1449_nl;
  wire[0:0] nor_1450_nl;
  wire[0:0] nor_1451_nl;
  wire[0:0] mux_283_nl;
  wire[0:0] mux_282_nl;
  wire[0:0] mux_280_nl;
  wire[0:0] mux_279_nl;
  wire[0:0] mux_278_nl;
  wire[0:0] mux_281_nl;
  wire[0:0] or_480_nl;
  wire[0:0] mux_287_nl;
  wire[0:0] mux_284_nl;
  wire[0:0] or_484_nl;
  wire[0:0] mux_286_nl;
  wire[0:0] or_491_nl;
  wire[0:0] mux_291_nl;
  wire[0:0] mux_290_nl;
  wire[0:0] and_2241_nl;
  wire[0:0] mux_289_nl;
  wire[0:0] nor_1445_nl;
  wire[0:0] nor_1446_nl;
  wire[0:0] nor_1447_nl;
  wire[0:0] mux_298_nl;
  wire[0:0] mux_297_nl;
  wire[0:0] mux_295_nl;
  wire[0:0] mux_294_nl;
  wire[0:0] mux_293_nl;
  wire[0:0] mux_296_nl;
  wire[0:0] or_508_nl;
  wire[0:0] mux_302_nl;
  wire[0:0] mux_299_nl;
  wire[0:0] or_512_nl;
  wire[0:0] mux_301_nl;
  wire[0:0] or_520_nl;
  wire[0:0] mux_306_nl;
  wire[0:0] mux_305_nl;
  wire[0:0] and_2240_nl;
  wire[0:0] mux_304_nl;
  wire[0:0] nor_1441_nl;
  wire[0:0] nor_1442_nl;
  wire[0:0] nor_1443_nl;
  wire[0:0] mux_313_nl;
  wire[0:0] mux_312_nl;
  wire[0:0] mux_310_nl;
  wire[0:0] mux_309_nl;
  wire[0:0] mux_308_nl;
  wire[0:0] mux_311_nl;
  wire[0:0] or_537_nl;
  wire[0:0] mux_317_nl;
  wire[0:0] mux_314_nl;
  wire[0:0] or_541_nl;
  wire[0:0] mux_316_nl;
  wire[0:0] mux_321_nl;
  wire[0:0] mux_320_nl;
  wire[0:0] and_2239_nl;
  wire[0:0] mux_319_nl;
  wire[0:0] nor_1437_nl;
  wire[0:0] nor_1438_nl;
  wire[0:0] nor_1439_nl;
  wire[0:0] mux_328_nl;
  wire[0:0] mux_327_nl;
  wire[0:0] mux_325_nl;
  wire[0:0] mux_324_nl;
  wire[0:0] mux_323_nl;
  wire[0:0] mux_326_nl;
  wire[0:0] or_566_nl;
  wire[0:0] mux_331_nl;
  wire[0:0] nor_1435_nl;
  wire[0:0] mux_330_nl;
  wire[0:0] nor_1436_nl;
  wire[0:0] mux_335_nl;
  wire[0:0] mux_334_nl;
  wire[0:0] and_2238_nl;
  wire[0:0] mux_333_nl;
  wire[0:0] nor_1431_nl;
  wire[0:0] nor_1432_nl;
  wire[0:0] nor_1433_nl;
  wire[0:0] mux_342_nl;
  wire[0:0] mux_341_nl;
  wire[0:0] mux_339_nl;
  wire[0:0] mux_338_nl;
  wire[0:0] mux_337_nl;
  wire[0:0] mux_340_nl;
  wire[0:0] or_589_nl;
  wire[0:0] mux_345_nl;
  wire[0:0] nor_1429_nl;
  wire[0:0] mux_344_nl;
  wire[0:0] nor_1430_nl;
  wire[0:0] mux_349_nl;
  wire[0:0] mux_348_nl;
  wire[0:0] and_2237_nl;
  wire[0:0] mux_347_nl;
  wire[0:0] nor_1425_nl;
  wire[0:0] nor_1426_nl;
  wire[0:0] nor_1427_nl;
  wire[0:0] mux_356_nl;
  wire[0:0] mux_355_nl;
  wire[0:0] mux_353_nl;
  wire[0:0] mux_352_nl;
  wire[0:0] mux_351_nl;
  wire[0:0] mux_354_nl;
  wire[0:0] or_612_nl;
  wire[0:0] mux_359_nl;
  wire[0:0] nor_1423_nl;
  wire[0:0] mux_358_nl;
  wire[0:0] nor_1424_nl;
  wire[0:0] mux_363_nl;
  wire[0:0] mux_362_nl;
  wire[0:0] and_2236_nl;
  wire[0:0] mux_361_nl;
  wire[0:0] nor_1419_nl;
  wire[0:0] nor_1420_nl;
  wire[0:0] nor_1421_nl;
  wire[0:0] mux_370_nl;
  wire[0:0] mux_369_nl;
  wire[0:0] mux_367_nl;
  wire[0:0] mux_366_nl;
  wire[0:0] mux_365_nl;
  wire[0:0] mux_368_nl;
  wire[0:0] or_635_nl;
  wire[0:0] mux_373_nl;
  wire[0:0] nor_1417_nl;
  wire[0:0] mux_372_nl;
  wire[0:0] nor_1418_nl;
  wire[0:0] mux_377_nl;
  wire[0:0] mux_376_nl;
  wire[0:0] and_2235_nl;
  wire[0:0] mux_375_nl;
  wire[0:0] nor_1414_nl;
  wire[0:0] nor_1415_nl;
  wire[0:0] mux_384_nl;
  wire[0:0] mux_383_nl;
  wire[0:0] mux_381_nl;
  wire[0:0] mux_380_nl;
  wire[0:0] mux_379_nl;
  wire[0:0] mux_382_nl;
  wire[0:0] or_658_nl;
  wire[0:0] mux_387_nl;
  wire[0:0] nor_1411_nl;
  wire[0:0] mux_386_nl;
  wire[0:0] nor_1412_nl;
  wire[0:0] mux_391_nl;
  wire[0:0] mux_390_nl;
  wire[0:0] and_2234_nl;
  wire[0:0] mux_389_nl;
  wire[0:0] nor_1407_nl;
  wire[0:0] nor_1408_nl;
  wire[0:0] nor_1409_nl;
  wire[0:0] mux_398_nl;
  wire[0:0] mux_397_nl;
  wire[0:0] mux_395_nl;
  wire[0:0] mux_394_nl;
  wire[0:0] mux_393_nl;
  wire[0:0] mux_396_nl;
  wire[0:0] or_681_nl;
  wire[0:0] mux_402_nl;
  wire[0:0] mux_399_nl;
  wire[0:0] or_685_nl;
  wire[0:0] mux_401_nl;
  wire[0:0] or_692_nl;
  wire[0:0] mux_404_nl;
  wire[0:0] mux_405_nl;
  wire[0:0] mux_408_nl;
  wire[0:0] or_707_nl;
  wire[0:0] mux_412_nl;
  wire[0:0] or_713_nl;
  wire[0:0] mux_411_nl;
  wire[0:0] mux_415_nl;
  wire[0:0] or_726_nl;
  wire[0:0] mux_418_nl;
  wire[0:0] or_732_nl;
  wire[0:0] mux_417_nl;
  wire[0:0] mux_421_nl;
  wire[0:0] or_742_nl;
  wire[0:0] mux_424_nl;
  wire[0:0] or_751_nl;
  wire[0:0] mux_427_nl;
  wire[0:0] or_760_nl;
  wire[0:0] mux_430_nl;
  wire[0:0] or_769_nl;
  wire[0:0] mux_433_nl;
  wire[0:0] or_778_nl;
  wire[0:0] mux_436_nl;
  wire[0:0] or_787_nl;
  wire[0:0] mux_439_nl;
  wire[0:0] or_796_nl;
  wire[0:0] mux_442_nl;
  wire[0:0] or_805_nl;
  wire[0:0] mux_445_nl;
  wire[0:0] or_814_nl;
  wire[0:0] mux_448_nl;
  wire[0:0] or_823_nl;
  wire[0:0] mux_451_nl;
  wire[0:0] or_832_nl;
  wire[0:0] mux_454_nl;
  wire[0:0] or_841_nl;
  wire[0:0] mux_457_nl;
  wire[0:0] or_850_nl;
  wire[0:0] mux_460_nl;
  wire[0:0] or_859_nl;
  wire[0:0] mux_463_nl;
  wire[0:0] or_868_nl;
  wire[0:0] mux_466_nl;
  wire[0:0] or_877_nl;
  wire[0:0] mux_469_nl;
  wire[0:0] or_886_nl;
  wire[0:0] mux_472_nl;
  wire[0:0] or_892_nl;
  wire[0:0] mux_471_nl;
  wire[0:0] mux_475_nl;
  wire[0:0] or_902_nl;
  wire[0:0] mux_478_nl;
  wire[0:0] or_908_nl;
  wire[0:0] mux_477_nl;
  wire[0:0] mux_481_nl;
  wire[0:0] or_918_nl;
  wire[0:0] mux_484_nl;
  wire[0:0] or_924_nl;
  wire[0:0] mux_483_nl;
  wire[0:0] mux_487_nl;
  wire[0:0] or_934_nl;
  wire[0:0] mux_490_nl;
  wire[0:0] or_940_nl;
  wire[0:0] mux_489_nl;
  wire[0:0] mux_493_nl;
  wire[0:0] or_950_nl;
  wire[0:0] mux_496_nl;
  wire[0:0] or_956_nl;
  wire[0:0] mux_495_nl;
  wire[0:0] mux_499_nl;
  wire[0:0] or_966_nl;
  wire[0:0] mux_502_nl;
  wire[0:0] or_975_nl;
  wire[0:0] and_718_nl;
  wire[0:0] and_719_nl;
  wire[0:0] mux_1616_nl;
  wire[0:0] or_4735_nl;
  wire[0:0] mux_1689_nl;
  wire[0:0] and_2512_nl;
  wire[0:0] mux_1693_nl;
  wire[0:0] nor_1676_nl;
  wire[0:0] or_4963_nl;
  wire[0:0] mux_512_nl;
  wire[0:0] and_2230_nl;
  wire[0:0] mux_511_nl;
  wire[0:0] mux_510_nl;
  wire[0:0] nor_1393_nl;
  wire[0:0] nor_1395_nl;
  wire[0:0] nor_1396_nl;
  wire[0:0] nor_1397_nl;
  wire[0:0] mux_514_nl;
  wire[0:0] nor_1390_nl;
  wire[0:0] mux_515_nl;
  wire[0:0] or_1023_nl;
  wire[0:0] mux_516_nl;
  wire[0:0] nor_1387_nl;
  wire[0:0] nor_1388_nl;
  wire[0:0] mux_520_nl;
  wire[0:0] mux_519_nl;
  wire[0:0] nor_1381_nl;
  wire[0:0] mux_518_nl;
  wire[0:0] and_2229_nl;
  wire[0:0] mux_517_nl;
  wire[0:0] nor_1382_nl;
  wire[0:0] nor_1384_nl;
  wire[0:0] nor_1385_nl;
  wire[0:0] nor_1386_nl;
  wire[0:0] mux_521_nl;
  wire[0:0] nor_1379_nl;
  wire[0:0] nor_1380_nl;
  wire[0:0] mux_526_nl;
  wire[0:0] mux_525_nl;
  wire[0:0] and_2228_nl;
  wire[0:0] mux_524_nl;
  wire[0:0] nor_1373_nl;
  wire[0:0] nor_1375_nl;
  wire[0:0] nor_1376_nl;
  wire[0:0] nor_1377_nl;
  wire[0:0] and_723_nl;
  wire[0:0] and_724_nl;
  wire[0:0] mux_1617_nl;
  wire[0:0] or_4747_nl;
  wire[0:0] mux_1694_nl;
  wire[0:0] and_2534_nl;
  wire[0:0] mux_1698_nl;
  wire[0:0] nor_1671_nl;
  wire[0:0] or_4960_nl;
  wire[0:0] mux_536_nl;
  wire[0:0] and_2224_nl;
  wire[0:0] mux_535_nl;
  wire[0:0] mux_534_nl;
  wire[0:0] nor_1359_nl;
  wire[0:0] nor_1361_nl;
  wire[0:0] nor_1362_nl;
  wire[0:0] nor_1363_nl;
  wire[0:0] mux_538_nl;
  wire[0:0] or_1098_nl;
  wire[0:0] mux_539_nl;
  wire[0:0] or_1103_nl;
  wire[0:0] mux_540_nl;
  wire[0:0] nor_1355_nl;
  wire[0:0] nor_1356_nl;
  wire[0:0] mux_544_nl;
  wire[0:0] mux_543_nl;
  wire[0:0] nor_1349_nl;
  wire[0:0] mux_542_nl;
  wire[0:0] and_2223_nl;
  wire[0:0] mux_541_nl;
  wire[0:0] nor_1350_nl;
  wire[0:0] nor_1352_nl;
  wire[0:0] nor_1353_nl;
  wire[0:0] nor_1354_nl;
  wire[0:0] mux_545_nl;
  wire[0:0] nor_1347_nl;
  wire[0:0] nor_1348_nl;
  wire[0:0] mux_550_nl;
  wire[0:0] mux_549_nl;
  wire[0:0] and_2222_nl;
  wire[0:0] mux_548_nl;
  wire[0:0] nor_1341_nl;
  wire[0:0] nor_1343_nl;
  wire[0:0] nor_1344_nl;
  wire[0:0] nor_1345_nl;
  wire[0:0] and_728_nl;
  wire[0:0] and_729_nl;
  wire[0:0] mux_1618_nl;
  wire[0:0] or_4759_nl;
  wire[0:0] mux_1699_nl;
  wire[0:0] and_2556_nl;
  wire[0:0] mux_1703_nl;
  wire[0:0] nor_1666_nl;
  wire[0:0] or_4957_nl;
  wire[0:0] mux_560_nl;
  wire[0:0] and_2218_nl;
  wire[0:0] mux_559_nl;
  wire[0:0] mux_558_nl;
  wire[0:0] nor_1327_nl;
  wire[0:0] nor_1329_nl;
  wire[0:0] nor_1330_nl;
  wire[0:0] nor_1331_nl;
  wire[0:0] mux_562_nl;
  wire[0:0] nor_1323_nl;
  wire[0:0] nor_1324_nl;
  wire[0:0] mux_563_nl;
  wire[0:0] or_1185_nl;
  wire[0:0] mux_564_nl;
  wire[0:0] nor_1321_nl;
  wire[0:0] nor_1322_nl;
  wire[0:0] mux_568_nl;
  wire[0:0] mux_567_nl;
  wire[0:0] nor_1315_nl;
  wire[0:0] mux_566_nl;
  wire[0:0] and_2217_nl;
  wire[0:0] mux_565_nl;
  wire[0:0] nor_1316_nl;
  wire[0:0] nor_1318_nl;
  wire[0:0] nor_1319_nl;
  wire[0:0] nor_1320_nl;
  wire[0:0] mux_569_nl;
  wire[0:0] nor_1313_nl;
  wire[0:0] nor_1314_nl;
  wire[0:0] mux_574_nl;
  wire[0:0] mux_573_nl;
  wire[0:0] and_2216_nl;
  wire[0:0] mux_572_nl;
  wire[0:0] nor_1307_nl;
  wire[0:0] nor_1309_nl;
  wire[0:0] nor_1310_nl;
  wire[0:0] nor_1311_nl;
  wire[0:0] and_733_nl;
  wire[0:0] and_734_nl;
  wire[0:0] mux_1619_nl;
  wire[0:0] or_4771_nl;
  wire[0:0] mux_1704_nl;
  wire[0:0] and_2578_nl;
  wire[0:0] mux_1708_nl;
  wire[0:0] nor_1661_nl;
  wire[0:0] or_4954_nl;
  wire[0:0] mux_584_nl;
  wire[0:0] and_2212_nl;
  wire[0:0] mux_583_nl;
  wire[0:0] mux_582_nl;
  wire[0:0] nor_1293_nl;
  wire[0:0] nor_1295_nl;
  wire[0:0] nor_1296_nl;
  wire[0:0] nor_1297_nl;
  wire[0:0] mux_588_nl;
  wire[0:0] or_1260_nl;
  wire[0:0] mux_587_nl;
  wire[0:0] or_1263_nl;
  wire[0:0] mux_589_nl;
  wire[0:0] or_1268_nl;
  wire[0:0] mux_590_nl;
  wire[0:0] nor_1291_nl;
  wire[0:0] nor_1292_nl;
  wire[0:0] mux_594_nl;
  wire[0:0] mux_593_nl;
  wire[0:0] nor_1285_nl;
  wire[0:0] mux_592_nl;
  wire[0:0] and_2211_nl;
  wire[0:0] mux_591_nl;
  wire[0:0] nor_1286_nl;
  wire[0:0] nor_1288_nl;
  wire[0:0] nor_1289_nl;
  wire[0:0] nor_1290_nl;
  wire[0:0] mux_595_nl;
  wire[0:0] nor_1283_nl;
  wire[0:0] nor_1284_nl;
  wire[0:0] mux_600_nl;
  wire[0:0] mux_599_nl;
  wire[0:0] and_2210_nl;
  wire[0:0] mux_598_nl;
  wire[0:0] nor_1277_nl;
  wire[0:0] nor_1279_nl;
  wire[0:0] nor_1280_nl;
  wire[0:0] nor_1281_nl;
  wire[0:0] and_738_nl;
  wire[0:0] and_739_nl;
  wire[0:0] mux_1620_nl;
  wire[0:0] or_4783_nl;
  wire[0:0] mux_1709_nl;
  wire[0:0] and_2600_nl;
  wire[0:0] mux_1713_nl;
  wire[0:0] nor_1656_nl;
  wire[0:0] or_4951_nl;
  wire[0:0] mux_610_nl;
  wire[0:0] and_2206_nl;
  wire[0:0] mux_609_nl;
  wire[0:0] mux_608_nl;
  wire[0:0] nor_1263_nl;
  wire[0:0] nor_1265_nl;
  wire[0:0] nor_1266_nl;
  wire[0:0] nor_1267_nl;
  wire[0:0] mux_612_nl;
  wire[0:0] or_1343_nl;
  wire[0:0] mux_613_nl;
  wire[0:0] or_1348_nl;
  wire[0:0] mux_614_nl;
  wire[0:0] nor_1259_nl;
  wire[0:0] nor_1260_nl;
  wire[0:0] mux_618_nl;
  wire[0:0] mux_617_nl;
  wire[0:0] nor_1253_nl;
  wire[0:0] mux_616_nl;
  wire[0:0] and_2205_nl;
  wire[0:0] mux_615_nl;
  wire[0:0] nor_1254_nl;
  wire[0:0] nor_1256_nl;
  wire[0:0] nor_1257_nl;
  wire[0:0] nor_1258_nl;
  wire[0:0] mux_619_nl;
  wire[0:0] nor_1251_nl;
  wire[0:0] nor_1252_nl;
  wire[0:0] mux_624_nl;
  wire[0:0] mux_623_nl;
  wire[0:0] and_2204_nl;
  wire[0:0] mux_622_nl;
  wire[0:0] nor_1245_nl;
  wire[0:0] nor_1247_nl;
  wire[0:0] nor_1248_nl;
  wire[0:0] nor_1249_nl;
  wire[0:0] and_743_nl;
  wire[0:0] and_744_nl;
  wire[0:0] mux_1621_nl;
  wire[0:0] or_4795_nl;
  wire[0:0] mux_1714_nl;
  wire[0:0] and_2622_nl;
  wire[0:0] mux_1718_nl;
  wire[0:0] nor_1651_nl;
  wire[0:0] or_4948_nl;
  wire[0:0] mux_634_nl;
  wire[0:0] and_2200_nl;
  wire[0:0] mux_633_nl;
  wire[0:0] mux_632_nl;
  wire[0:0] nor_1231_nl;
  wire[0:0] nor_1233_nl;
  wire[0:0] nor_1234_nl;
  wire[0:0] nor_1235_nl;
  wire[0:0] mux_636_nl;
  wire[0:0] nor_1227_nl;
  wire[0:0] nor_1228_nl;
  wire[0:0] mux_637_nl;
  wire[0:0] or_1430_nl;
  wire[0:0] mux_638_nl;
  wire[0:0] nor_1225_nl;
  wire[0:0] nor_1226_nl;
  wire[0:0] mux_642_nl;
  wire[0:0] mux_641_nl;
  wire[0:0] nor_1219_nl;
  wire[0:0] mux_640_nl;
  wire[0:0] and_2199_nl;
  wire[0:0] mux_639_nl;
  wire[0:0] nor_1220_nl;
  wire[0:0] nor_1222_nl;
  wire[0:0] nor_1223_nl;
  wire[0:0] nor_1224_nl;
  wire[0:0] mux_643_nl;
  wire[0:0] nor_1217_nl;
  wire[0:0] nor_1218_nl;
  wire[0:0] mux_648_nl;
  wire[0:0] mux_647_nl;
  wire[0:0] and_2198_nl;
  wire[0:0] mux_646_nl;
  wire[0:0] nor_1211_nl;
  wire[0:0] nor_1213_nl;
  wire[0:0] nor_1214_nl;
  wire[0:0] nor_1215_nl;
  wire[0:0] and_748_nl;
  wire[0:0] and_749_nl;
  wire[0:0] mux_1622_nl;
  wire[0:0] or_4807_nl;
  wire[0:0] mux_1719_nl;
  wire[0:0] and_2644_nl;
  wire[0:0] mux_1723_nl;
  wire[0:0] nor_1646_nl;
  wire[0:0] or_4945_nl;
  wire[0:0] mux_658_nl;
  wire[0:0] and_2194_nl;
  wire[0:0] mux_657_nl;
  wire[0:0] mux_656_nl;
  wire[0:0] nor_1197_nl;
  wire[0:0] nor_1199_nl;
  wire[0:0] nor_1200_nl;
  wire[0:0] nor_1201_nl;
  wire[0:0] mux_660_nl;
  wire[0:0] nor_1193_nl;
  wire[0:0] nor_1194_nl;
  wire[0:0] mux_661_nl;
  wire[0:0] or_1512_nl;
  wire[0:0] mux_662_nl;
  wire[0:0] nor_1191_nl;
  wire[0:0] nor_1192_nl;
  wire[0:0] mux_666_nl;
  wire[0:0] mux_665_nl;
  wire[0:0] nor_1185_nl;
  wire[0:0] mux_664_nl;
  wire[0:0] and_2193_nl;
  wire[0:0] mux_663_nl;
  wire[0:0] nor_1186_nl;
  wire[0:0] nor_1188_nl;
  wire[0:0] nor_1189_nl;
  wire[0:0] nor_1190_nl;
  wire[0:0] mux_667_nl;
  wire[0:0] nor_1183_nl;
  wire[0:0] nor_1184_nl;
  wire[0:0] mux_672_nl;
  wire[0:0] mux_671_nl;
  wire[0:0] and_2192_nl;
  wire[0:0] mux_670_nl;
  wire[0:0] nor_1177_nl;
  wire[0:0] nor_1179_nl;
  wire[0:0] nor_1180_nl;
  wire[0:0] nor_1181_nl;
  wire[0:0] and_753_nl;
  wire[0:0] and_754_nl;
  wire[0:0] mux_1623_nl;
  wire[0:0] or_4819_nl;
  wire[0:0] mux_1724_nl;
  wire[0:0] and_2666_nl;
  wire[0:0] mux_1728_nl;
  wire[0:0] nor_1641_nl;
  wire[0:0] or_4942_nl;
  wire[0:0] mux_682_nl;
  wire[0:0] and_2188_nl;
  wire[0:0] mux_681_nl;
  wire[0:0] mux_680_nl;
  wire[0:0] nor_1163_nl;
  wire[0:0] nor_1165_nl;
  wire[0:0] nor_1166_nl;
  wire[0:0] nor_1167_nl;
  wire[0:0] mux_684_nl;
  wire[0:0] or_1587_nl;
  wire[0:0] mux_685_nl;
  wire[0:0] or_1592_nl;
  wire[0:0] mux_686_nl;
  wire[0:0] nor_1159_nl;
  wire[0:0] nor_1160_nl;
  wire[0:0] mux_690_nl;
  wire[0:0] mux_689_nl;
  wire[0:0] nor_1153_nl;
  wire[0:0] mux_688_nl;
  wire[0:0] and_2187_nl;
  wire[0:0] mux_687_nl;
  wire[0:0] nor_1154_nl;
  wire[0:0] nor_1156_nl;
  wire[0:0] nor_1157_nl;
  wire[0:0] nor_1158_nl;
  wire[0:0] mux_691_nl;
  wire[0:0] nor_1151_nl;
  wire[0:0] nor_1152_nl;
  wire[0:0] mux_696_nl;
  wire[0:0] mux_695_nl;
  wire[0:0] and_2186_nl;
  wire[0:0] mux_694_nl;
  wire[0:0] nor_1145_nl;
  wire[0:0] nor_1147_nl;
  wire[0:0] nor_1148_nl;
  wire[0:0] nor_1149_nl;
  wire[0:0] and_758_nl;
  wire[0:0] and_759_nl;
  wire[0:0] mux_1624_nl;
  wire[0:0] or_4831_nl;
  wire[0:0] mux_1729_nl;
  wire[0:0] and_2688_nl;
  wire[0:0] mux_1733_nl;
  wire[0:0] nor_1636_nl;
  wire[0:0] or_4939_nl;
  wire[0:0] mux_706_nl;
  wire[0:0] and_2182_nl;
  wire[0:0] mux_705_nl;
  wire[0:0] mux_704_nl;
  wire[0:0] nor_1131_nl;
  wire[0:0] nor_1133_nl;
  wire[0:0] nor_1134_nl;
  wire[0:0] nor_1135_nl;
  wire[0:0] mux_708_nl;
  wire[0:0] or_1667_nl;
  wire[0:0] mux_709_nl;
  wire[0:0] or_1672_nl;
  wire[0:0] mux_710_nl;
  wire[0:0] nor_1127_nl;
  wire[0:0] nor_1128_nl;
  wire[0:0] mux_714_nl;
  wire[0:0] mux_713_nl;
  wire[0:0] nor_1121_nl;
  wire[0:0] mux_712_nl;
  wire[0:0] and_2181_nl;
  wire[0:0] mux_711_nl;
  wire[0:0] nor_1122_nl;
  wire[0:0] nor_1124_nl;
  wire[0:0] nor_1125_nl;
  wire[0:0] nor_1126_nl;
  wire[0:0] mux_715_nl;
  wire[0:0] nor_1119_nl;
  wire[0:0] nor_1120_nl;
  wire[0:0] mux_720_nl;
  wire[0:0] mux_719_nl;
  wire[0:0] and_2180_nl;
  wire[0:0] mux_718_nl;
  wire[0:0] nor_1113_nl;
  wire[0:0] nor_1115_nl;
  wire[0:0] nor_1116_nl;
  wire[0:0] nor_1117_nl;
  wire[0:0] and_763_nl;
  wire[0:0] and_764_nl;
  wire[0:0] mux_1625_nl;
  wire[0:0] or_4843_nl;
  wire[0:0] mux_1734_nl;
  wire[0:0] and_2710_nl;
  wire[0:0] mux_1738_nl;
  wire[0:0] nor_1631_nl;
  wire[0:0] or_4936_nl;
  wire[0:0] mux_730_nl;
  wire[0:0] and_2175_nl;
  wire[0:0] mux_729_nl;
  wire[0:0] mux_728_nl;
  wire[0:0] nor_1098_nl;
  wire[0:0] nor_1100_nl;
  wire[0:0] nor_1101_nl;
  wire[0:0] and_2176_nl;
  wire[0:0] mux_732_nl;
  wire[0:0] or_1747_nl;
  wire[0:0] mux_733_nl;
  wire[0:0] or_1752_nl;
  wire[0:0] mux_734_nl;
  wire[0:0] nor_1094_nl;
  wire[0:0] nor_1095_nl;
  wire[0:0] mux_738_nl;
  wire[0:0] mux_737_nl;
  wire[0:0] nor_1088_nl;
  wire[0:0] mux_736_nl;
  wire[0:0] and_2174_nl;
  wire[0:0] mux_735_nl;
  wire[0:0] nor_1089_nl;
  wire[0:0] nor_1091_nl;
  wire[0:0] nor_1092_nl;
  wire[0:0] nor_1093_nl;
  wire[0:0] mux_739_nl;
  wire[0:0] nor_1086_nl;
  wire[0:0] nor_1087_nl;
  wire[0:0] mux_744_nl;
  wire[0:0] mux_743_nl;
  wire[0:0] and_2173_nl;
  wire[0:0] mux_742_nl;
  wire[0:0] nor_1080_nl;
  wire[0:0] nor_1082_nl;
  wire[0:0] nor_1083_nl;
  wire[0:0] nor_1084_nl;
  wire[0:0] and_768_nl;
  wire[0:0] and_769_nl;
  wire[0:0] mux_1626_nl;
  wire[0:0] mux_1739_nl;
  wire[0:0] or_4854_nl;
  wire[0:0] mux_1740_nl;
  wire[0:0] and_2732_nl;
  wire[0:0] mux_1745_nl;
  wire[0:0] nor_1627_nl;
  wire[0:0] or_4935_nl;
  wire[0:0] mux_754_nl;
  wire[0:0] and_2166_nl;
  wire[0:0] mux_753_nl;
  wire[0:0] mux_752_nl;
  wire[0:0] nor_1065_nl;
  wire[0:0] nor_1067_nl;
  wire[0:0] nor_1068_nl;
  wire[0:0] and_2167_nl;
  wire[0:0] mux_759_nl;
  wire[0:0] or_1830_nl;
  wire[0:0] mux_758_nl;
  wire[0:0] mux_760_nl;
  wire[0:0] or_1835_nl;
  wire[0:0] mux_761_nl;
  wire[0:0] nor_1063_nl;
  wire[0:0] nor_1064_nl;
  wire[0:0] mux_765_nl;
  wire[0:0] mux_764_nl;
  wire[0:0] nor_1057_nl;
  wire[0:0] mux_763_nl;
  wire[0:0] and_2165_nl;
  wire[0:0] mux_762_nl;
  wire[0:0] nor_1058_nl;
  wire[0:0] nor_1060_nl;
  wire[0:0] nor_1061_nl;
  wire[0:0] nor_1062_nl;
  wire[0:0] mux_766_nl;
  wire[0:0] nor_1055_nl;
  wire[0:0] nor_1056_nl;
  wire[0:0] mux_770_nl;
  wire[0:0] mux_769_nl;
  wire[0:0] and_2164_nl;
  wire[0:0] mux_768_nl;
  wire[0:0] nor_1049_nl;
  wire[0:0] nor_1051_nl;
  wire[0:0] nor_1052_nl;
  wire[0:0] nor_1053_nl;
  wire[0:0] and_773_nl;
  wire[0:0] and_774_nl;
  wire[0:0] mux_1627_nl;
  wire[0:0] or_4865_nl;
  wire[0:0] mux_1746_nl;
  wire[0:0] and_2754_nl;
  wire[0:0] mux_1750_nl;
  wire[0:0] nor_1622_nl;
  wire[0:0] or_4932_nl;
  wire[0:0] mux_781_nl;
  wire[0:0] and_2160_nl;
  wire[0:0] mux_780_nl;
  wire[0:0] mux_779_nl;
  wire[0:0] nor_1032_nl;
  wire[0:0] nor_1034_nl;
  wire[0:0] nor_1035_nl;
  wire[0:0] and_2161_nl;
  wire[0:0] mux_785_nl;
  wire[0:0] or_1905_nl;
  wire[0:0] mux_784_nl;
  wire[0:0] or_1908_nl;
  wire[0:0] mux_786_nl;
  wire[0:0] or_1913_nl;
  wire[0:0] mux_787_nl;
  wire[0:0] nor_1030_nl;
  wire[0:0] nor_1031_nl;
  wire[0:0] mux_791_nl;
  wire[0:0] mux_790_nl;
  wire[0:0] nor_1024_nl;
  wire[0:0] mux_789_nl;
  wire[0:0] and_2159_nl;
  wire[0:0] mux_788_nl;
  wire[0:0] nor_1025_nl;
  wire[0:0] nor_1027_nl;
  wire[0:0] nor_1028_nl;
  wire[0:0] nor_1029_nl;
  wire[0:0] mux_792_nl;
  wire[0:0] nor_1022_nl;
  wire[0:0] nor_1023_nl;
  wire[0:0] mux_797_nl;
  wire[0:0] mux_796_nl;
  wire[0:0] and_2158_nl;
  wire[0:0] mux_795_nl;
  wire[0:0] nor_1016_nl;
  wire[0:0] nor_1018_nl;
  wire[0:0] nor_1019_nl;
  wire[0:0] nor_1020_nl;
  wire[0:0] and_778_nl;
  wire[0:0] and_779_nl;
  wire[0:0] mux_1628_nl;
  wire[0:0] or_4877_nl;
  wire[0:0] mux_1751_nl;
  wire[0:0] and_2776_nl;
  wire[0:0] mux_1755_nl;
  wire[0:0] nor_1617_nl;
  wire[0:0] or_4929_nl;
  wire[0:0] mux_808_nl;
  wire[0:0] and_2154_nl;
  wire[0:0] mux_807_nl;
  wire[0:0] mux_806_nl;
  wire[0:0] nor_999_nl;
  wire[0:0] nor_1001_nl;
  wire[0:0] nor_1002_nl;
  wire[0:0] and_2155_nl;
  wire[0:0] mux_812_nl;
  wire[0:0] or_1988_nl;
  wire[0:0] mux_811_nl;
  wire[0:0] or_1991_nl;
  wire[0:0] mux_813_nl;
  wire[0:0] or_1996_nl;
  wire[0:0] mux_814_nl;
  wire[0:0] nor_997_nl;
  wire[0:0] nor_998_nl;
  wire[0:0] mux_818_nl;
  wire[0:0] mux_817_nl;
  wire[0:0] nor_991_nl;
  wire[0:0] mux_816_nl;
  wire[0:0] and_2153_nl;
  wire[0:0] mux_815_nl;
  wire[0:0] nor_992_nl;
  wire[0:0] nor_994_nl;
  wire[0:0] nor_995_nl;
  wire[0:0] nor_996_nl;
  wire[0:0] mux_819_nl;
  wire[0:0] nor_989_nl;
  wire[0:0] nor_990_nl;
  wire[0:0] mux_824_nl;
  wire[0:0] mux_823_nl;
  wire[0:0] and_2152_nl;
  wire[0:0] mux_822_nl;
  wire[0:0] nor_983_nl;
  wire[0:0] nor_985_nl;
  wire[0:0] nor_986_nl;
  wire[0:0] nor_987_nl;
  wire[0:0] and_783_nl;
  wire[0:0] and_784_nl;
  wire[0:0] mux_1629_nl;
  wire[0:0] mux_1756_nl;
  wire[0:0] or_4888_nl;
  wire[0:0] mux_1757_nl;
  wire[0:0] and_2798_nl;
  wire[0:0] mux_1762_nl;
  wire[0:0] nor_1612_nl;
  wire[0:0] or_4928_nl;
  wire[0:0] mux_835_nl;
  wire[0:0] and_2149_nl;
  wire[0:0] mux_834_nl;
  wire[0:0] mux_833_nl;
  wire[0:0] nor_967_nl;
  wire[0:0] nor_969_nl;
  wire[0:0] nor_970_nl;
  wire[0:0] and_2150_nl;
  wire[0:0] mux_837_nl;
  wire[0:0] nor_963_nl;
  wire[0:0] nor_964_nl;
  wire[0:0] mux_838_nl;
  wire[0:0] or_2082_nl;
  wire[0:0] mux_839_nl;
  wire[0:0] nor_961_nl;
  wire[0:0] nor_962_nl;
  wire[0:0] mux_843_nl;
  wire[0:0] mux_842_nl;
  wire[0:0] nor_955_nl;
  wire[0:0] mux_841_nl;
  wire[0:0] and_2148_nl;
  wire[0:0] mux_840_nl;
  wire[0:0] nor_956_nl;
  wire[0:0] nor_958_nl;
  wire[0:0] nor_959_nl;
  wire[0:0] nor_960_nl;
  wire[0:0] mux_844_nl;
  wire[0:0] nor_953_nl;
  wire[0:0] nor_954_nl;
  wire[0:0] mux_849_nl;
  wire[0:0] mux_848_nl;
  wire[0:0] and_2147_nl;
  wire[0:0] mux_847_nl;
  wire[0:0] nor_947_nl;
  wire[0:0] nor_949_nl;
  wire[0:0] nor_950_nl;
  wire[0:0] nor_951_nl;
  wire[0:0] and_788_nl;
  wire[0:0] and_789_nl;
  wire[0:0] mux_1630_nl;
  wire[0:0] or_4900_nl;
  wire[0:0] mux_1763_nl;
  wire[0:0] and_2819_nl;
  wire[0:0] mux_1767_nl;
  wire[0:0] nor_1607_nl;
  wire[0:0] or_4925_nl;
  wire[0:0] mux_860_nl;
  wire[0:0] and_2143_nl;
  wire[0:0] mux_859_nl;
  wire[0:0] mux_858_nl;
  wire[0:0] nor_930_nl;
  wire[0:0] nor_932_nl;
  wire[0:0] nor_933_nl;
  wire[0:0] and_2144_nl;
  wire[0:0] mux_862_nl;
  wire[0:0] nor_926_nl;
  wire[0:0] nor_927_nl;
  wire[0:0] mux_863_nl;
  wire[0:0] or_2162_nl;
  wire[0:0] mux_864_nl;
  wire[0:0] nor_924_nl;
  wire[0:0] nor_925_nl;
  wire[0:0] mux_868_nl;
  wire[0:0] mux_867_nl;
  wire[0:0] nor_918_nl;
  wire[0:0] mux_866_nl;
  wire[0:0] and_2142_nl;
  wire[0:0] mux_865_nl;
  wire[0:0] nor_919_nl;
  wire[0:0] nor_921_nl;
  wire[0:0] nor_922_nl;
  wire[0:0] nor_923_nl;
  wire[0:0] mux_869_nl;
  wire[0:0] nor_916_nl;
  wire[0:0] nor_917_nl;
  wire[0:0] mux_874_nl;
  wire[0:0] mux_873_nl;
  wire[0:0] and_2141_nl;
  wire[0:0] mux_872_nl;
  wire[0:0] nor_910_nl;
  wire[0:0] nor_912_nl;
  wire[0:0] nor_913_nl;
  wire[0:0] nor_914_nl;
  wire[0:0] and_793_nl;
  wire[0:0] and_794_nl;
  wire[0:0] mux_1631_nl;
  wire[0:0] or_4912_nl;
  wire[0:0] mux_1768_nl;
  wire[0:0] and_2841_nl;
  wire[0:0] mux_1772_nl;
  wire[0:0] nor_1602_nl;
  wire[0:0] or_4922_nl;
  wire[0:0] mux_885_nl;
  wire[0:0] and_2137_nl;
  wire[0:0] mux_884_nl;
  wire[0:0] mux_883_nl;
  wire[0:0] nor_893_nl;
  wire[0:0] nor_895_nl;
  wire[0:0] nor_896_nl;
  wire[0:0] and_2138_nl;
  wire[0:0] mux_887_nl;
  wire[0:0] or_2237_nl;
  wire[0:0] mux_888_nl;
  wire[0:0] or_2242_nl;
  wire[0:0] mux_889_nl;
  wire[0:0] nor_889_nl;
  wire[0:0] nor_890_nl;
  wire[0:0] mux_893_nl;
  wire[0:0] mux_892_nl;
  wire[0:0] nor_883_nl;
  wire[0:0] mux_891_nl;
  wire[0:0] and_2136_nl;
  wire[0:0] mux_890_nl;
  wire[0:0] nor_884_nl;
  wire[0:0] nor_886_nl;
  wire[0:0] nor_887_nl;
  wire[0:0] nor_888_nl;
  wire[0:0] mux_894_nl;
  wire[0:0] nor_881_nl;
  wire[0:0] nor_882_nl;
  wire[0:0] mux_899_nl;
  wire[0:0] mux_898_nl;
  wire[0:0] and_2135_nl;
  wire[0:0] mux_897_nl;
  wire[0:0] nor_875_nl;
  wire[0:0] nor_877_nl;
  wire[0:0] nor_878_nl;
  wire[0:0] nor_879_nl;
  wire[0:0] mux_900_nl;
  wire[0:0] or_2278_nl;
  wire[0:0] mux_902_nl;
  wire[0:0] mux_901_nl;
  wire[0:0] or_2282_nl;
  wire[0:0] nor_873_nl;
  wire[0:0] mux_905_nl;
  wire[0:0] mux_904_nl;
  wire[0:0] and_323_nl;
  wire[0:0] mux_903_nl;
  wire[0:0] or_2286_nl;
  wire[0:0] mux_907_nl;
  wire[0:0] mux_906_nl;
  wire[0:0] or_2293_nl;
  wire[0:0] nor_870_nl;
  wire[0:0] mux_910_nl;
  wire[0:0] mux_909_nl;
  wire[0:0] and_324_nl;
  wire[0:0] mux_908_nl;
  wire[0:0] or_2297_nl;
  wire[0:0] mux_912_nl;
  wire[0:0] mux_911_nl;
  wire[0:0] or_2304_nl;
  wire[0:0] nor_867_nl;
  wire[0:0] mux_915_nl;
  wire[0:0] mux_914_nl;
  wire[0:0] and_325_nl;
  wire[0:0] mux_913_nl;
  wire[0:0] or_2308_nl;
  wire[0:0] mux_917_nl;
  wire[0:0] mux_916_nl;
  wire[0:0] or_2317_nl;
  wire[0:0] nor_865_nl;
  wire[0:0] mux_920_nl;
  wire[0:0] mux_919_nl;
  wire[0:0] and_326_nl;
  wire[0:0] mux_918_nl;
  wire[0:0] or_2318_nl;
  wire[0:0] mux_922_nl;
  wire[0:0] mux_921_nl;
  wire[0:0] or_2325_nl;
  wire[0:0] nor_863_nl;
  wire[0:0] mux_925_nl;
  wire[0:0] mux_924_nl;
  wire[0:0] and_327_nl;
  wire[0:0] mux_923_nl;
  wire[0:0] or_2329_nl;
  wire[0:0] mux_927_nl;
  wire[0:0] mux_926_nl;
  wire[0:0] or_2336_nl;
  wire[0:0] nor_860_nl;
  wire[0:0] mux_932_nl;
  wire[0:0] mux_931_nl;
  wire[0:0] mux_930_nl;
  wire[0:0] mux_928_nl;
  wire[0:0] nor_385_nl;
  wire[0:0] mux_929_nl;
  wire[0:0] mux_934_nl;
  wire[0:0] mux_933_nl;
  wire[0:0] or_2347_nl;
  wire[0:0] nor_857_nl;
  wire[0:0] mux_937_nl;
  wire[0:0] mux_936_nl;
  wire[0:0] and_329_nl;
  wire[0:0] mux_935_nl;
  wire[0:0] or_2351_nl;
  wire[0:0] mux_939_nl;
  wire[0:0] mux_938_nl;
  wire[0:0] or_2358_nl;
  wire[0:0] nor_854_nl;
  wire[0:0] mux_942_nl;
  wire[0:0] mux_941_nl;
  wire[0:0] and_330_nl;
  wire[0:0] mux_940_nl;
  wire[0:0] or_2362_nl;
  wire[0:0] mux_944_nl;
  wire[0:0] mux_943_nl;
  wire[0:0] or_2369_nl;
  wire[0:0] nor_851_nl;
  wire[0:0] mux_947_nl;
  wire[0:0] mux_946_nl;
  wire[0:0] and_331_nl;
  wire[0:0] mux_945_nl;
  wire[0:0] or_2373_nl;
  wire[0:0] mux_949_nl;
  wire[0:0] mux_948_nl;
  wire[0:0] or_2380_nl;
  wire[0:0] nor_848_nl;
  wire[0:0] mux_954_nl;
  wire[0:0] mux_953_nl;
  wire[0:0] mux_952_nl;
  wire[0:0] mux_950_nl;
  wire[0:0] nor_392_nl;
  wire[0:0] mux_951_nl;
  wire[0:0] mux_956_nl;
  wire[0:0] mux_955_nl;
  wire[0:0] or_2391_nl;
  wire[0:0] nor_846_nl;
  wire[0:0] mux_959_nl;
  wire[0:0] mux_958_nl;
  wire[0:0] and_333_nl;
  wire[0:0] mux_957_nl;
  wire[0:0] or_4652_nl;
  wire[0:0] or_2392_nl;
  wire[0:0] mux_961_nl;
  wire[0:0] mux_960_nl;
  wire[0:0] or_2400_nl;
  wire[0:0] and_2132_nl;
  wire[0:0] or_2396_nl;
  wire[0:0] mux_964_nl;
  wire[0:0] mux_963_nl;
  wire[0:0] and_334_nl;
  wire[0:0] mux_962_nl;
  wire[0:0] or_2401_nl;
  wire[0:0] mux_966_nl;
  wire[0:0] mux_965_nl;
  wire[0:0] or_2409_nl;
  wire[0:0] and_2131_nl;
  wire[0:0] or_2405_nl;
  wire[0:0] mux_969_nl;
  wire[0:0] mux_968_nl;
  wire[0:0] and_335_nl;
  wire[0:0] mux_967_nl;
  wire[0:0] or_2410_nl;
  wire[0:0] mux_971_nl;
  wire[0:0] mux_970_nl;
  wire[0:0] or_2417_nl;
  wire[0:0] nor_844_nl;
  wire[0:0] mux_974_nl;
  wire[0:0] mux_973_nl;
  wire[0:0] and_336_nl;
  wire[0:0] mux_972_nl;
  wire[0:0] or_2423_nl;
  wire[0:0] or_2421_nl;
  wire[0:0] mux_976_nl;
  wire[0:0] mux_975_nl;
  wire[0:0] or_2428_nl;
  wire[0:0] nor_841_nl;
  wire[0:0] mux_979_nl;
  wire[0:0] mux_978_nl;
  wire[0:0] and_337_nl;
  wire[0:0] mux_977_nl;
  wire[0:0] or_2432_nl;
  wire[0:0] mux_982_nl;
  wire[0:0] mux_981_nl;
  wire[0:0] mux_980_nl;
  wire[0:0] or_2439_nl;
  wire[0:0] nor_899_nl;
  wire[0:0] mux_985_nl;
  wire[0:0] mux_984_nl;
  wire[0:0] and_338_nl;
  wire[0:0] mux_983_nl;
  wire[0:0] or_2442_nl;
  wire[0:0] mux_992_nl;
  wire[0:0] mux_991_nl;
  wire[0:0] mux_989_nl;
  wire[0:0] mux_988_nl;
  wire[0:0] mux_987_nl;
  wire[0:0] mux_990_nl;
  wire[0:0] or_2453_nl;
  wire[0:0] mux_999_nl;
  wire[0:0] mux_998_nl;
  wire[0:0] mux_996_nl;
  wire[0:0] mux_995_nl;
  wire[0:0] mux_994_nl;
  wire[0:0] mux_997_nl;
  wire[0:0] or_2461_nl;
  wire[0:0] mux_1008_nl;
  wire[0:0] mux_1006_nl;
  wire[0:0] mux_1005_nl;
  wire[0:0] mux_1003_nl;
  wire[0:0] mux_1002_nl;
  wire[0:0] mux_1001_nl;
  wire[0:0] mux_1004_nl;
  wire[0:0] mux_1007_nl;
  wire[0:0] nor_838_nl;
  wire[0:0] or_2467_nl;
  wire[0:0] mux_1017_nl;
  wire[0:0] mux_1015_nl;
  wire[0:0] mux_1014_nl;
  wire[0:0] mux_1012_nl;
  wire[0:0] mux_1011_nl;
  wire[0:0] mux_1010_nl;
  wire[0:0] mux_1013_nl;
  wire[0:0] mux_1016_nl;
  wire[0:0] nor_837_nl;
  wire[0:0] or_2475_nl;
  wire[0:0] mux_1026_nl;
  wire[0:0] mux_1024_nl;
  wire[0:0] mux_1023_nl;
  wire[0:0] mux_1021_nl;
  wire[0:0] mux_1020_nl;
  wire[0:0] mux_1019_nl;
  wire[0:0] mux_1022_nl;
  wire[0:0] mux_1025_nl;
  wire[0:0] nor_836_nl;
  wire[0:0] or_2483_nl;
  wire[0:0] mux_1035_nl;
  wire[0:0] mux_1033_nl;
  wire[0:0] mux_1032_nl;
  wire[0:0] mux_1030_nl;
  wire[0:0] mux_1029_nl;
  wire[0:0] mux_1028_nl;
  wire[0:0] mux_1031_nl;
  wire[0:0] mux_1034_nl;
  wire[0:0] nor_835_nl;
  wire[0:0] or_2491_nl;
  wire[0:0] mux_1044_nl;
  wire[0:0] mux_1042_nl;
  wire[0:0] mux_1041_nl;
  wire[0:0] mux_1039_nl;
  wire[0:0] mux_1038_nl;
  wire[0:0] mux_1037_nl;
  wire[0:0] mux_1040_nl;
  wire[0:0] mux_1043_nl;
  wire[0:0] nor_834_nl;
  wire[0:0] or_2499_nl;
  wire[0:0] mux_1051_nl;
  wire[0:0] mux_1050_nl;
  wire[0:0] mux_1048_nl;
  wire[0:0] mux_1047_nl;
  wire[0:0] mux_1046_nl;
  wire[0:0] mux_1049_nl;
  wire[0:0] or_2509_nl;
  wire[0:0] mux_1060_nl;
  wire[0:0] mux_1058_nl;
  wire[0:0] mux_1057_nl;
  wire[0:0] mux_1055_nl;
  wire[0:0] mux_1054_nl;
  wire[0:0] mux_1053_nl;
  wire[0:0] mux_1056_nl;
  wire[0:0] mux_1059_nl;
  wire[0:0] nor_833_nl;
  wire[0:0] or_2515_nl;
  wire[0:0] mux_1069_nl;
  wire[0:0] mux_1067_nl;
  wire[0:0] mux_1066_nl;
  wire[0:0] mux_1064_nl;
  wire[0:0] mux_1063_nl;
  wire[0:0] mux_1062_nl;
  wire[0:0] mux_1065_nl;
  wire[0:0] mux_1068_nl;
  wire[0:0] nor_832_nl;
  wire[0:0] or_2523_nl;
  wire[0:0] mux_1078_nl;
  wire[0:0] mux_1076_nl;
  wire[0:0] mux_1075_nl;
  wire[0:0] mux_1073_nl;
  wire[0:0] mux_1072_nl;
  wire[0:0] mux_1071_nl;
  wire[0:0] mux_1074_nl;
  wire[0:0] mux_1077_nl;
  wire[0:0] nor_831_nl;
  wire[0:0] or_2531_nl;
  wire[0:0] mux_1087_nl;
  wire[0:0] mux_1085_nl;
  wire[0:0] mux_1084_nl;
  wire[0:0] mux_1082_nl;
  wire[0:0] mux_1081_nl;
  wire[0:0] mux_1080_nl;
  wire[0:0] mux_1083_nl;
  wire[0:0] mux_1086_nl;
  wire[0:0] nor_830_nl;
  wire[0:0] or_2539_nl;
  wire[0:0] mux_1096_nl;
  wire[0:0] mux_1094_nl;
  wire[0:0] mux_1093_nl;
  wire[0:0] mux_1091_nl;
  wire[0:0] mux_1090_nl;
  wire[0:0] mux_1089_nl;
  wire[0:0] mux_1092_nl;
  wire[0:0] mux_1095_nl;
  wire[0:0] nor_829_nl;
  wire[0:0] or_2547_nl;
  wire[0:0] mux_1105_nl;
  wire[0:0] mux_1103_nl;
  wire[0:0] mux_1102_nl;
  wire[0:0] mux_1100_nl;
  wire[0:0] mux_1099_nl;
  wire[0:0] mux_1098_nl;
  wire[0:0] mux_1101_nl;
  wire[0:0] mux_1104_nl;
  wire[0:0] nor_828_nl;
  wire[0:0] or_2555_nl;
  wire[0:0] mux_1114_nl;
  wire[0:0] mux_1112_nl;
  wire[0:0] mux_1111_nl;
  wire[0:0] mux_1109_nl;
  wire[0:0] mux_1108_nl;
  wire[0:0] mux_1107_nl;
  wire[0:0] mux_1110_nl;
  wire[0:0] mux_1113_nl;
  wire[0:0] nor_827_nl;
  wire[0:0] or_2563_nl;
  wire[0:0] mux_1122_nl;
  wire[0:0] mux_1120_nl;
  wire[0:0] mux_1118_nl;
  wire[0:0] mux_1117_nl;
  wire[0:0] mux_1115_nl;
  wire[0:0] mux_1116_nl;
  wire[0:0] or_2570_nl;
  wire[0:0] mux_1119_nl;
  wire[0:0] or_2571_nl;
  wire[0:0] mux_1121_nl;
  wire[0:0] nor_826_nl;
  wire[0:0] or_2572_nl;
  wire[0:0] nor_825_nl;
  wire[0:0] mux_1140_nl;
  wire[0:0] mux_1139_nl;
  wire[0:0] mux_1137_nl;
  wire[0:0] mux_1124_nl;
  wire[0:0] mux_1123_nl;
  wire[0:0] mux_1136_nl;
  wire[0:0] mux_1132_nl;
  wire[0:0] mux_1128_nl;
  wire[0:0] mux_1131_nl;
  wire[0:0] and_344_nl;
  wire[0:0] nor_824_nl;
  wire[0:0] mux_1135_nl;
  wire[0:0] mux_1144_nl;
  wire[0:0] mux_1143_nl;
  wire[0:0] nand_133_nl;
  wire[0:0] and_2129_nl;
  wire[0:0] mux_1142_nl;
  wire[0:0] nor_822_nl;
  wire[0:0] nor_818_nl;
  wire[0:0] mux_1162_nl;
  wire[0:0] mux_1161_nl;
  wire[0:0] mux_1159_nl;
  wire[0:0] mux_1146_nl;
  wire[0:0] mux_1145_nl;
  wire[0:0] mux_1158_nl;
  wire[0:0] mux_1154_nl;
  wire[0:0] mux_1150_nl;
  wire[0:0] mux_1153_nl;
  wire[0:0] and_348_nl;
  wire[0:0] nor_817_nl;
  wire[0:0] mux_1157_nl;
  wire[0:0] and_2128_nl;
  wire[0:0] mux_1167_nl;
  wire[0:0] mux_1166_nl;
  wire[0:0] mux_1165_nl;
  wire[0:0] mux_1164_nl;
  wire[0:0] and_350_nl;
  wire[0:0] nor_816_nl;
  wire[0:0] mux_1185_nl;
  wire[0:0] mux_1184_nl;
  wire[0:0] mux_1182_nl;
  wire[0:0] mux_1169_nl;
  wire[0:0] mux_1168_nl;
  wire[0:0] mux_1181_nl;
  wire[0:0] mux_1177_nl;
  wire[0:0] mux_1173_nl;
  wire[0:0] mux_1176_nl;
  wire[0:0] and_353_nl;
  wire[0:0] nor_815_nl;
  wire[0:0] mux_1180_nl;
  wire[0:0] and_2127_nl;
  wire[0:0] mux_1189_nl;
  wire[0:0] mux_1188_nl;
  wire[0:0] nand_135_nl;
  wire[0:0] and_2126_nl;
  wire[0:0] mux_1187_nl;
  wire[0:0] nor_813_nl;
  wire[0:0] mux_1194_nl;
  wire[0:0] mux_1193_nl;
  wire[0:0] or_2667_nl;
  wire[0:0] nor_808_nl;
  wire[0:0] mux_1192_nl;
  wire[0:0] or_2672_nl;
  wire[0:0] nor_806_nl;
  wire[0:0] mux_1212_nl;
  wire[0:0] mux_1211_nl;
  wire[0:0] mux_1209_nl;
  wire[0:0] mux_1196_nl;
  wire[0:0] mux_1195_nl;
  wire[0:0] mux_1208_nl;
  wire[0:0] mux_1204_nl;
  wire[0:0] mux_1200_nl;
  wire[0:0] mux_1203_nl;
  wire[0:0] and_357_nl;
  wire[0:0] nor_805_nl;
  wire[0:0] mux_1207_nl;
  wire[0:0] and_2125_nl;
  wire[0:0] mux_1218_nl;
  wire[0:0] mux_1217_nl;
  wire[0:0] mux_1216_nl;
  wire[0:0] mux_1214_nl;
  wire[0:0] and_359_nl;
  wire[0:0] mux_1223_nl;
  wire[0:0] mux_1222_nl;
  wire[0:0] or_2701_nl;
  wire[0:0] nor_803_nl;
  wire[0:0] mux_1221_nl;
  wire[0:0] or_2706_nl;
  wire[0:0] mux_1228_nl;
  wire[0:0] mux_1227_nl;
  wire[0:0] or_2714_nl;
  wire[0:0] nor_800_nl;
  wire[0:0] mux_1226_nl;
  wire[0:0] or_2719_nl;
  wire[0:0] nor_798_nl;
  wire[0:0] mux_1246_nl;
  wire[0:0] mux_1245_nl;
  wire[0:0] mux_1243_nl;
  wire[0:0] mux_1230_nl;
  wire[0:0] mux_1229_nl;
  wire[0:0] mux_1242_nl;
  wire[0:0] mux_1238_nl;
  wire[0:0] mux_1234_nl;
  wire[0:0] mux_1237_nl;
  wire[0:0] and_362_nl;
  wire[0:0] nor_797_nl;
  wire[0:0] mux_1241_nl;
  wire[0:0] and_2124_nl;
  wire[0:0] mux_1251_nl;
  wire[0:0] mux_1250_nl;
  wire[0:0] mux_1249_nl;
  wire[0:0] mux_1248_nl;
  wire[0:0] and_364_nl;
  wire[0:0] nor_796_nl;
  wire[0:0] mux_1269_nl;
  wire[0:0] mux_1268_nl;
  wire[0:0] mux_1266_nl;
  wire[0:0] mux_1253_nl;
  wire[0:0] mux_1252_nl;
  wire[0:0] mux_1265_nl;
  wire[0:0] mux_1261_nl;
  wire[0:0] mux_1257_nl;
  wire[0:0] mux_1260_nl;
  wire[0:0] and_367_nl;
  wire[0:0] nor_795_nl;
  wire[0:0] mux_1264_nl;
  wire[0:0] and_2123_nl;
  wire[0:0] mux_1275_nl;
  wire[0:0] mux_1274_nl;
  wire[0:0] mux_1273_nl;
  wire[0:0] mux_1271_nl;
  wire[0:0] and_369_nl;
  wire[0:0] mux_1280_nl;
  wire[0:0] mux_1279_nl;
  wire[0:0] mux_1278_nl;
  wire[0:0] mux_1277_nl;
  wire[0:0] or_2769_nl;
  wire[0:0] mux_1285_nl;
  wire[0:0] mux_1284_nl;
  wire[0:0] or_2777_nl;
  wire[0:0] nor_793_nl;
  wire[0:0] mux_1283_nl;
  wire[0:0] or_2782_nl;
  wire[0:0] mux_1290_nl;
  wire[0:0] mux_1289_nl;
  wire[0:0] or_2790_nl;
  wire[0:0] nor_790_nl;
  wire[0:0] mux_1288_nl;
  wire[0:0] or_2795_nl;
  wire[0:0] nor_788_nl;
  wire[0:0] mux_1308_nl;
  wire[0:0] mux_1307_nl;
  wire[0:0] mux_1305_nl;
  wire[0:0] mux_1292_nl;
  wire[0:0] mux_1291_nl;
  wire[0:0] mux_1304_nl;
  wire[0:0] mux_1300_nl;
  wire[0:0] mux_1296_nl;
  wire[0:0] mux_1299_nl;
  wire[0:0] and_372_nl;
  wire[0:0] nor_787_nl;
  wire[0:0] mux_1303_nl;
  wire[0:0] and_2122_nl;
  wire[0:0] mux_1313_nl;
  wire[0:0] mux_1312_nl;
  wire[0:0] mux_1311_nl;
  wire[0:0] mux_1310_nl;
  wire[0:0] and_374_nl;
  wire[0:0] mux_1318_nl;
  wire[0:0] mux_1317_nl;
  wire[0:0] or_2826_nl;
  wire[0:0] nor_785_nl;
  wire[0:0] mux_1316_nl;
  wire[0:0] or_2831_nl;
  wire[0:0] nor_783_nl;
  wire[0:0] mux_1336_nl;
  wire[0:0] mux_1335_nl;
  wire[0:0] mux_1333_nl;
  wire[0:0] mux_1320_nl;
  wire[0:0] mux_1319_nl;
  wire[0:0] mux_1332_nl;
  wire[0:0] mux_1328_nl;
  wire[0:0] mux_1324_nl;
  wire[0:0] mux_1327_nl;
  wire[0:0] and_377_nl;
  wire[0:0] nor_782_nl;
  wire[0:0] mux_1331_nl;
  wire[0:0] and_2121_nl;
  wire[0:0] mux_1340_nl;
  wire[0:0] mux_1339_nl;
  wire[0:0] nand_143_nl;
  wire[0:0] and_2120_nl;
  wire[0:0] mux_1338_nl;
  wire[0:0] nor_780_nl;
  wire[0:0] nor_776_nl;
  wire[0:0] mux_1358_nl;
  wire[0:0] mux_1357_nl;
  wire[0:0] mux_1355_nl;
  wire[0:0] mux_1342_nl;
  wire[0:0] mux_1341_nl;
  wire[0:0] mux_1354_nl;
  wire[0:0] mux_1350_nl;
  wire[0:0] mux_1346_nl;
  wire[0:0] mux_1349_nl;
  wire[0:0] and_381_nl;
  wire[0:0] nor_775_nl;
  wire[0:0] mux_1353_nl;
  wire[0:0] and_2119_nl;
  wire[0:0] mux_1363_nl;
  wire[0:0] mux_1362_nl;
  wire[0:0] mux_1361_nl;
  wire[0:0] mux_1360_nl;
  wire[0:0] and_383_nl;
  wire[0:0] mux_1446_nl;
  wire[0:0] or_2967_nl;
  wire[0:0] mux_1447_nl;
  wire[0:0] or_2970_nl;
  wire[0:0] mux_1448_nl;
  wire[0:0] or_2973_nl;
  wire[0:0] mux_1449_nl;
  wire[0:0] or_2976_nl;
  wire[0:0] mux_1450_nl;
  wire[0:0] or_2979_nl;
  wire[0:0] mux_1452_nl;
  wire[0:0] or_2984_nl;
  wire[0:0] mux_1453_nl;
  wire[0:0] or_2987_nl;
  wire[0:0] mux_1454_nl;
  wire[0:0] or_2990_nl;
  wire[0:0] mux_1456_nl;
  wire[0:0] or_2995_nl;
  wire[0:0] mux_1457_nl;
  wire[0:0] or_2998_nl;
  wire[0:0] mux_1458_nl;
  wire[0:0] or_3001_nl;
  wire[0:0] mux_1460_nl;
  wire[0:0] or_3006_nl;
  wire[0:0] mux_1461_nl;
  wire[0:0] or_3009_nl;
  wire[0:0] mux_1462_nl;
  wire[0:0] or_3012_nl;
  wire[0:0] mux_1464_nl;
  wire[0:0] or_3017_nl;
  wire[0:0] mux_1465_nl;
  wire[0:0] or_3020_nl;
  wire[0:0] mux_1466_nl;
  wire[0:0] or_3023_nl;
  wire[0:0] mux_1468_nl;
  wire[0:0] or_3028_nl;
  wire[0:0] mux_1469_nl;
  wire[0:0] or_3031_nl;
  wire[0:0] mux_1470_nl;
  wire[0:0] or_3034_nl;
  wire[0:0] mux_1472_nl;
  wire[0:0] or_3039_nl;
  wire[0:0] mux_1473_nl;
  wire[0:0] or_3042_nl;
  wire[0:0] mux_1474_nl;
  wire[0:0] or_3045_nl;
  wire[0:0] mux_1476_nl;
  wire[0:0] or_3050_nl;
  wire[0:0] mux_1477_nl;
  wire[0:0] or_3053_nl;
  wire[0:0] mux_1478_nl;
  wire[0:0] or_3056_nl;
  wire[0:0] mux_1480_nl;
  wire[0:0] or_3061_nl;
  wire[0:0] mux_1481_nl;
  wire[0:0] or_3064_nl;
  wire[0:0] mux_1482_nl;
  wire[0:0] or_3067_nl;
  wire[0:0] mux_1484_nl;
  wire[0:0] or_3072_nl;
  wire[0:0] mux_1485_nl;
  wire[0:0] or_3075_nl;
  wire[0:0] mux_1486_nl;
  wire[0:0] or_3078_nl;
  wire[0:0] mux_1488_nl;
  wire[0:0] or_3083_nl;
  wire[0:0] mux_1489_nl;
  wire[0:0] or_3086_nl;
  wire[0:0] mux_1490_nl;
  wire[0:0] or_3089_nl;
  wire[0:0] mux_1492_nl;
  wire[0:0] or_3094_nl;
  wire[0:0] mux_1493_nl;
  wire[0:0] or_3097_nl;
  wire[0:0] mux_1494_nl;
  wire[0:0] or_3100_nl;
  wire[0:0] mux_1496_nl;
  wire[0:0] or_3105_nl;
  wire[0:0] mux_1497_nl;
  wire[0:0] or_3108_nl;
  wire[0:0] mux_1498_nl;
  wire[0:0] or_3111_nl;
  wire[0:0] mux_1500_nl;
  wire[0:0] or_3116_nl;
  wire[0:0] mux_1501_nl;
  wire[0:0] or_3119_nl;
  wire[0:0] mux_1502_nl;
  wire[0:0] or_3122_nl;
  wire[0:0] mux_1504_nl;
  wire[0:0] or_3127_nl;
  wire[0:0] mux_1505_nl;
  wire[0:0] or_3130_nl;
  wire[0:0] mux_1506_nl;
  wire[0:0] or_3133_nl;
  wire[0:0] mux_1508_nl;
  wire[0:0] or_3138_nl;
  wire[0:0] mux_1510_nl;
  wire[0:0] or_3143_nl;
  wire[0:0] mux_1513_nl;
  wire[0:0] or_4633_nl;
  wire[0:0] mux_1512_nl;
  wire[0:0] mux_1516_nl;
  wire[0:0] or_4632_nl;
  wire[0:0] mux_1515_nl;
  wire[0:0] mux_1519_nl;
  wire[0:0] or_4631_nl;
  wire[0:0] mux_1518_nl;
  wire[0:0] mux_1522_nl;
  wire[0:0] or_4630_nl;
  wire[0:0] mux_1521_nl;
  wire[0:0] mux_1525_nl;
  wire[0:0] or_4629_nl;
  wire[0:0] mux_1524_nl;
  wire[0:0] mux_1527_nl;
  wire[0:0] or_3178_nl;
  wire[0:0] mux_1529_nl;
  wire[0:0] or_3183_nl;
  wire[0:0] mux_1531_nl;
  wire[0:0] or_3188_nl;
  wire[0:0] mux_1533_nl;
  wire[0:0] or_3193_nl;
  wire[0:0] mux_1535_nl;
  wire[0:0] or_3198_nl;
  wire[0:0] mux_1537_nl;
  wire[0:0] or_3203_nl;
  wire[0:0] mux_1539_nl;
  wire[0:0] or_3208_nl;
  wire[0:0] mux_1541_nl;
  wire[0:0] or_3213_nl;
  wire[0:0] mux_1544_nl;
  wire[0:0] or_4628_nl;
  wire[0:0] mux_1543_nl;
  wire[0:0] mux_1547_nl;
  wire[0:0] or_4627_nl;
  wire[0:0] mux_1546_nl;
  wire[0:0] mux_1445_nl;
  wire[0:0] mux_1440_nl;
  wire[0:0] mux_1430_nl;
  wire[0:0] mux_1439_nl;
  wire[0:0] mux_1438_nl;
  wire[0:0] and_385_nl;
  wire[0:0] mux_1444_nl;
  wire[0:0] mux_1441_nl;
  wire[0:0] or_2963_nl;
  wire[0:0] and_2500_nl;
  wire[0:0] mux_1548_nl;
  wire[0:0] and_2099_nl;
  wire[0:0] nor_750_nl;
  wire[0:0] mux_1549_nl;
  wire[0:0] and_2096_nl;
  wire[0:0] nor_747_nl;
  wire[0:0] mux_1550_nl;
  wire[0:0] and_2093_nl;
  wire[0:0] nor_744_nl;
  wire[0:0] mux_1551_nl;
  wire[0:0] and_2090_nl;
  wire[0:0] nor_741_nl;
  wire[0:0] mux_1552_nl;
  wire[0:0] and_2087_nl;
  wire[0:0] nor_738_nl;
  wire[0:0] mux_1553_nl;
  wire[0:0] and_2084_nl;
  wire[0:0] nor_735_nl;
  wire[0:0] mux_1554_nl;
  wire[0:0] and_2081_nl;
  wire[0:0] nor_732_nl;
  wire[0:0] mux_1555_nl;
  wire[0:0] and_2078_nl;
  wire[0:0] nor_729_nl;
  wire[0:0] mux_1556_nl;
  wire[0:0] and_2075_nl;
  wire[0:0] nor_726_nl;
  wire[0:0] mux_1557_nl;
  wire[0:0] and_2072_nl;
  wire[0:0] nor_723_nl;
  wire[0:0] mux_1558_nl;
  wire[0:0] and_2069_nl;
  wire[0:0] nor_720_nl;
  wire[0:0] mux_1559_nl;
  wire[0:0] and_2066_nl;
  wire[0:0] nor_717_nl;
  wire[0:0] mux_1560_nl;
  wire[0:0] and_2063_nl;
  wire[0:0] nor_714_nl;
  wire[0:0] mux_1561_nl;
  wire[0:0] and_2060_nl;
  wire[0:0] nor_711_nl;
  wire[0:0] mux_1562_nl;
  wire[0:0] and_2057_nl;
  wire[0:0] nor_708_nl;
  wire[0:0] mux_1563_nl;
  wire[0:0] and_2054_nl;
  wire[0:0] nor_705_nl;
  wire[0:0] mux_1565_nl;
  wire[0:0] mux_1564_nl;
  wire[0:0] and_2052_nl;
  wire[0:0] and_2053_nl;
  wire[0:0] nor_702_nl;
  wire[0:0] mux_1567_nl;
  wire[0:0] mux_1566_nl;
  wire[0:0] and_2050_nl;
  wire[0:0] and_2051_nl;
  wire[0:0] nor_701_nl;
  wire[0:0] mux_1569_nl;
  wire[0:0] mux_1568_nl;
  wire[0:0] and_2048_nl;
  wire[0:0] and_2049_nl;
  wire[0:0] nor_700_nl;
  wire[0:0] mux_1571_nl;
  wire[0:0] mux_1570_nl;
  wire[0:0] and_2046_nl;
  wire[0:0] and_2047_nl;
  wire[0:0] nor_699_nl;
  wire[0:0] mux_1573_nl;
  wire[0:0] mux_1572_nl;
  wire[0:0] and_2044_nl;
  wire[0:0] and_2045_nl;
  wire[0:0] nor_698_nl;
  wire[0:0] mux_1575_nl;
  wire[0:0] mux_1574_nl;
  wire[0:0] and_2042_nl;
  wire[0:0] and_2043_nl;
  wire[0:0] nor_697_nl;
  wire[0:0] mux_1577_nl;
  wire[0:0] mux_1576_nl;
  wire[0:0] and_2040_nl;
  wire[0:0] and_2041_nl;
  wire[0:0] nor_696_nl;
  wire[0:0] mux_1579_nl;
  wire[0:0] mux_1578_nl;
  wire[0:0] and_2038_nl;
  wire[0:0] and_2039_nl;
  wire[0:0] nor_695_nl;
  wire[0:0] mux_1581_nl;
  wire[0:0] mux_1580_nl;
  wire[0:0] and_2036_nl;
  wire[0:0] and_2037_nl;
  wire[0:0] nor_694_nl;
  wire[0:0] mux_1583_nl;
  wire[0:0] mux_1582_nl;
  wire[0:0] and_2034_nl;
  wire[0:0] and_2035_nl;
  wire[0:0] nor_693_nl;
  wire[0:0] mux_1585_nl;
  wire[0:0] mux_1584_nl;
  wire[0:0] and_2032_nl;
  wire[0:0] and_2033_nl;
  wire[0:0] nor_692_nl;
  wire[0:0] mux_1587_nl;
  wire[0:0] mux_1586_nl;
  wire[0:0] and_2030_nl;
  wire[0:0] and_2031_nl;
  wire[0:0] nor_691_nl;
  wire[0:0] mux_1589_nl;
  wire[0:0] mux_1588_nl;
  wire[0:0] and_2028_nl;
  wire[0:0] and_2029_nl;
  wire[0:0] nor_690_nl;
  wire[0:0] mux_1591_nl;
  wire[0:0] mux_1590_nl;
  wire[0:0] and_2026_nl;
  wire[0:0] and_2027_nl;
  wire[0:0] nor_689_nl;
  wire[0:0] mux_1593_nl;
  wire[0:0] mux_1592_nl;
  wire[0:0] and_2024_nl;
  wire[0:0] and_2025_nl;
  wire[0:0] nor_688_nl;
  wire[0:0] mux_1595_nl;
  wire[0:0] mux_1594_nl;
  wire[0:0] and_2022_nl;
  wire[0:0] and_2023_nl;
  wire[0:0] nor_687_nl;
  wire[0:0] mux_1596_nl;
  wire[0:0] nor_684_nl;
  wire[0:0] nor_686_nl;
  wire[0:0] mux_1597_nl;
  wire[0:0] nor_681_nl;
  wire[0:0] nor_683_nl;
  wire[0:0] mux_1598_nl;
  wire[0:0] nor_678_nl;
  wire[0:0] nor_680_nl;
  wire[0:0] mux_1599_nl;
  wire[0:0] nor_675_nl;
  wire[0:0] nor_677_nl;
  wire[0:0] mux_1600_nl;
  wire[0:0] nor_672_nl;
  wire[0:0] nor_674_nl;
  wire[0:0] mux_1601_nl;
  wire[0:0] nor_669_nl;
  wire[0:0] nor_671_nl;
  wire[0:0] mux_1602_nl;
  wire[0:0] nor_666_nl;
  wire[0:0] nor_668_nl;
  wire[0:0] mux_1603_nl;
  wire[0:0] nor_663_nl;
  wire[0:0] nor_665_nl;
  wire[0:0] mux_1604_nl;
  wire[0:0] nor_660_nl;
  wire[0:0] nor_662_nl;
  wire[0:0] mux_1605_nl;
  wire[0:0] nor_657_nl;
  wire[0:0] nor_659_nl;
  wire[0:0] mux_1606_nl;
  wire[0:0] nor_654_nl;
  wire[0:0] nor_656_nl;
  wire[0:0] mux_1607_nl;
  wire[0:0] nor_651_nl;
  wire[0:0] nor_653_nl;
  wire[0:0] mux_1608_nl;
  wire[0:0] nor_648_nl;
  wire[0:0] nor_650_nl;
  wire[0:0] mux_1609_nl;
  wire[0:0] nor_645_nl;
  wire[0:0] nor_647_nl;
  wire[0:0] mux_1610_nl;
  wire[0:0] nor_642_nl;
  wire[0:0] nor_644_nl;
  wire[0:0] mux_1611_nl;
  wire[0:0] nor_639_nl;
  wire[0:0] nor_641_nl;
  wire[0:0] and_552_nl;
  wire[0:0] and_554_nl;
  wire[0:0] and_556_nl;
  wire[0:0] and_558_nl;
  wire[0:0] and_560_nl;
  wire[0:0] and_562_nl;
  wire[0:0] and_564_nl;
  wire[0:0] and_566_nl;
  wire[0:0] and_568_nl;
  wire[0:0] and_570_nl;
  wire[0:0] and_572_nl;
  wire[0:0] and_574_nl;
  wire[0:0] and_576_nl;
  wire[0:0] and_578_nl;
  wire[0:0] and_580_nl;
  wire[0:0] and_582_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_178_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_65_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_144_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_2_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_182_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_67_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_146_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_6_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_1_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_186_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_69_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_148_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_10_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_2_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_190_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_71_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_150_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_14_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_3_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_194_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_73_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_152_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_18_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_4_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_198_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_75_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_154_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_22_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_5_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_202_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_77_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_156_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_26_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_6_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_206_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_79_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_158_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_30_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_7_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_210_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_81_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_160_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_34_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_8_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_214_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_83_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_162_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_38_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_9_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_218_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_85_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_164_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_42_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_10_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_222_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_87_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_166_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_46_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_11_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_226_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_89_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_168_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_50_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_12_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_230_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_91_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_170_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_54_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_13_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_234_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_93_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_172_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_58_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_14_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_238_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_95_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_174_nl;
  wire[1:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_62_nl;
  wire[3:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_15_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_2_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_2_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_3_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_3_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_4_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_4_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_5_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_5_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_6_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_6_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_7_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_7_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_8_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_8_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_9_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_9_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_10_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_10_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_11_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_11_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_12_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_12_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_13_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_13_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_14_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_14_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_15_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_15_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_16_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_16_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_177_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_239_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_181_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_145_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_1_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_66_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_1_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_185_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_147_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_68_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_2_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_189_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_149_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_3_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_70_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_3_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_193_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_151_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_72_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_4_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_197_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_153_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_5_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_74_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_5_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_201_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_155_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_76_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_6_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_205_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_157_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_7_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_78_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_7_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_209_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_159_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_80_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_8_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_213_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_161_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_9_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_82_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_9_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_217_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_163_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_84_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_10_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_221_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_165_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_11_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_86_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_11_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_225_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_167_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_88_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_12_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_229_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_169_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_13_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_90_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_13_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_233_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_171_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_92_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_14_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_237_nl;
  wire[9:0] FpExpoWidthInc_5U_8U_23U_1U_1U_mux_173_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_nor_15_nl;
  wire[2:0] FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_94_nl;
  wire[0:0] FpExpoWidthInc_5U_8U_23U_1U_1U_not_15_nl;
  wire[0:0] mul_loop_mul_16_FpMul_8U_23U_xor_nl;
  wire[0:0] mul_loop_mul_15_FpMul_8U_23U_xor_nl;
  wire[0:0] mul_loop_mul_14_FpMul_8U_23U_xor_nl;
  wire[0:0] mul_loop_mul_13_FpMul_8U_23U_xor_nl;
  wire[0:0] mul_loop_mul_12_FpMul_8U_23U_xor_nl;
  wire[0:0] mul_loop_mul_11_FpMul_8U_23U_xor_nl;
  wire[0:0] mul_loop_mul_10_FpMul_8U_23U_xor_nl;
  wire[0:0] mul_loop_mul_9_FpMul_8U_23U_xor_nl;
  wire[0:0] mul_loop_mul_8_FpMul_8U_23U_xor_nl;
  wire[0:0] mul_loop_mul_7_FpMul_8U_23U_xor_nl;
  wire[0:0] mul_loop_mul_6_FpMul_8U_23U_xor_nl;
  wire[0:0] mul_loop_mul_5_FpMul_8U_23U_xor_nl;
  wire[0:0] mul_loop_mul_4_FpMul_8U_23U_xor_nl;
  wire[0:0] mul_loop_mul_3_FpMul_8U_23U_xor_nl;
  wire[0:0] mul_loop_mul_2_FpMul_8U_23U_xor_nl;
  wire[0:0] mul_loop_mul_1_FpMul_8U_23U_xor_nl;
  wire[0:0] FpMul_8U_23U_p_mant_p1_and_31_nl;
  wire[8:0] mul_loop_mul_1_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_mul_loop_mul_1_FpMul_8U_23U_else_2_if_acc_nl;
  wire[8:0] mul_loop_mul_1_FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_mul_loop_mul_1_FpMul_8U_23U_else_2_acc_1_nl;
  wire[0:0] FpMul_8U_23U_p_mant_p1_and_30_nl;
  wire[8:0] mul_loop_mul_2_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_mul_loop_mul_2_FpMul_8U_23U_else_2_if_acc_nl;
  wire[8:0] mul_loop_mul_2_FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_mul_loop_mul_2_FpMul_8U_23U_else_2_acc_1_nl;
  wire[0:0] FpMul_8U_23U_p_mant_p1_and_29_nl;
  wire[8:0] mul_loop_mul_3_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_mul_loop_mul_3_FpMul_8U_23U_else_2_if_acc_nl;
  wire[8:0] mul_loop_mul_3_FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_mul_loop_mul_3_FpMul_8U_23U_else_2_acc_1_nl;
  wire[0:0] FpMul_8U_23U_p_mant_p1_and_28_nl;
  wire[8:0] mul_loop_mul_4_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_mul_loop_mul_4_FpMul_8U_23U_else_2_if_acc_nl;
  wire[8:0] mul_loop_mul_4_FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_mul_loop_mul_4_FpMul_8U_23U_else_2_acc_1_nl;
  wire[0:0] FpMul_8U_23U_p_mant_p1_and_27_nl;
  wire[8:0] mul_loop_mul_5_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_mul_loop_mul_5_FpMul_8U_23U_else_2_if_acc_nl;
  wire[8:0] mul_loop_mul_5_FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_mul_loop_mul_5_FpMul_8U_23U_else_2_acc_1_nl;
  wire[0:0] FpMul_8U_23U_p_mant_p1_and_26_nl;
  wire[8:0] mul_loop_mul_6_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_mul_loop_mul_6_FpMul_8U_23U_else_2_if_acc_nl;
  wire[8:0] mul_loop_mul_6_FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_mul_loop_mul_6_FpMul_8U_23U_else_2_acc_1_nl;
  wire[0:0] FpMul_8U_23U_p_mant_p1_and_25_nl;
  wire[8:0] mul_loop_mul_7_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_mul_loop_mul_7_FpMul_8U_23U_else_2_if_acc_nl;
  wire[8:0] mul_loop_mul_7_FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_mul_loop_mul_7_FpMul_8U_23U_else_2_acc_1_nl;
  wire[0:0] FpMul_8U_23U_p_mant_p1_and_24_nl;
  wire[8:0] mul_loop_mul_8_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_mul_loop_mul_8_FpMul_8U_23U_else_2_if_acc_nl;
  wire[8:0] mul_loop_mul_8_FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_mul_loop_mul_8_FpMul_8U_23U_else_2_acc_1_nl;
  wire[0:0] FpMul_8U_23U_p_mant_p1_and_23_nl;
  wire[8:0] mul_loop_mul_9_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_mul_loop_mul_9_FpMul_8U_23U_else_2_if_acc_nl;
  wire[8:0] mul_loop_mul_9_FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_mul_loop_mul_9_FpMul_8U_23U_else_2_acc_1_nl;
  wire[0:0] FpMul_8U_23U_p_mant_p1_and_22_nl;
  wire[8:0] mul_loop_mul_10_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_mul_loop_mul_10_FpMul_8U_23U_else_2_if_acc_nl;
  wire[8:0] mul_loop_mul_10_FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_mul_loop_mul_10_FpMul_8U_23U_else_2_acc_1_nl;
  wire[0:0] FpMul_8U_23U_p_mant_p1_and_21_nl;
  wire[8:0] mul_loop_mul_11_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_mul_loop_mul_11_FpMul_8U_23U_else_2_if_acc_nl;
  wire[8:0] mul_loop_mul_11_FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_mul_loop_mul_11_FpMul_8U_23U_else_2_acc_1_nl;
  wire[0:0] FpMul_8U_23U_p_mant_p1_and_20_nl;
  wire[8:0] mul_loop_mul_12_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_mul_loop_mul_12_FpMul_8U_23U_else_2_if_acc_nl;
  wire[8:0] mul_loop_mul_12_FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_mul_loop_mul_12_FpMul_8U_23U_else_2_acc_1_nl;
  wire[0:0] FpMul_8U_23U_p_mant_p1_and_19_nl;
  wire[8:0] mul_loop_mul_13_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_mul_loop_mul_13_FpMul_8U_23U_else_2_if_acc_nl;
  wire[8:0] mul_loop_mul_13_FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_mul_loop_mul_13_FpMul_8U_23U_else_2_acc_1_nl;
  wire[0:0] FpMul_8U_23U_p_mant_p1_and_18_nl;
  wire[8:0] mul_loop_mul_14_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_mul_loop_mul_14_FpMul_8U_23U_else_2_if_acc_nl;
  wire[8:0] mul_loop_mul_14_FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_mul_loop_mul_14_FpMul_8U_23U_else_2_acc_1_nl;
  wire[0:0] FpMul_8U_23U_p_mant_p1_and_17_nl;
  wire[8:0] mul_loop_mul_15_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_mul_loop_mul_15_FpMul_8U_23U_else_2_if_acc_nl;
  wire[8:0] mul_loop_mul_15_FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_mul_loop_mul_15_FpMul_8U_23U_else_2_acc_1_nl;
  wire[0:0] FpMul_8U_23U_p_mant_p1_and_16_nl;
  wire[8:0] mul_loop_mul_16_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_mul_loop_mul_16_FpMul_8U_23U_else_2_if_acc_nl;
  wire[8:0] mul_loop_mul_16_FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_mul_loop_mul_16_FpMul_8U_23U_else_2_acc_1_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_110_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_48_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_108_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_50_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_106_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_52_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_104_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_54_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_102_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_56_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_100_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_58_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_98_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_60_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_96_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_62_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_94_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_64_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_92_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_66_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_90_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_68_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_88_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_70_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_86_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_72_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_84_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_74_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_82_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_76_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_80_nl;
  wire[0:0] mul_nan_to_zero_aelse_not_78_nl;
  wire[9:0] mul_loop_mul_1_FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_mul_loop_mul_1_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_nl;
  wire[9:0] mul_loop_mul_2_FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_mul_loop_mul_2_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_1_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_1_nl;
  wire[9:0] mul_loop_mul_3_FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_mul_loop_mul_3_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_2_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_2_nl;
  wire[9:0] mul_loop_mul_4_FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_mul_loop_mul_4_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_3_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_3_nl;
  wire[9:0] mul_loop_mul_5_FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_mul_loop_mul_5_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_4_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_4_nl;
  wire[9:0] mul_loop_mul_6_FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_mul_loop_mul_6_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_5_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_5_nl;
  wire[9:0] mul_loop_mul_7_FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_mul_loop_mul_7_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_6_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_6_nl;
  wire[9:0] mul_loop_mul_8_FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_mul_loop_mul_8_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_7_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_7_nl;
  wire[9:0] mul_loop_mul_9_FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_mul_loop_mul_9_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_8_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_8_nl;
  wire[9:0] mul_loop_mul_10_FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_mul_loop_mul_10_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_9_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_9_nl;
  wire[9:0] mul_loop_mul_11_FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_mul_loop_mul_11_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_10_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_10_nl;
  wire[9:0] mul_loop_mul_12_FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_mul_loop_mul_12_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_11_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_11_nl;
  wire[9:0] mul_loop_mul_13_FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_mul_loop_mul_13_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_12_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_12_nl;
  wire[9:0] mul_loop_mul_14_FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_mul_loop_mul_14_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_13_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_13_nl;
  wire[9:0] mul_loop_mul_15_FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_mul_loop_mul_15_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_14_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_14_nl;
  wire[9:0] mul_loop_mul_16_FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_mul_loop_mul_16_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_15_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_15_nl;
  wire[7:0] mul_loop_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_mul_loop_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_63_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_1_nl;
  wire[7:0] mul_loop_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_mul_loop_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_62_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_2_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_3_nl;
  wire[7:0] mul_loop_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_mul_loop_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_61_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_4_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_5_nl;
  wire[7:0] mul_loop_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_mul_loop_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_60_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_6_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_7_nl;
  wire[7:0] mul_loop_mul_5_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_mul_loop_mul_5_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_59_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_8_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_9_nl;
  wire[7:0] mul_loop_mul_6_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_mul_loop_mul_6_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_58_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_10_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_11_nl;
  wire[7:0] mul_loop_mul_7_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_mul_loop_mul_7_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_57_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_12_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_13_nl;
  wire[7:0] mul_loop_mul_8_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_mul_loop_mul_8_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_56_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_14_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_15_nl;
  wire[7:0] mul_loop_mul_9_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_mul_loop_mul_9_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_55_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_16_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_17_nl;
  wire[7:0] mul_loop_mul_10_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_mul_loop_mul_10_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_54_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_18_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_19_nl;
  wire[7:0] mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_53_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_20_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_21_nl;
  wire[7:0] mul_loop_mul_12_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_mul_loop_mul_12_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_52_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_22_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_23_nl;
  wire[7:0] mul_loop_mul_13_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_mul_loop_mul_13_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_51_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_24_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_25_nl;
  wire[7:0] mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_50_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_26_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_27_nl;
  wire[7:0] mul_loop_mul_15_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_mul_loop_mul_15_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_49_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_28_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_29_nl;
  wire[7:0] mul_loop_mul_16_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_mul_loop_mul_16_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_48_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_30_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_31_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_32_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_33_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_34_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_35_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_36_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_37_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_38_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_39_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_40_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_41_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_42_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_43_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_44_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_45_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_46_nl;
  wire[0:0] IsNaN_5U_23U_aelse_not_47_nl;
  wire[7:0] mul_loop_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_mul_loop_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[0:0] mux_1664_nl;
  wire[7:0] mul_loop_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_mul_loop_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[0:0] mux_1665_nl;
  wire[7:0] mul_loop_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_mul_loop_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[0:0] mux_1666_nl;
  wire[7:0] mul_loop_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_mul_loop_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[0:0] mux_1667_nl;
  wire[7:0] mul_loop_mul_5_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_mul_loop_mul_5_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[0:0] mux_1668_nl;
  wire[7:0] mul_loop_mul_6_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_mul_loop_mul_6_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[0:0] mux_1669_nl;
  wire[7:0] mul_loop_mul_7_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_mul_loop_mul_7_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[0:0] mux_1670_nl;
  wire[7:0] mul_loop_mul_8_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_mul_loop_mul_8_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[0:0] mux_1671_nl;
  wire[7:0] mul_loop_mul_9_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_mul_loop_mul_9_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[0:0] mux_1672_nl;
  wire[7:0] mul_loop_mul_10_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_mul_loop_mul_10_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[0:0] mux_1673_nl;
  wire[7:0] mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[0:0] mux_1674_nl;
  wire[0:0] nor_606_nl;
  wire[0:0] nand_170_nl;
  wire[7:0] mul_loop_mul_12_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_mul_loop_mul_12_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[0:0] mux_1675_nl;
  wire[7:0] mul_loop_mul_13_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_mul_loop_mul_13_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[0:0] mux_1676_nl;
  wire[7:0] mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[0:0] mux_1677_nl;
  wire[7:0] mul_loop_mul_15_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_mul_loop_mul_15_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[0:0] mux_1678_nl;
  wire[7:0] mul_loop_mul_16_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_mul_loop_mul_16_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[0:0] mux_1679_nl;
  wire[0:0] mux_7_nl;
  wire[0:0] or_4664_nl;
  wire[0:0] mux_11_nl;
  wire[0:0] mux_14_nl;
  wire[0:0] mux_10_nl;
  wire[0:0] mux_13_nl;
  wire[0:0] mux_20_nl;
  wire[0:0] or_4662_nl;
  wire[0:0] mux_24_nl;
  wire[0:0] mux_22_nl;
  wire[0:0] mux_23_nl;
  wire[0:0] mux_30_nl;
  wire[0:0] or_4661_nl;
  wire[0:0] mux_34_nl;
  wire[0:0] mux_32_nl;
  wire[0:0] mux_33_nl;
  wire[0:0] or_117_nl;
  wire[0:0] mux_44_nl;
  wire[0:0] mux_50_nl;
  wire[0:0] or_4660_nl;
  wire[0:0] mux_54_nl;
  wire[0:0] mux_52_nl;
  wire[0:0] mux_53_nl;
  wire[0:0] or_132_nl;
  wire[0:0] mux_61_nl;
  wire[0:0] or_138_nl;
  wire[0:0] mux_68_nl;
  wire[0:0] mux_74_nl;
  wire[0:0] or_4659_nl;
  wire[0:0] mux_78_nl;
  wire[0:0] mux_76_nl;
  wire[0:0] mux_77_nl;
  wire[0:0] mux_84_nl;
  wire[0:0] or_4658_nl;
  wire[0:0] mux_88_nl;
  wire[0:0] mux_86_nl;
  wire[0:0] mux_87_nl;
  wire[0:0] or_158_nl;
  wire[0:0] mux_95_nl;
  wire[0:0] or_164_nl;
  wire[0:0] mux_102_nl;
  wire[0:0] or_170_nl;
  wire[0:0] mux_109_nl;
  wire[0:0] mux_115_nl;
  wire[0:0] or_4657_nl;
  wire[0:0] mux_119_nl;
  wire[0:0] mux_117_nl;
  wire[0:0] mux_118_nl;
  wire[0:0] or_183_nl;
  wire[0:0] mux_126_nl;
  wire[0:0] mux_132_nl;
  wire[0:0] or_4656_nl;
  wire[0:0] mux_136_nl;
  wire[0:0] mux_134_nl;
  wire[0:0] mux_135_nl;
  wire[0:0] mux_142_nl;
  wire[0:0] or_4655_nl;
  wire[0:0] mux_146_nl;
  wire[0:0] mux_144_nl;
  wire[0:0] mux_145_nl;
  wire[0:0] and_2250_nl;
  wire[0:0] or_210_nl;
  wire[0:0] or_216_nl;
  wire[0:0] or_222_nl;
  wire[0:0] or_229_nl;
  wire[0:0] or_235_nl;
  wire[0:0] or_239_nl;
  wire[0:0] or_243_nl;
  wire[0:0] or_249_nl;
  wire[0:0] or_255_nl;
  wire[0:0] or_259_nl;
  wire[0:0] or_263_nl;
  wire[0:0] or_267_nl;
  wire[0:0] or_273_nl;
  wire[0:0] or_277_nl;
  wire[0:0] or_283_nl;
  wire[0:0] or_289_nl;
  wire[0:0] or_1044_nl;
  wire[0:0] or_1049_nl;
  wire[0:0] or_1124_nl;
  wire[0:0] or_1129_nl;
  wire[0:0] or_1206_nl;
  wire[0:0] or_1211_nl;
  wire[0:0] or_1289_nl;
  wire[0:0] or_1294_nl;
  wire[0:0] or_1369_nl;
  wire[0:0] or_1374_nl;
  wire[0:0] or_1451_nl;
  wire[0:0] or_1456_nl;
  wire[0:0] or_1533_nl;
  wire[0:0] or_1538_nl;
  wire[0:0] or_1613_nl;
  wire[0:0] or_1618_nl;
  wire[0:0] or_1693_nl;
  wire[0:0] or_1698_nl;
  wire[0:0] or_1773_nl;
  wire[0:0] or_1778_nl;
  wire[0:0] or_1828_nl;
  wire[0:0] or_1856_nl;
  wire[0:0] or_1934_nl;
  wire[0:0] or_1939_nl;
  wire[0:0] or_2017_nl;
  wire[0:0] or_2022_nl;
  wire[0:0] or_2101_nl;
  wire[0:0] or_2106_nl;
  wire[0:0] or_2183_nl;
  wire[0:0] or_2188_nl;
  wire[0:0] or_2263_nl;
  wire[0:0] or_2268_nl;
  wire[0:0] mux_1138_nl;
  wire[0:0] or_2591_nl;
  wire[0:0] mux_1160_nl;
  wire[0:0] or_2622_nl;
  wire[0:0] mux_1183_nl;
  wire[0:0] or_2645_nl;
  wire[0:0] mux_1210_nl;
  wire[0:0] or_2689_nl;
  wire[0:0] mux_1244_nl;
  wire[0:0] or_2736_nl;
  wire[0:0] mux_1267_nl;
  wire[0:0] or_2759_nl;
  wire[0:0] mux_1306_nl;
  wire[0:0] or_2812_nl;
  wire[0:0] mux_1334_nl;
  wire[0:0] or_2848_nl;
  wire[0:0] mux_1356_nl;
  wire[0:0] or_2879_nl;
  wire[0:0] or_2950_nl;
  wire[0:0] mux_1428_nl;
  wire[0:0] or_2958_nl;
  wire[0:0] mux_1431_nl;
  wire[0:0] or_2961_nl;
  wire[0:0] mux_1632_nl;
  wire[0:0] and_1042_nl;
  wire[0:0] mux_1633_nl;
  wire[0:0] and_1046_nl;
  wire[0:0] mux_1634_nl;
  wire[0:0] and_1050_nl;
  wire[0:0] mux_1635_nl;
  wire[0:0] and_1054_nl;
  wire[0:0] mux_1636_nl;
  wire[0:0] and_1058_nl;
  wire[0:0] mux_1637_nl;
  wire[0:0] and_1062_nl;
  wire[0:0] mux_1638_nl;
  wire[0:0] and_1066_nl;
  wire[0:0] mux_1639_nl;
  wire[0:0] and_1070_nl;
  wire[0:0] mux_1640_nl;
  wire[0:0] and_1074_nl;
  wire[0:0] mux_1641_nl;
  wire[0:0] and_1078_nl;
  wire[0:0] mux_1642_nl;
  wire[0:0] and_1082_nl;
  wire[0:0] mux_1643_nl;
  wire[0:0] and_1086_nl;
  wire[0:0] mux_1644_nl;
  wire[0:0] and_1090_nl;
  wire[0:0] mux_1645_nl;
  wire[0:0] and_1094_nl;
  wire[0:0] mux_1646_nl;
  wire[0:0] and_1098_nl;
  wire[0:0] mux_1647_nl;
  wire[0:0] and_1102_nl;
// Interconnect Declarations for Component Instantiations
  wire [21:0] nl_mul_loop_mul_1_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_mul_loop_mul_1_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a = {(mul_nan_to_zero_op_mant_1_lpi_1_dfm[8:0])
      , 13'b0};
  wire [6:0] nl_mul_loop_mul_1_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_mul_loop_mul_1_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_16)
      + 6'b1;
  wire [22:0] nl_mul_loop_mul_1_leading_sign_23_0_rg_mantissa;
  assign nl_mul_loop_mul_1_leading_sign_23_0_rg_mantissa = {mul_nan_to_zero_op_mant_1_lpi_1_dfm
      , 13'b0};
  wire [21:0] nl_mul_loop_mul_2_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_mul_loop_mul_2_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a = {(mul_nan_to_zero_op_mant_2_lpi_1_dfm[8:0])
      , 13'b0};
  wire [6:0] nl_mul_loop_mul_2_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_mul_loop_mul_2_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_17)
      + 6'b1;
  wire [22:0] nl_mul_loop_mul_2_leading_sign_23_0_rg_mantissa;
  assign nl_mul_loop_mul_2_leading_sign_23_0_rg_mantissa = {mul_nan_to_zero_op_mant_2_lpi_1_dfm
      , 13'b0};
  wire [21:0] nl_mul_loop_mul_3_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_mul_loop_mul_3_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a = {(mul_nan_to_zero_op_mant_3_lpi_1_dfm[8:0])
      , 13'b0};
  wire [6:0] nl_mul_loop_mul_3_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_mul_loop_mul_3_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_18)
      + 6'b1;
  wire [22:0] nl_mul_loop_mul_3_leading_sign_23_0_rg_mantissa;
  assign nl_mul_loop_mul_3_leading_sign_23_0_rg_mantissa = {mul_nan_to_zero_op_mant_3_lpi_1_dfm
      , 13'b0};
  wire [21:0] nl_mul_loop_mul_4_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_mul_loop_mul_4_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a = {(mul_nan_to_zero_op_mant_4_lpi_1_dfm[8:0])
      , 13'b0};
  wire [6:0] nl_mul_loop_mul_4_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_mul_loop_mul_4_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_19)
      + 6'b1;
  wire [22:0] nl_mul_loop_mul_4_leading_sign_23_0_rg_mantissa;
  assign nl_mul_loop_mul_4_leading_sign_23_0_rg_mantissa = {mul_nan_to_zero_op_mant_4_lpi_1_dfm
      , 13'b0};
  wire [21:0] nl_mul_loop_mul_5_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_mul_loop_mul_5_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a = {(mul_nan_to_zero_op_mant_5_lpi_1_dfm[8:0])
      , 13'b0};
  wire [6:0] nl_mul_loop_mul_5_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_mul_loop_mul_5_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_20)
      + 6'b1;
  wire [22:0] nl_mul_loop_mul_5_leading_sign_23_0_rg_mantissa;
  assign nl_mul_loop_mul_5_leading_sign_23_0_rg_mantissa = {mul_nan_to_zero_op_mant_5_lpi_1_dfm
      , 13'b0};
  wire [21:0] nl_mul_loop_mul_6_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_mul_loop_mul_6_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a = {(mul_nan_to_zero_op_mant_6_lpi_1_dfm[8:0])
      , 13'b0};
  wire [6:0] nl_mul_loop_mul_6_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_mul_loop_mul_6_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_21)
      + 6'b1;
  wire [22:0] nl_mul_loop_mul_6_leading_sign_23_0_rg_mantissa;
  assign nl_mul_loop_mul_6_leading_sign_23_0_rg_mantissa = {mul_nan_to_zero_op_mant_6_lpi_1_dfm
      , 13'b0};
  wire [21:0] nl_mul_loop_mul_7_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_mul_loop_mul_7_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a = {(mul_nan_to_zero_op_mant_7_lpi_1_dfm[8:0])
      , 13'b0};
  wire [6:0] nl_mul_loop_mul_7_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_mul_loop_mul_7_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_22)
      + 6'b1;
  wire [22:0] nl_mul_loop_mul_7_leading_sign_23_0_rg_mantissa;
  assign nl_mul_loop_mul_7_leading_sign_23_0_rg_mantissa = {mul_nan_to_zero_op_mant_7_lpi_1_dfm
      , 13'b0};
  wire [21:0] nl_mul_loop_mul_8_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_mul_loop_mul_8_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a = {(mul_nan_to_zero_op_mant_8_lpi_1_dfm[8:0])
      , 13'b0};
  wire [6:0] nl_mul_loop_mul_8_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_mul_loop_mul_8_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_23)
      + 6'b1;
  wire [22:0] nl_mul_loop_mul_8_leading_sign_23_0_rg_mantissa;
  assign nl_mul_loop_mul_8_leading_sign_23_0_rg_mantissa = {mul_nan_to_zero_op_mant_8_lpi_1_dfm
      , 13'b0};
  wire [21:0] nl_mul_loop_mul_9_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_mul_loop_mul_9_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a = {(mul_nan_to_zero_op_mant_9_lpi_1_dfm[8:0])
      , 13'b0};
  wire [6:0] nl_mul_loop_mul_9_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_mul_loop_mul_9_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_24)
      + 6'b1;
  wire [22:0] nl_mul_loop_mul_9_leading_sign_23_0_rg_mantissa;
  assign nl_mul_loop_mul_9_leading_sign_23_0_rg_mantissa = {mul_nan_to_zero_op_mant_9_lpi_1_dfm
      , 13'b0};
  wire [21:0] nl_mul_loop_mul_10_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_mul_loop_mul_10_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a =
      {(mul_nan_to_zero_op_mant_10_lpi_1_dfm[8:0]) , 13'b0};
  wire [6:0] nl_mul_loop_mul_10_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_mul_loop_mul_10_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s =
      conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_25)
      + 6'b1;
  wire [22:0] nl_mul_loop_mul_10_leading_sign_23_0_rg_mantissa;
  assign nl_mul_loop_mul_10_leading_sign_23_0_rg_mantissa = {mul_nan_to_zero_op_mant_10_lpi_1_dfm
      , 13'b0};
  wire [21:0] nl_mul_loop_mul_11_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_mul_loop_mul_11_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a =
      {(mul_nan_to_zero_op_mant_11_lpi_1_dfm[8:0]) , 13'b0};
  wire [6:0] nl_mul_loop_mul_11_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_mul_loop_mul_11_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s =
      conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_26)
      + 6'b1;
  wire [22:0] nl_mul_loop_mul_11_leading_sign_23_0_rg_mantissa;
  assign nl_mul_loop_mul_11_leading_sign_23_0_rg_mantissa = {mul_nan_to_zero_op_mant_11_lpi_1_dfm
      , 13'b0};
  wire [21:0] nl_mul_loop_mul_12_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_mul_loop_mul_12_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a =
      {(mul_nan_to_zero_op_mant_12_lpi_1_dfm[8:0]) , 13'b0};
  wire [6:0] nl_mul_loop_mul_12_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_mul_loop_mul_12_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s =
      conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_27)
      + 6'b1;
  wire [22:0] nl_mul_loop_mul_12_leading_sign_23_0_rg_mantissa;
  assign nl_mul_loop_mul_12_leading_sign_23_0_rg_mantissa = {mul_nan_to_zero_op_mant_12_lpi_1_dfm
      , 13'b0};
  wire [21:0] nl_mul_loop_mul_13_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_mul_loop_mul_13_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a =
      {(mul_nan_to_zero_op_mant_13_lpi_1_dfm[8:0]) , 13'b0};
  wire [6:0] nl_mul_loop_mul_13_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_mul_loop_mul_13_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s =
      conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_28)
      + 6'b1;
  wire [22:0] nl_mul_loop_mul_13_leading_sign_23_0_rg_mantissa;
  assign nl_mul_loop_mul_13_leading_sign_23_0_rg_mantissa = {mul_nan_to_zero_op_mant_13_lpi_1_dfm
      , 13'b0};
  wire [21:0] nl_mul_loop_mul_14_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_mul_loop_mul_14_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a =
      {(mul_nan_to_zero_op_mant_14_lpi_1_dfm[8:0]) , 13'b0};
  wire [6:0] nl_mul_loop_mul_14_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_mul_loop_mul_14_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s =
      conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_29)
      + 6'b1;
  wire [22:0] nl_mul_loop_mul_14_leading_sign_23_0_rg_mantissa;
  assign nl_mul_loop_mul_14_leading_sign_23_0_rg_mantissa = {mul_nan_to_zero_op_mant_14_lpi_1_dfm
      , 13'b0};
  wire [21:0] nl_mul_loop_mul_15_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_mul_loop_mul_15_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a =
      {(mul_nan_to_zero_op_mant_15_lpi_1_dfm[8:0]) , 13'b0};
  wire [6:0] nl_mul_loop_mul_15_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_mul_loop_mul_15_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s =
      conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_30)
      + 6'b1;
  wire [22:0] nl_mul_loop_mul_15_leading_sign_23_0_rg_mantissa;
  assign nl_mul_loop_mul_15_leading_sign_23_0_rg_mantissa = {mul_nan_to_zero_op_mant_15_lpi_1_dfm
      , 13'b0};
  wire [21:0] nl_mul_loop_mul_16_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_mul_loop_mul_16_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a =
      {(mul_nan_to_zero_op_mant_lpi_1_dfm[8:0]) , 13'b0};
  wire [6:0] nl_mul_loop_mul_16_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_mul_loop_mul_16_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s =
      conv_u2u_5_6(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_31)
      + 6'b1;
  wire [22:0] nl_mul_loop_mul_16_leading_sign_23_0_rg_mantissa;
  assign nl_mul_loop_mul_16_leading_sign_23_0_rg_mantissa = {mul_nan_to_zero_op_mant_lpi_1_dfm
      , 13'b0};
  wire [799:0] nl_X_mul_core_chn_mul_out_rsci_inst_chn_mul_out_rsci_d;
  assign nl_X_mul_core_chn_mul_out_rsci_inst_chn_mul_out_rsci_d = {chn_mul_out_rsci_d_799
      , chn_mul_out_rsci_d_798 , chn_mul_out_rsci_d_797 , chn_mul_out_rsci_d_796
      , chn_mul_out_rsci_d_795 , chn_mul_out_rsci_d_794 , chn_mul_out_rsci_d_793
      , chn_mul_out_rsci_d_792 , chn_mul_out_rsci_d_791 , chn_mul_out_rsci_d_790
      , chn_mul_out_rsci_d_789 , chn_mul_out_rsci_d_788 , chn_mul_out_rsci_d_787
      , chn_mul_out_rsci_d_786 , chn_mul_out_rsci_d_785 , chn_mul_out_rsci_d_784
      , chn_mul_out_rsci_d_783_766 , chn_mul_out_rsci_d_765_764 , chn_mul_out_rsci_d_763_762
      , chn_mul_out_rsci_d_761_758 , chn_mul_out_rsci_d_757_748 , chn_mul_out_rsci_d_747_745
      , chn_mul_out_rsci_d_744_735 , chn_mul_out_rsci_d_734_717 , chn_mul_out_rsci_d_716_715
      , chn_mul_out_rsci_d_714_713 , chn_mul_out_rsci_d_712_709 , chn_mul_out_rsci_d_708_699
      , chn_mul_out_rsci_d_698_696 , chn_mul_out_rsci_d_695_686 , chn_mul_out_rsci_d_685_668
      , chn_mul_out_rsci_d_667_666 , chn_mul_out_rsci_d_665_664 , chn_mul_out_rsci_d_663_660
      , chn_mul_out_rsci_d_659_650 , chn_mul_out_rsci_d_649_647 , chn_mul_out_rsci_d_646_637
      , chn_mul_out_rsci_d_636_619 , chn_mul_out_rsci_d_618_617 , chn_mul_out_rsci_d_616_615
      , chn_mul_out_rsci_d_614_611 , chn_mul_out_rsci_d_610_601 , chn_mul_out_rsci_d_600_598
      , chn_mul_out_rsci_d_597_588 , chn_mul_out_rsci_d_587_570 , chn_mul_out_rsci_d_569_568
      , chn_mul_out_rsci_d_567_566 , chn_mul_out_rsci_d_565_562 , chn_mul_out_rsci_d_561_552
      , chn_mul_out_rsci_d_551_549 , chn_mul_out_rsci_d_548_539 , chn_mul_out_rsci_d_538_521
      , chn_mul_out_rsci_d_520_519 , chn_mul_out_rsci_d_518_517 , chn_mul_out_rsci_d_516_513
      , chn_mul_out_rsci_d_512_503 , chn_mul_out_rsci_d_502_500 , chn_mul_out_rsci_d_499_490
      , chn_mul_out_rsci_d_489_472 , chn_mul_out_rsci_d_471_470 , chn_mul_out_rsci_d_469_468
      , chn_mul_out_rsci_d_467_464 , chn_mul_out_rsci_d_463_454 , chn_mul_out_rsci_d_453_451
      , chn_mul_out_rsci_d_450_441 , chn_mul_out_rsci_d_440_423 , chn_mul_out_rsci_d_422_421
      , chn_mul_out_rsci_d_420_419 , chn_mul_out_rsci_d_418_415 , chn_mul_out_rsci_d_414_405
      , chn_mul_out_rsci_d_404_402 , chn_mul_out_rsci_d_401_392 , chn_mul_out_rsci_d_391_374
      , chn_mul_out_rsci_d_373_372 , chn_mul_out_rsci_d_371_370 , chn_mul_out_rsci_d_369_366
      , chn_mul_out_rsci_d_365_356 , chn_mul_out_rsci_d_355_353 , chn_mul_out_rsci_d_352_343
      , chn_mul_out_rsci_d_342_325 , chn_mul_out_rsci_d_324_323 , chn_mul_out_rsci_d_322_321
      , chn_mul_out_rsci_d_320_317 , chn_mul_out_rsci_d_316_307 , chn_mul_out_rsci_d_306_304
      , chn_mul_out_rsci_d_303_294 , chn_mul_out_rsci_d_293_276 , chn_mul_out_rsci_d_275_274
      , chn_mul_out_rsci_d_273_272 , chn_mul_out_rsci_d_271_268 , chn_mul_out_rsci_d_267_258
      , chn_mul_out_rsci_d_257_255 , chn_mul_out_rsci_d_254_245 , chn_mul_out_rsci_d_244_227
      , chn_mul_out_rsci_d_226_225 , chn_mul_out_rsci_d_224_223 , chn_mul_out_rsci_d_222_219
      , chn_mul_out_rsci_d_218_209 , chn_mul_out_rsci_d_208_206 , chn_mul_out_rsci_d_205_196
      , chn_mul_out_rsci_d_195_178 , chn_mul_out_rsci_d_177_176 , chn_mul_out_rsci_d_175_174
      , chn_mul_out_rsci_d_173_170 , chn_mul_out_rsci_d_169_160 , chn_mul_out_rsci_d_159_157
      , chn_mul_out_rsci_d_156_147 , chn_mul_out_rsci_d_146_129 , chn_mul_out_rsci_d_128_127
      , chn_mul_out_rsci_d_126_125 , chn_mul_out_rsci_d_124_121 , chn_mul_out_rsci_d_120_111
      , chn_mul_out_rsci_d_110_108 , chn_mul_out_rsci_d_107_98 , chn_mul_out_rsci_d_97_80
      , chn_mul_out_rsci_d_79_78 , chn_mul_out_rsci_d_77_76 , chn_mul_out_rsci_d_75_72
      , chn_mul_out_rsci_d_71_62 , chn_mul_out_rsci_d_61_59 , chn_mul_out_rsci_d_58_49
      , chn_mul_out_rsci_d_48_31 , chn_mul_out_rsci_d_30_29 , chn_mul_out_rsci_d_28_27
      , chn_mul_out_rsci_d_26_23 , chn_mul_out_rsci_d_22_13 , chn_mul_out_rsci_d_12_10
      , chn_mul_out_rsci_d_9_0};
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) mul_loop_mul_1_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_mul_loop_mul_1_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_mul_loop_mul_1_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_sva_2)
    );
  SDP_X_leading_sign_23_0 mul_loop_mul_1_leading_sign_23_0_rg (
      .mantissa(nl_mul_loop_mul_1_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_16)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) mul_loop_mul_2_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_mul_loop_mul_2_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_mul_loop_mul_2_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_sva_2)
    );
  SDP_X_leading_sign_23_0 mul_loop_mul_2_leading_sign_23_0_rg (
      .mantissa(nl_mul_loop_mul_2_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_17)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) mul_loop_mul_3_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_mul_loop_mul_3_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_mul_loop_mul_3_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_sva_2)
    );
  SDP_X_leading_sign_23_0 mul_loop_mul_3_leading_sign_23_0_rg (
      .mantissa(nl_mul_loop_mul_3_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_18)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) mul_loop_mul_4_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_mul_loop_mul_4_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_mul_loop_mul_4_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_sva_2)
    );
  SDP_X_leading_sign_23_0 mul_loop_mul_4_leading_sign_23_0_rg (
      .mantissa(nl_mul_loop_mul_4_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_19)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) mul_loop_mul_5_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_mul_loop_mul_5_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_mul_loop_mul_5_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_sva_2)
    );
  SDP_X_leading_sign_23_0 mul_loop_mul_5_leading_sign_23_0_rg (
      .mantissa(nl_mul_loop_mul_5_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_20)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) mul_loop_mul_6_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_mul_loop_mul_6_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_mul_loop_mul_6_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_sva_2)
    );
  SDP_X_leading_sign_23_0 mul_loop_mul_6_leading_sign_23_0_rg (
      .mantissa(nl_mul_loop_mul_6_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_21)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) mul_loop_mul_7_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_mul_loop_mul_7_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_mul_loop_mul_7_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_sva_2)
    );
  SDP_X_leading_sign_23_0 mul_loop_mul_7_leading_sign_23_0_rg (
      .mantissa(nl_mul_loop_mul_7_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_22)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) mul_loop_mul_8_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_mul_loop_mul_8_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_mul_loop_mul_8_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_sva_2)
    );
  SDP_X_leading_sign_23_0 mul_loop_mul_8_leading_sign_23_0_rg (
      .mantissa(nl_mul_loop_mul_8_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_23)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) mul_loop_mul_9_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_mul_loop_mul_9_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_mul_loop_mul_9_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_sva_2)
    );
  SDP_X_leading_sign_23_0 mul_loop_mul_9_leading_sign_23_0_rg (
      .mantissa(nl_mul_loop_mul_9_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_24)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) mul_loop_mul_10_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_mul_loop_mul_10_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_mul_loop_mul_10_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_sva_2)
    );
  SDP_X_leading_sign_23_0 mul_loop_mul_10_leading_sign_23_0_rg (
      .mantissa(nl_mul_loop_mul_10_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_25)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) mul_loop_mul_11_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_mul_loop_mul_11_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_mul_loop_mul_11_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_sva_2)
    );
  SDP_X_leading_sign_23_0 mul_loop_mul_11_leading_sign_23_0_rg (
      .mantissa(nl_mul_loop_mul_11_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_26)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) mul_loop_mul_12_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_mul_loop_mul_12_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_mul_loop_mul_12_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_sva_2)
    );
  SDP_X_leading_sign_23_0 mul_loop_mul_12_leading_sign_23_0_rg (
      .mantissa(nl_mul_loop_mul_12_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_27)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) mul_loop_mul_13_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_mul_loop_mul_13_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_mul_loop_mul_13_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_sva_2)
    );
  SDP_X_leading_sign_23_0 mul_loop_mul_13_leading_sign_23_0_rg (
      .mantissa(nl_mul_loop_mul_13_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_28)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) mul_loop_mul_14_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_mul_loop_mul_14_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_mul_loop_mul_14_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_sva_2)
    );
  SDP_X_leading_sign_23_0 mul_loop_mul_14_leading_sign_23_0_rg (
      .mantissa(nl_mul_loop_mul_14_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_29)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) mul_loop_mul_15_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_mul_loop_mul_15_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_mul_loop_mul_15_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_sva_2)
    );
  SDP_X_leading_sign_23_0 mul_loop_mul_15_leading_sign_23_0_rg (
      .mantissa(nl_mul_loop_mul_15_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_30)
    );
  SDP_X_mgc_shift_l_v4 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd23)) mul_loop_mul_16_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_mul_loop_mul_16_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_a[21:0]),
      .s(nl_mul_loop_mul_16_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_lshift_rg_s[5:0]),
      .z(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_sva_2)
    );
  SDP_X_leading_sign_23_0 mul_loop_mul_16_leading_sign_23_0_rg (
      .mantissa(nl_mul_loop_mul_16_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_31)
    );
  SDP_X_X_mul_core_chn_mul_in_rsci X_mul_core_chn_mul_in_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_in_rsc_slz(chn_mul_in_rsc_slz),
      .chn_mul_in_rsc_sz(chn_mul_in_rsc_sz),
      .chn_mul_in_rsc_z(chn_mul_in_rsc_z),
      .chn_mul_in_rsc_vz(chn_mul_in_rsc_vz),
      .chn_mul_in_rsc_lz(chn_mul_in_rsc_lz),
      .chn_mul_in_rsci_oswt(chn_mul_in_rsci_oswt),
      .core_wen(core_wen),
      .chn_mul_in_rsci_iswt0(chn_mul_in_rsci_iswt0),
      .chn_mul_in_rsci_bawt(chn_mul_in_rsci_bawt),
      .chn_mul_in_rsci_wen_comp(chn_mul_in_rsci_wen_comp),
      .chn_mul_in_rsci_ld_core_psct(chn_mul_in_rsci_ld_core_psct),
      .chn_mul_in_rsci_d_mxwt(chn_mul_in_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  SDP_X_X_mul_core_chn_mul_op_rsci X_mul_core_chn_mul_op_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_op_rsc_z(chn_mul_op_rsc_z),
      .chn_mul_op_rsc_vz(chn_mul_op_rsc_vz),
      .chn_mul_op_rsc_lz(chn_mul_op_rsc_lz),
      .chn_mul_op_rsci_oswt(chn_mul_op_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_mul_op_rsci_iswt0(chn_mul_op_rsci_iswt0),
      .chn_mul_op_rsci_bawt(chn_mul_op_rsci_bawt),
      .chn_mul_op_rsci_wen_comp(chn_mul_op_rsci_wen_comp),
      .chn_mul_op_rsci_ld_core_psct(chn_mul_op_rsci_ld_core_psct),
      .chn_mul_op_rsci_d_mxwt(chn_mul_op_rsci_d_mxwt)
    );
  SDP_X_X_mul_core_chn_mul_out_rsci X_mul_core_chn_mul_out_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_out_rsc_z(chn_mul_out_rsc_z),
      .chn_mul_out_rsc_vz(chn_mul_out_rsc_vz),
      .chn_mul_out_rsc_lz(chn_mul_out_rsc_lz),
      .chn_mul_out_rsci_oswt(chn_mul_out_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_mul_out_rsci_iswt0(chn_mul_out_rsci_iswt0),
      .chn_mul_out_rsci_bawt(chn_mul_out_rsci_bawt),
      .chn_mul_out_rsci_wen_comp(chn_mul_out_rsci_wen_comp),
      .chn_mul_out_rsci_ld_core_psct(reg_chn_mul_out_rsci_ld_core_psct_cse),
      .chn_mul_out_rsci_d(nl_X_mul_core_chn_mul_out_rsci_inst_chn_mul_out_rsci_d[799:0])
    );
  SDP_X_X_mul_core_cfg_mul_op_rsc_triosy_obj X_mul_core_cfg_mul_op_rsc_triosy_obj_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_mul_op_rsc_triosy_lz(cfg_mul_op_rsc_triosy_lz),
      .cfg_mul_op_rsc_triosy_obj_oswt(cfg_mul_op_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_mul_op_rsc_triosy_obj_iswt0(reg_cfg_mul_src_rsc_triosy_obj_ld_core_psct_cse),
      .cfg_mul_op_rsc_triosy_obj_bawt(cfg_mul_op_rsc_triosy_obj_bawt)
    );
  SDP_X_X_mul_core_cfg_mul_bypass_rsc_triosy_obj X_mul_core_cfg_mul_bypass_rsc_triosy_obj_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_mul_bypass_rsc_triosy_lz(cfg_mul_bypass_rsc_triosy_lz),
      .cfg_mul_bypass_rsc_triosy_obj_oswt(cfg_mul_bypass_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_mul_bypass_rsc_triosy_obj_iswt0(reg_cfg_mul_src_rsc_triosy_obj_ld_core_psct_cse),
      .cfg_mul_bypass_rsc_triosy_obj_bawt(cfg_mul_bypass_rsc_triosy_obj_bawt)
    );
  SDP_X_X_mul_core_cfg_mul_prelu_rsc_triosy_obj X_mul_core_cfg_mul_prelu_rsc_triosy_obj_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_mul_prelu_rsc_triosy_lz(cfg_mul_prelu_rsc_triosy_lz),
      .cfg_mul_prelu_rsc_triosy_obj_oswt(cfg_mul_prelu_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_mul_prelu_rsc_triosy_obj_iswt0(reg_cfg_mul_src_rsc_triosy_obj_ld_core_psct_cse),
      .cfg_mul_prelu_rsc_triosy_obj_bawt(cfg_mul_prelu_rsc_triosy_obj_bawt)
    );
  SDP_X_X_mul_core_cfg_mul_src_rsc_triosy_obj X_mul_core_cfg_mul_src_rsc_triosy_obj_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_mul_src_rsc_triosy_lz(cfg_mul_src_rsc_triosy_lz),
      .cfg_mul_src_rsc_triosy_obj_oswt(cfg_mul_src_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_mul_src_rsc_triosy_obj_iswt0(reg_cfg_mul_src_rsc_triosy_obj_ld_core_psct_cse),
      .cfg_mul_src_rsc_triosy_obj_bawt(cfg_mul_src_rsc_triosy_obj_bawt)
    );
  SDP_X_X_mul_core_staller X_mul_core_staller_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .chn_mul_in_rsci_wen_comp(chn_mul_in_rsci_wen_comp),
      .core_wten(core_wten),
      .chn_mul_op_rsci_wen_comp(chn_mul_op_rsci_wen_comp),
      .chn_mul_out_rsci_wen_comp(chn_mul_out_rsci_wen_comp)
    );
  SDP_X_X_mul_core_core_fsm X_mul_core_core_fsm_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign iExpoWidth_oExpoWidth_prb = mul_loop_mul_1_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL mul_loop_mul_1_X_mul_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb = mul_loop_mul_1_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL mul_loop_mul_1_X_mul_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_1 = mul_loop_mul_1_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL mul_loop_mul_1_X_mul_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_1 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_1 = mul_loop_mul_1_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL mul_loop_mul_1_X_mul_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_1 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_2 = mul_loop_mul_1_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL mul_loop_mul_1_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_2 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_2 = mul_loop_mul_2_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL mul_loop_mul_2_X_mul_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_2 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_3 = mul_loop_mul_2_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL mul_loop_mul_2_X_mul_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_3 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_4 = mul_loop_mul_2_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL mul_loop_mul_2_X_mul_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_4 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_3 = mul_loop_mul_2_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL mul_loop_mul_2_X_mul_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_3 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_5 = mul_loop_mul_2_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL mul_loop_mul_2_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_5 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_4 = mul_loop_mul_3_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL mul_loop_mul_3_X_mul_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_4 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_6 = mul_loop_mul_3_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL mul_loop_mul_3_X_mul_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_6 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_7 = mul_loop_mul_3_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL mul_loop_mul_3_X_mul_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_7 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_5 = mul_loop_mul_3_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL mul_loop_mul_3_X_mul_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_5 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_8 = mul_loop_mul_3_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL mul_loop_mul_3_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_8 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_6 = mul_loop_mul_4_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL mul_loop_mul_4_X_mul_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_6 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_9 = mul_loop_mul_4_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL mul_loop_mul_4_X_mul_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_9 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_10 = mul_loop_mul_4_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL mul_loop_mul_4_X_mul_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_10 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_7 = mul_loop_mul_4_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL mul_loop_mul_4_X_mul_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_7 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_11 = mul_loop_mul_4_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL mul_loop_mul_4_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_11 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_8 = mul_loop_mul_5_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL mul_loop_mul_5_X_mul_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_8 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_12 = mul_loop_mul_5_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL mul_loop_mul_5_X_mul_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_12 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_13 = mul_loop_mul_5_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL mul_loop_mul_5_X_mul_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_13 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_9 = mul_loop_mul_5_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL mul_loop_mul_5_X_mul_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_9 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_14 = mul_loop_mul_5_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL mul_loop_mul_5_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_14 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_10 = mul_loop_mul_6_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL mul_loop_mul_6_X_mul_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_10 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_15 = mul_loop_mul_6_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL mul_loop_mul_6_X_mul_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_15 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_16 = mul_loop_mul_6_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL mul_loop_mul_6_X_mul_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_16 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_11 = mul_loop_mul_6_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL mul_loop_mul_6_X_mul_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_11 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_17 = mul_loop_mul_6_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL mul_loop_mul_6_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_17 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_12 = mul_loop_mul_7_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL mul_loop_mul_7_X_mul_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_12 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_18 = mul_loop_mul_7_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL mul_loop_mul_7_X_mul_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_18 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_19 = mul_loop_mul_7_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL mul_loop_mul_7_X_mul_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_19 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_13 = mul_loop_mul_7_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL mul_loop_mul_7_X_mul_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_13 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_20 = mul_loop_mul_7_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL mul_loop_mul_7_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_20 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_14 = mul_loop_mul_8_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL mul_loop_mul_8_X_mul_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_14 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_21 = mul_loop_mul_8_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL mul_loop_mul_8_X_mul_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_21 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_22 = mul_loop_mul_8_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL mul_loop_mul_8_X_mul_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_22 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_15 = mul_loop_mul_8_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL mul_loop_mul_8_X_mul_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_15 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_23 = mul_loop_mul_8_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL mul_loop_mul_8_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_23 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_16 = mul_loop_mul_9_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL mul_loop_mul_9_X_mul_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_16 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_24 = mul_loop_mul_9_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL mul_loop_mul_9_X_mul_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_24 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_25 = mul_loop_mul_9_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL mul_loop_mul_9_X_mul_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_25 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_17 = mul_loop_mul_9_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL mul_loop_mul_9_X_mul_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_17 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_26 = mul_loop_mul_9_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL mul_loop_mul_9_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_26 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_18 = mul_loop_mul_10_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL mul_loop_mul_10_X_mul_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_18 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_27 = mul_loop_mul_10_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL mul_loop_mul_10_X_mul_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_27 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_28 = mul_loop_mul_10_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL mul_loop_mul_10_X_mul_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_28 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_19 = mul_loop_mul_10_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL mul_loop_mul_10_X_mul_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_19 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_29 = mul_loop_mul_10_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL mul_loop_mul_10_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_29 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_20 = mul_loop_mul_11_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL mul_loop_mul_11_X_mul_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_20 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_30 = mul_loop_mul_11_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL mul_loop_mul_11_X_mul_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_30 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_31 = mul_loop_mul_11_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL mul_loop_mul_11_X_mul_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_31 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_21 = mul_loop_mul_11_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL mul_loop_mul_11_X_mul_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_21 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_32 = mul_loop_mul_11_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL mul_loop_mul_11_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_32 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_22 = mul_loop_mul_12_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL mul_loop_mul_12_X_mul_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_22 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_33 = mul_loop_mul_12_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL mul_loop_mul_12_X_mul_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_33 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_34 = mul_loop_mul_12_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL mul_loop_mul_12_X_mul_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_34 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_23 = mul_loop_mul_12_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL mul_loop_mul_12_X_mul_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_23 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_35 = mul_loop_mul_12_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL mul_loop_mul_12_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_35 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_24 = mul_loop_mul_13_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL mul_loop_mul_13_X_mul_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_24 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_36 = mul_loop_mul_13_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL mul_loop_mul_13_X_mul_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_36 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_37 = mul_loop_mul_13_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL mul_loop_mul_13_X_mul_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_37 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_25 = mul_loop_mul_13_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL mul_loop_mul_13_X_mul_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_25 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_38 = mul_loop_mul_13_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL mul_loop_mul_13_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_38 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_26 = mul_loop_mul_14_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL mul_loop_mul_14_X_mul_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_26 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_39 = mul_loop_mul_14_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL mul_loop_mul_14_X_mul_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_39 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_40 = mul_loop_mul_14_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL mul_loop_mul_14_X_mul_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_40 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_27 = mul_loop_mul_14_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL mul_loop_mul_14_X_mul_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_27 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_41 = mul_loop_mul_14_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL mul_loop_mul_14_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_41 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_28 = mul_loop_mul_15_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL mul_loop_mul_15_X_mul_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_28 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_42 = mul_loop_mul_15_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL mul_loop_mul_15_X_mul_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_42 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_43 = mul_loop_mul_15_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL mul_loop_mul_15_X_mul_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_43 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_29 = mul_loop_mul_15_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL mul_loop_mul_15_X_mul_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_29 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_44 = mul_loop_mul_15_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL mul_loop_mul_15_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_44 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_30 = mul_loop_mul_16_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL mul_loop_mul_16_X_mul_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_30 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_45 = mul_loop_mul_16_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL mul_loop_mul_16_X_mul_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_45 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_46 = mul_loop_mul_16_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL mul_loop_mul_16_X_mul_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_46 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_31 = mul_loop_mul_16_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL mul_loop_mul_16_X_mul_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_31 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_47 = mul_loop_mul_16_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL mul_loop_mul_16_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_47 } @rose(nvdla_core_clk);
  assign and_2496_cse = (~(IsNaN_8U_23U_1_land_1_lpi_1_dfm_9 | IsNaN_8U_23U_land_1_lpi_1_dfm_11))
      & and_116_ssc;
  assign and_2497_cse = IsNaN_8U_23U_1_land_1_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_1_lpi_1_dfm_11)
      & and_116_ssc;
  assign or_4733_cse = (IsNaN_8U_23U_land_1_lpi_1_dfm_11 & and_116_ssc) | or_17_ssc;
  assign chn_mul_out_and_cse = core_wen & (~(and_dcpl_50 | (~ main_stage_v_4)));
  assign and_2488_cse = (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_9) & asn_1165;
  assign and_2489_cse = IsNaN_8U_23U_1_land_1_lpi_1_dfm_9 & asn_1165;
  assign and_2481_cse = (~(IsNaN_8U_23U_1_land_2_lpi_1_dfm_9 | IsNaN_8U_23U_land_2_lpi_1_dfm_11))
      & and_51_ssc;
  assign and_2482_cse = IsNaN_8U_23U_1_land_2_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_2_lpi_1_dfm_11)
      & and_51_ssc;
  assign or_4729_cse = (IsNaN_8U_23U_land_2_lpi_1_dfm_11 & and_51_ssc) | or_1_ssc;
  assign and_2473_cse = (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_9) & asn_1175;
  assign and_2474_cse = IsNaN_8U_23U_1_land_2_lpi_1_dfm_9 & asn_1175;
  assign and_2466_cse = (~(IsNaN_8U_23U_1_land_3_lpi_1_dfm_9 | IsNaN_8U_23U_land_3_lpi_1_dfm_11))
      & and_55_ssc;
  assign and_2467_cse = IsNaN_8U_23U_1_land_3_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_3_lpi_1_dfm_11)
      & and_55_ssc;
  assign or_4725_cse = (IsNaN_8U_23U_land_3_lpi_1_dfm_11 & and_55_ssc) | or_2_ssc;
  assign and_2458_cse = (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_9) & asn_1185;
  assign and_2459_cse = IsNaN_8U_23U_1_land_3_lpi_1_dfm_9 & asn_1185;
  assign and_2451_cse = (~(IsNaN_8U_23U_1_land_4_lpi_1_dfm_9 | IsNaN_8U_23U_land_4_lpi_1_dfm_11))
      & and_59_ssc;
  assign and_2452_cse = IsNaN_8U_23U_1_land_4_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_4_lpi_1_dfm_11)
      & and_59_ssc;
  assign or_4721_cse = (IsNaN_8U_23U_land_4_lpi_1_dfm_11 & and_59_ssc) | or_3_ssc;
  assign and_2443_cse = (~ IsNaN_8U_23U_1_land_4_lpi_1_dfm_9) & asn_1195;
  assign and_2444_cse = IsNaN_8U_23U_1_land_4_lpi_1_dfm_9 & asn_1195;
  assign and_2436_cse = (~(IsNaN_8U_23U_1_land_5_lpi_1_dfm_9 | IsNaN_8U_23U_land_5_lpi_1_dfm_11))
      & and_63_ssc;
  assign and_2437_cse = IsNaN_8U_23U_1_land_5_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_5_lpi_1_dfm_11)
      & and_63_ssc;
  assign or_4717_cse = (IsNaN_8U_23U_land_5_lpi_1_dfm_11 & and_63_ssc) | or_4_ssc;
  assign and_2428_cse = (~ IsNaN_8U_23U_1_land_5_lpi_1_dfm_9) & asn_1205;
  assign and_2429_cse = IsNaN_8U_23U_1_land_5_lpi_1_dfm_9 & asn_1205;
  assign and_2421_cse = (~(IsNaN_8U_23U_1_land_6_lpi_1_dfm_9 | IsNaN_8U_23U_land_6_lpi_1_dfm_11))
      & and_67_ssc;
  assign and_2422_cse = IsNaN_8U_23U_1_land_6_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_6_lpi_1_dfm_11)
      & and_67_ssc;
  assign or_4713_cse = (IsNaN_8U_23U_land_6_lpi_1_dfm_11 & and_67_ssc) | or_5_ssc;
  assign and_2413_cse = (~ IsNaN_8U_23U_1_land_6_lpi_1_dfm_9) & asn_1215;
  assign and_2414_cse = IsNaN_8U_23U_1_land_6_lpi_1_dfm_9 & asn_1215;
  assign and_2406_cse = (~(IsNaN_8U_23U_1_land_7_lpi_1_dfm_9 | IsNaN_8U_23U_land_7_lpi_1_dfm_11))
      & and_71_ssc;
  assign and_2407_cse = IsNaN_8U_23U_1_land_7_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_7_lpi_1_dfm_11)
      & and_71_ssc;
  assign or_4709_cse = (IsNaN_8U_23U_land_7_lpi_1_dfm_11 & and_71_ssc) | or_6_ssc;
  assign and_2398_cse = (~ IsNaN_8U_23U_1_land_7_lpi_1_dfm_9) & asn_1225;
  assign and_2399_cse = IsNaN_8U_23U_1_land_7_lpi_1_dfm_9 & asn_1225;
  assign and_2391_cse = (~(IsNaN_8U_23U_1_land_8_lpi_1_dfm_9 | IsNaN_8U_23U_land_8_lpi_1_dfm_11))
      & and_75_ssc;
  assign and_2392_cse = IsNaN_8U_23U_1_land_8_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_8_lpi_1_dfm_11)
      & and_75_ssc;
  assign or_4705_cse = (IsNaN_8U_23U_land_8_lpi_1_dfm_11 & and_75_ssc) | or_7_ssc;
  assign and_2383_cse = (~ IsNaN_8U_23U_1_land_8_lpi_1_dfm_9) & asn_1235;
  assign and_2384_cse = IsNaN_8U_23U_1_land_8_lpi_1_dfm_9 & asn_1235;
  assign and_2376_cse = (~(IsNaN_8U_23U_1_land_9_lpi_1_dfm_9 | IsNaN_8U_23U_land_9_lpi_1_dfm_11))
      & and_79_ssc;
  assign and_2377_cse = IsNaN_8U_23U_1_land_9_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_9_lpi_1_dfm_11)
      & and_79_ssc;
  assign or_4701_cse = (IsNaN_8U_23U_land_9_lpi_1_dfm_11 & and_79_ssc) | or_8_ssc;
  assign and_2368_cse = (~ IsNaN_8U_23U_1_land_9_lpi_1_dfm_9) & asn_1245;
  assign and_2369_cse = IsNaN_8U_23U_1_land_9_lpi_1_dfm_9 & asn_1245;
  assign and_2361_cse = (~(IsNaN_8U_23U_1_land_10_lpi_1_dfm_9 | IsNaN_8U_23U_land_10_lpi_1_dfm_11))
      & and_83_ssc;
  assign and_2362_cse = IsNaN_8U_23U_1_land_10_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_10_lpi_1_dfm_11)
      & and_83_ssc;
  assign or_4697_cse = (IsNaN_8U_23U_land_10_lpi_1_dfm_11 & and_83_ssc) | or_9_ssc;
  assign and_2353_cse = (~ IsNaN_8U_23U_1_land_10_lpi_1_dfm_9) & asn_1255;
  assign and_2354_cse = IsNaN_8U_23U_1_land_10_lpi_1_dfm_9 & asn_1255;
  assign and_2346_cse = (~(IsNaN_8U_23U_1_land_11_lpi_1_dfm_9 | IsNaN_8U_23U_land_11_lpi_1_dfm_11))
      & and_87_ssc;
  assign and_2347_cse = IsNaN_8U_23U_1_land_11_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_11_lpi_1_dfm_11)
      & and_87_ssc;
  assign or_4693_cse = (IsNaN_8U_23U_land_11_lpi_1_dfm_11 & and_87_ssc) | or_10_ssc;
  assign and_2338_cse = (~ IsNaN_8U_23U_1_land_11_lpi_1_dfm_9) & asn_1265;
  assign and_2339_cse = IsNaN_8U_23U_1_land_11_lpi_1_dfm_9 & asn_1265;
  assign and_2331_cse = (~(IsNaN_8U_23U_1_land_12_lpi_1_dfm_9 | IsNaN_8U_23U_land_12_lpi_1_dfm_11))
      & and_91_ssc;
  assign and_2332_cse = IsNaN_8U_23U_1_land_12_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_12_lpi_1_dfm_11)
      & and_91_ssc;
  assign or_4689_cse = (IsNaN_8U_23U_land_12_lpi_1_dfm_11 & and_91_ssc) | or_11_ssc;
  assign and_2323_cse = (~ IsNaN_8U_23U_1_land_12_lpi_1_dfm_9) & asn_1275;
  assign and_2324_cse = IsNaN_8U_23U_1_land_12_lpi_1_dfm_9 & asn_1275;
  assign and_2316_cse = (~(IsNaN_8U_23U_1_land_13_lpi_1_dfm_9 | IsNaN_8U_23U_land_13_lpi_1_dfm_11))
      & and_95_ssc;
  assign and_2317_cse = IsNaN_8U_23U_1_land_13_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_13_lpi_1_dfm_11)
      & and_95_ssc;
  assign or_4685_cse = (IsNaN_8U_23U_land_13_lpi_1_dfm_11 & and_95_ssc) | or_12_ssc;
  assign and_2308_cse = (~ IsNaN_8U_23U_1_land_13_lpi_1_dfm_9) & asn_1285;
  assign and_2309_cse = IsNaN_8U_23U_1_land_13_lpi_1_dfm_9 & asn_1285;
  assign and_2301_cse = (~(IsNaN_8U_23U_1_land_14_lpi_1_dfm_9 | IsNaN_8U_23U_land_14_lpi_1_dfm_11))
      & and_99_ssc;
  assign and_2302_cse = IsNaN_8U_23U_1_land_14_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_14_lpi_1_dfm_11)
      & and_99_ssc;
  assign or_4681_cse = (IsNaN_8U_23U_land_14_lpi_1_dfm_11 & and_99_ssc) | or_13_ssc;
  assign and_2293_cse = (~ IsNaN_8U_23U_1_land_14_lpi_1_dfm_9) & asn_1295;
  assign and_2294_cse = IsNaN_8U_23U_1_land_14_lpi_1_dfm_9 & asn_1295;
  assign and_2286_cse = (~(IsNaN_8U_23U_1_land_15_lpi_1_dfm_9 | IsNaN_8U_23U_land_15_lpi_1_dfm_11))
      & and_103_ssc;
  assign and_2287_cse = IsNaN_8U_23U_1_land_15_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_15_lpi_1_dfm_11)
      & and_103_ssc;
  assign or_4677_cse = (IsNaN_8U_23U_land_15_lpi_1_dfm_11 & and_103_ssc) | or_14_ssc;
  assign and_2278_cse = (~ IsNaN_8U_23U_1_land_15_lpi_1_dfm_9) & asn_1305;
  assign and_2279_cse = IsNaN_8U_23U_1_land_15_lpi_1_dfm_9 & asn_1305;
  assign and_2271_cse = (~(IsNaN_8U_23U_1_land_lpi_1_dfm_9 | IsNaN_8U_23U_land_lpi_1_dfm_11))
      & and_107_ssc;
  assign and_2272_cse = IsNaN_8U_23U_1_land_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_lpi_1_dfm_11)
      & and_107_ssc;
  assign or_4673_cse = (IsNaN_8U_23U_land_lpi_1_dfm_11 & and_107_ssc) | or_15_ssc;
  assign and_2263_cse = (~ IsNaN_8U_23U_1_land_lpi_1_dfm_9) & asn_1315;
  assign and_2264_cse = IsNaN_8U_23U_1_land_lpi_1_dfm_9 & asn_1315;
  assign or_90_cse = (cfg_precision!=2'b10);
  assign nor_21_cse = ~((chn_mul_in_rsci_d_mxwt[31]) | (~ cfg_mul_prelu_rsci_d));
  assign IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_31_cse = (and_dcpl_7 & and_dcpl_85)
      | and_dcpl_87;
  assign nor_23_cse = ~((chn_mul_in_rsci_d_mxwt[64]) | (~ cfg_mul_prelu_rsci_d));
  assign nor_25_cse = ~((chn_mul_in_rsci_d_mxwt[97]) | (~ cfg_mul_prelu_rsci_d));
  assign nor_26_cse = ~((chn_mul_in_rsci_d_mxwt[130]) | (~ cfg_mul_prelu_rsci_d));
  assign nor_28_cse = ~((chn_mul_in_rsci_d_mxwt[163]) | (~ cfg_mul_prelu_rsci_d));
  assign nor_29_cse = ~((chn_mul_in_rsci_d_mxwt[196]) | (~ cfg_mul_prelu_rsci_d));
  assign nor_30_cse = ~((chn_mul_in_rsci_d_mxwt[229]) | (~ cfg_mul_prelu_rsci_d));
  assign nor_32_cse = ~((chn_mul_in_rsci_d_mxwt[262]) | (~ cfg_mul_prelu_rsci_d));
  assign nor_34_cse = ~((chn_mul_in_rsci_d_mxwt[295]) | (~ cfg_mul_prelu_rsci_d));
  assign nor_35_cse = ~((chn_mul_in_rsci_d_mxwt[328]) | (~ cfg_mul_prelu_rsci_d));
  assign nor_36_cse = ~((chn_mul_in_rsci_d_mxwt[361]) | (~ cfg_mul_prelu_rsci_d));
  assign nor_37_cse = ~((chn_mul_in_rsci_d_mxwt[394]) | (~ cfg_mul_prelu_rsci_d));
  assign nor_39_cse = ~((chn_mul_in_rsci_d_mxwt[427]) | (~ cfg_mul_prelu_rsci_d));
  assign nor_40_cse = ~((chn_mul_in_rsci_d_mxwt[460]) | (~ cfg_mul_prelu_rsci_d));
  assign nor_42_cse = ~((chn_mul_in_rsci_d_mxwt[493]) | (~ cfg_mul_prelu_rsci_d));
  assign nor_44_cse = ~((chn_mul_in_rsci_d_mxwt[526]) | (~ cfg_mul_prelu_rsci_d));
  assign nand_26_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 & (~(cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & or_309_cse)));
  assign mux_152_nl = MUX_s_1_2_2(or_309_cse, (nand_26_nl), main_stage_v_1);
  assign mux_153_nl = MUX_s_1_2_2(or_tmp_115, (~ (mux_152_nl)), chn_mul_in_rsci_bawt);
  assign mux_154_nl = MUX_s_1_2_2((mux_153_nl), or_tmp_115, cfg_mul_bypass_rsci_d);
  assign mul_loop_mul_if_aelse_and_16_cse = core_wen & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_31_cse
      & (~ (mux_154_nl));
  assign cfg_mul_op_and_cse = core_wen & (~ or_dcpl_46);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_48_cse = core_wen & ((and_dcpl_100
      & (~ mul_loop_mul_if_land_1_lpi_1_dfm_st_5) & (cfg_precision==2'b10)) | and_dcpl_102)
      & mux_tmp_148;
  assign MulIn_data_and_cse = core_wen & (~ and_dcpl_50) & mux_tmp_148;
  assign FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse = (or_309_cse & and_dcpl_85)
      | and_dcpl_104;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_51_cse = core_wen & ((and_dcpl_100
      & (~ mul_loop_mul_if_land_2_lpi_1_dfm_st_5) & (cfg_precision==2'b10)) | and_dcpl_108)
      & mux_tmp_148;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_54_cse = core_wen & ((and_dcpl_100
      & (~ mul_loop_mul_if_land_3_lpi_1_dfm_st_5) & (cfg_precision==2'b10)) | and_dcpl_112)
      & mux_tmp_148;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_57_cse = core_wen & ((and_dcpl_100
      & (~ mul_loop_mul_if_land_4_lpi_1_dfm_st_5) & (cfg_precision==2'b10)) | and_dcpl_116)
      & mux_tmp_148;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_60_cse = core_wen & ((and_dcpl_100
      & (~ mul_loop_mul_if_land_5_lpi_1_dfm_st_5) & (cfg_precision==2'b10)) | and_dcpl_120)
      & mux_tmp_148;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_63_cse = core_wen & ((and_dcpl_100
      & (~ mul_loop_mul_if_land_6_lpi_1_dfm_st_5) & (cfg_precision==2'b10)) | and_dcpl_124)
      & mux_tmp_148;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_66_cse = core_wen & ((and_dcpl_100
      & (~ mul_loop_mul_if_land_7_lpi_1_dfm_st_5) & (cfg_precision==2'b10)) | and_dcpl_128)
      & mux_tmp_148;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_69_cse = core_wen & ((and_dcpl_100
      & (~ mul_loop_mul_if_land_8_lpi_1_dfm_st_5) & (cfg_precision==2'b10)) | and_dcpl_132)
      & mux_tmp_148;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_72_cse = core_wen & ((and_dcpl_100
      & (~ mul_loop_mul_if_land_9_lpi_1_dfm_st_5) & (cfg_precision==2'b10)) | and_dcpl_136)
      & mux_tmp_148;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_75_cse = core_wen & ((and_dcpl_100
      & (~ mul_loop_mul_if_land_10_lpi_1_dfm_st_5) & (cfg_precision==2'b10)) | and_dcpl_140)
      & mux_tmp_148;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_78_cse = core_wen & ((and_dcpl_100
      & (~ mul_loop_mul_if_land_11_lpi_1_dfm_st_5) & (cfg_precision==2'b10)) | and_dcpl_144)
      & mux_tmp_148;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_81_cse = core_wen & ((and_dcpl_100
      & (~ mul_loop_mul_if_land_12_lpi_1_dfm_st_5) & (cfg_precision==2'b10)) | and_dcpl_148)
      & mux_tmp_148;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_84_cse = core_wen & ((and_dcpl_100
      & (~ mul_loop_mul_if_land_13_lpi_1_dfm_st_5) & (cfg_precision==2'b10)) | and_dcpl_152)
      & mux_tmp_148;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_87_cse = core_wen & ((and_dcpl_100
      & (~ mul_loop_mul_if_land_14_lpi_1_dfm_st_5) & (cfg_precision==2'b10)) | and_dcpl_156)
      & mux_tmp_148;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_90_cse = core_wen & ((and_dcpl_100
      & (~ mul_loop_mul_if_land_15_lpi_1_dfm_st_5) & (cfg_precision==2'b10)) | and_dcpl_160)
      & mux_tmp_148;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_93_cse = core_wen & ((and_dcpl_100
      & (~ mul_loop_mul_if_land_lpi_1_dfm_st_5) & (cfg_precision==2'b10)) | and_dcpl_164)
      & mux_tmp_148;
  assign mux_172_nl = MUX_s_1_2_2(or_tmp_204, or_tmp_139, or_309_cse);
  assign mul_loop_mul_if_aelse_and_32_cse = core_wen & (~ and_dcpl_50) & (~ (mux_172_nl));
  assign nor_1492_nl = ~(mul_loop_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_1_lpi_1_dfm_st_6);
  assign mux_173_nl = MUX_s_1_2_2((nor_1492_nl), nor_821_cse, reg_FpMul_8U_23U_lor_3_lpi_1_dfm_4_cse);
  assign and_2249_nl = nor_50_cse & (mux_173_nl);
  assign nor_1493_nl = ~((~ mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_18_lpi_1_dfm_st | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_1_lpi_1_dfm_st_6);
  assign mux_174_nl = MUX_s_1_2_2((nor_1493_nl), (and_2249_nl), nor_53_cse);
  assign mux_175_nl = MUX_s_1_2_2(nor_129_cse, (mux_174_nl), or_309_cse);
  assign IsZero_8U_23U_aelse_and_32_cse = core_wen & (~ and_dcpl_50) & (mux_175_nl);
  assign mux_176_nl = MUX_s_1_2_2(main_stage_v_3, main_stage_v_2, or_309_cse);
  assign MulIn_data_and_1_cse = core_wen & (~ and_dcpl_50) & (mux_176_nl);
  assign mux_178_nl = MUX_s_1_2_2(or_2576_cse, or_tmp_213, mul_loop_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_179_nl = MUX_s_1_2_2((mux_178_nl), or_2576_cse, reg_FpMul_8U_23U_lor_3_lpi_1_dfm_4_cse);
  assign mux_180_nl = MUX_s_1_2_2(or_tmp_213, (mux_179_nl), nor_50_cse);
  assign mux_181_nl = MUX_s_1_2_2(or_2576_cse, or_tmp_213, or_2577_cse);
  assign mux_182_nl = MUX_s_1_2_2((mux_181_nl), (mux_180_nl), nor_53_cse);
  assign or_308_nl = (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_1_lpi_1_dfm_st_7
      | ((IsNaN_8U_23U_land_1_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | (~
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_8) | mul_loop_mul_if_land_1_lpi_1_dfm_9) &
      or_4383_cse);
  assign mux_183_nl = MUX_s_1_2_2((or_308_nl), (mux_182_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_48_cse = core_wen & (~ and_dcpl_50)
      & (~ (mux_183_nl));
  assign or_309_cse = (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt;
  assign nor_53_cse = ~((cfg_precision!=2'b10));
  assign nor_1490_cse = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_1_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_18_lpi_1_dfm_st_3);
  assign or_312_cse = mul_loop_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_3_lpi_1_dfm_4_cse;
  assign FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_31_cse = MUX_s_1_2_2(or_312_cse,
      FpMul_8U_23U_lor_18_lpi_1_dfm_st, and_dcpl_104);
  assign nor_1481_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_2_lpi_1_dfm_st_6);
  assign nor_1482_nl = ~(mul_loop_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_2_lpi_1_dfm_st_6);
  assign mux_188_nl = MUX_s_1_2_2((nor_1482_nl), (nor_1481_nl), reg_FpMul_8U_23U_lor_4_lpi_1_dfm_4_cse);
  assign and_2248_nl = nor_55_cse & (mux_188_nl);
  assign nor_1483_nl = ~((~ mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_19_lpi_1_dfm_st | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_2_lpi_1_dfm_st_6);
  assign mux_189_nl = MUX_s_1_2_2((nor_1483_nl), (and_2248_nl), nor_53_cse);
  assign mux_190_nl = MUX_s_1_2_2(nor_145_cse, (mux_189_nl), or_309_cse);
  assign IsZero_8U_23U_aelse_and_33_cse = core_wen & (~ and_dcpl_50) & (mux_190_nl);
  assign mux_192_nl = MUX_s_1_2_2(or_2607_cse, or_tmp_236, mul_loop_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_193_nl = MUX_s_1_2_2((mux_192_nl), or_2607_cse, reg_FpMul_8U_23U_lor_4_lpi_1_dfm_4_cse);
  assign mux_194_nl = MUX_s_1_2_2(or_tmp_236, (mux_193_nl), nor_55_cse);
  assign mux_195_nl = MUX_s_1_2_2(or_2607_cse, or_tmp_236, or_2608_cse);
  assign mux_196_nl = MUX_s_1_2_2((mux_195_nl), (mux_194_nl), nor_53_cse);
  assign or_331_nl = (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_2_lpi_1_dfm_st_7
      | ((IsNaN_8U_23U_land_2_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | (~
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_8) | mul_loop_mul_if_land_2_lpi_1_dfm_9) &
      or_4384_cse);
  assign mux_197_nl = MUX_s_1_2_2((or_331_nl), (mux_196_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_51_cse = core_wen & (~ and_dcpl_50)
      & (~ (mux_197_nl));
  assign FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_30_cse = MUX_s_1_2_2(or_2628_cse,
      FpMul_8U_23U_lor_19_lpi_1_dfm_st, and_dcpl_104);
  assign nor_1477_cse = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_3_lpi_1_dfm_st_6);
  assign nor_1478_nl = ~(mul_loop_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_3_lpi_1_dfm_st_6);
  assign mux_203_nl = MUX_s_1_2_2((nor_1478_nl), nor_1477_cse, reg_FpMul_8U_23U_lor_5_lpi_1_dfm_4_cse);
  assign and_2247_nl = nor_59_cse & (mux_203_nl);
  assign nor_1479_nl = ~((~ mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_20_lpi_1_dfm_st | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_3_lpi_1_dfm_st_6);
  assign mux_204_nl = MUX_s_1_2_2((nor_1479_nl), (and_2247_nl), nor_53_cse);
  assign mux_205_nl = MUX_s_1_2_2(nor_161_cse, (mux_204_nl), or_309_cse);
  assign IsZero_8U_23U_aelse_and_34_cse = core_wen & (~ and_dcpl_50) & (mux_205_nl);
  assign mux_207_nl = MUX_s_1_2_2(or_2630_cse, or_tmp_264, mul_loop_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_208_nl = MUX_s_1_2_2((mux_207_nl), or_2630_cse, reg_FpMul_8U_23U_lor_5_lpi_1_dfm_4_cse);
  assign mux_209_nl = MUX_s_1_2_2(or_tmp_264, (mux_208_nl), nor_59_cse);
  assign mux_210_nl = MUX_s_1_2_2(or_2630_cse, or_tmp_264, or_2631_cse);
  assign mux_211_nl = MUX_s_1_2_2((mux_210_nl), (mux_209_nl), nor_53_cse);
  assign or_359_nl = (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_3_lpi_1_dfm_st_7
      | ((IsNaN_8U_23U_land_3_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | (~
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_8) | mul_loop_mul_if_land_3_lpi_1_dfm_9) &
      or_4385_cse);
  assign mux_212_nl = MUX_s_1_2_2((or_359_nl), (mux_211_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_54_cse = core_wen & (~ and_dcpl_50)
      & (~ (mux_212_nl));
  assign or_363_cse = mul_loop_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_5_lpi_1_dfm_4_cse;
  assign FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_29_cse = MUX_s_1_2_2(or_363_cse,
      FpMul_8U_23U_lor_20_lpi_1_dfm_st, and_dcpl_104);
  assign nor_1471_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_4_lpi_1_dfm_st_6);
  assign nor_1472_nl = ~(mul_loop_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_4_lpi_1_dfm_st_6);
  assign mux_217_nl = MUX_s_1_2_2((nor_1472_nl), (nor_1471_nl), reg_FpMul_8U_23U_lor_6_lpi_1_dfm_4_cse);
  assign and_2246_nl = nor_64_cse & (mux_217_nl);
  assign nor_1473_nl = ~((~ mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_21_lpi_1_dfm_st | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_4_lpi_1_dfm_st_6);
  assign mux_218_nl = MUX_s_1_2_2((nor_1473_nl), (and_2246_nl), nor_53_cse);
  assign mux_219_nl = MUX_s_1_2_2(nor_177_cse, (mux_218_nl), or_309_cse);
  assign IsZero_8U_23U_aelse_and_35_cse = core_wen & (~ and_dcpl_50) & (mux_219_nl);
  assign mux_221_nl = MUX_s_1_2_2(or_2664_cse, or_tmp_287, mul_loop_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_222_nl = MUX_s_1_2_2((mux_221_nl), or_2664_cse, reg_FpMul_8U_23U_lor_6_lpi_1_dfm_4_cse);
  assign mux_223_nl = MUX_s_1_2_2(or_tmp_287, (mux_222_nl), nor_64_cse);
  assign mux_224_nl = MUX_s_1_2_2(or_2664_cse, or_tmp_287, or_378_cse);
  assign mux_225_nl = MUX_s_1_2_2((mux_224_nl), (mux_223_nl), nor_53_cse);
  assign or_382_nl = (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_4_lpi_1_dfm_st_7
      | ((IsNaN_8U_23U_land_4_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | (~
      IsNaN_8U_23U_1_land_4_lpi_1_dfm_8) | mul_loop_mul_if_land_4_lpi_1_dfm_9) &
      or_1253_cse);
  assign mux_226_nl = MUX_s_1_2_2((or_382_nl), (mux_225_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_57_cse = core_wen & (~ and_dcpl_50)
      & (~ (mux_226_nl));
  assign or_386_cse = mul_loop_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_6_lpi_1_dfm_4_cse;
  assign FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_28_cse = MUX_s_1_2_2(or_386_cse,
      FpMul_8U_23U_lor_21_lpi_1_dfm_st, and_dcpl_104);
  assign nor_1465_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_5_lpi_1_dfm_st_6);
  assign nor_1466_nl = ~(mul_loop_mul_5_FpMul_8U_23U_oelse_1_acc_itm_9_1 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_5_lpi_1_dfm_st_6);
  assign mux_231_nl = MUX_s_1_2_2((nor_1466_nl), (nor_1465_nl), reg_FpMul_8U_23U_lor_7_lpi_1_dfm_4_cse);
  assign and_2245_nl = nor_69_cse & (mux_231_nl);
  assign nor_1467_nl = ~((~ mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_22_lpi_1_dfm_st | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_5_lpi_1_dfm_st_6);
  assign mux_232_nl = MUX_s_1_2_2((nor_1467_nl), (and_2245_nl), nor_53_cse);
  assign mux_233_nl = MUX_s_1_2_2(nor_193_cse, (mux_232_nl), or_309_cse);
  assign IsZero_8U_23U_aelse_and_36_cse = core_wen & (~ and_dcpl_50) & (mux_233_nl);
  assign mux_235_nl = MUX_s_1_2_2(or_414_cse, or_tmp_310, mul_loop_mul_5_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_236_nl = MUX_s_1_2_2((mux_235_nl), or_414_cse, reg_FpMul_8U_23U_lor_7_lpi_1_dfm_4_cse);
  assign mux_237_nl = MUX_s_1_2_2(or_tmp_310, (mux_236_nl), nor_69_cse);
  assign mux_238_nl = MUX_s_1_2_2(or_414_cse, or_tmp_310, or_2675_cse);
  assign mux_239_nl = MUX_s_1_2_2((mux_238_nl), (mux_237_nl), nor_53_cse);
  assign or_405_nl = (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_5_lpi_1_dfm_st_7
      | ((IsNaN_8U_23U_land_5_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | (~
      IsNaN_8U_23U_1_land_5_lpi_1_dfm_8) | mul_loop_mul_if_land_5_lpi_1_dfm_9) &
      or_4387_cse);
  assign mux_240_nl = MUX_s_1_2_2((or_405_nl), (mux_239_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_60_cse = core_wen & (~ and_dcpl_50)
      & (~ (mux_240_nl));
  assign or_414_cse = mul_loop_mul_if_land_5_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_27_cse = MUX_s_1_2_2(FpMul_8U_23U_lor_22_lpi_1_dfm_mx0w0,
      FpMul_8U_23U_lor_22_lpi_1_dfm_st, and_dcpl_104);
  assign nor_1461_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_6_lpi_1_dfm_st_6);
  assign nor_1462_nl = ~(mul_loop_mul_6_FpMul_8U_23U_oelse_1_acc_itm_9_1 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_6_lpi_1_dfm_st_6);
  assign mux_246_nl = MUX_s_1_2_2((nor_1462_nl), (nor_1461_nl), reg_FpMul_8U_23U_lor_8_lpi_1_dfm_4_cse);
  assign and_2244_nl = nor_73_cse & (mux_246_nl);
  assign nor_1463_nl = ~((~ mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_23_lpi_1_dfm_st | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_6_lpi_1_dfm_st_6);
  assign mux_247_nl = MUX_s_1_2_2((nor_1463_nl), (and_2244_nl), nor_53_cse);
  assign mux_248_nl = MUX_s_1_2_2(nor_209_cse, (mux_247_nl), or_309_cse);
  assign IsZero_8U_23U_aelse_and_37_cse = core_wen & (~ and_dcpl_50) & (mux_248_nl);
  assign mux_250_nl = MUX_s_1_2_2(or_2698_cse, or_tmp_339, mul_loop_mul_6_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_251_nl = MUX_s_1_2_2((mux_250_nl), or_2698_cse, reg_FpMul_8U_23U_lor_8_lpi_1_dfm_4_cse);
  assign mux_252_nl = MUX_s_1_2_2(or_tmp_339, (mux_251_nl), nor_73_cse);
  assign mux_253_nl = MUX_s_1_2_2(or_2698_cse, or_tmp_339, or_430_cse);
  assign mux_254_nl = MUX_s_1_2_2((mux_253_nl), (mux_252_nl), nor_53_cse);
  assign or_434_nl = (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_6_lpi_1_dfm_st_7
      | ((IsNaN_8U_23U_land_6_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | (~
      IsNaN_8U_23U_1_land_6_lpi_1_dfm_8) | mul_loop_mul_if_land_6_lpi_1_dfm_9) &
      or_2342_cse);
  assign mux_255_nl = MUX_s_1_2_2((or_434_nl), (mux_254_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_63_cse = core_wen & (~ and_dcpl_50)
      & (~ (mux_255_nl));
  assign or_438_cse = mul_loop_mul_6_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_8_lpi_1_dfm_4_cse;
  assign FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_26_cse = MUX_s_1_2_2(or_438_cse,
      FpMul_8U_23U_lor_23_lpi_1_dfm_st, and_dcpl_104);
  assign nor_1455_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_7_lpi_1_dfm_st_6);
  assign nor_1456_nl = ~(mul_loop_mul_7_FpMul_8U_23U_oelse_1_acc_itm_9_1 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_7_lpi_1_dfm_st_6);
  assign mux_260_nl = MUX_s_1_2_2((nor_1456_nl), (nor_1455_nl), reg_FpMul_8U_23U_lor_9_lpi_1_dfm_4_cse);
  assign and_2243_nl = nor_78_cse & (mux_260_nl);
  assign nor_1457_nl = ~((~ mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_24_lpi_1_dfm_st | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_7_lpi_1_dfm_st_6);
  assign mux_261_nl = MUX_s_1_2_2((nor_1457_nl), (and_2243_nl), nor_53_cse);
  assign mux_262_nl = MUX_s_1_2_2(nor_225_cse, (mux_261_nl), or_309_cse);
  assign IsZero_8U_23U_aelse_and_38_cse = core_wen & (~ and_dcpl_50) & (mux_262_nl);
  assign mux_264_nl = MUX_s_1_2_2(or_2711_cse, or_tmp_362, mul_loop_mul_7_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_265_nl = MUX_s_1_2_2((mux_264_nl), or_2711_cse, reg_FpMul_8U_23U_lor_9_lpi_1_dfm_4_cse);
  assign mux_266_nl = MUX_s_1_2_2(or_tmp_362, (mux_265_nl), nor_78_cse);
  assign mux_267_nl = MUX_s_1_2_2(or_2711_cse, or_tmp_362, or_453_cse);
  assign mux_268_nl = MUX_s_1_2_2((mux_267_nl), (mux_266_nl), nor_53_cse);
  assign or_457_nl = (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_7_lpi_1_dfm_st_7
      | ((IsNaN_8U_23U_land_7_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | (~
      IsNaN_8U_23U_1_land_7_lpi_1_dfm_8) | mul_loop_mul_if_land_7_lpi_1_dfm_9) &
      or_4389_cse);
  assign mux_269_nl = MUX_s_1_2_2((or_457_nl), (mux_268_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_66_cse = core_wen & (~ and_dcpl_50)
      & (~ (mux_269_nl));
  assign or_461_cse = mul_loop_mul_7_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_9_lpi_1_dfm_4_cse;
  assign FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_25_cse = MUX_s_1_2_2(or_461_cse,
      FpMul_8U_23U_lor_24_lpi_1_dfm_st, and_dcpl_104);
  assign nor_1449_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_8_lpi_1_dfm_st_6);
  assign nor_1450_nl = ~(mul_loop_mul_8_FpMul_8U_23U_oelse_1_acc_itm_9_1 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_8_lpi_1_dfm_st_6);
  assign mux_274_nl = MUX_s_1_2_2((nor_1450_nl), (nor_1449_nl), reg_FpMul_8U_23U_lor_10_lpi_1_dfm_4_cse);
  assign and_2242_nl = nor_83_cse & (mux_274_nl);
  assign nor_1451_nl = ~((~ mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_25_lpi_1_dfm_st | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_8_lpi_1_dfm_st_6);
  assign mux_275_nl = MUX_s_1_2_2((nor_1451_nl), (and_2242_nl), nor_53_cse);
  assign mux_276_nl = MUX_s_1_2_2(nor_241_cse, (mux_275_nl), or_309_cse);
  assign IsZero_8U_23U_aelse_and_39_cse = core_wen & (~ and_dcpl_50) & (mux_276_nl);
  assign mux_278_nl = MUX_s_1_2_2(or_2721_cse, or_tmp_385, mul_loop_mul_8_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_279_nl = MUX_s_1_2_2((mux_278_nl), or_2721_cse, reg_FpMul_8U_23U_lor_10_lpi_1_dfm_4_cse);
  assign mux_280_nl = MUX_s_1_2_2(or_tmp_385, (mux_279_nl), nor_83_cse);
  assign mux_281_nl = MUX_s_1_2_2(or_2721_cse, or_tmp_385, or_2722_cse);
  assign mux_282_nl = MUX_s_1_2_2((mux_281_nl), (mux_280_nl), nor_53_cse);
  assign or_480_nl = (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_8_lpi_1_dfm_st_7
      | ((IsNaN_8U_23U_land_8_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | (~
      IsNaN_8U_23U_1_land_8_lpi_1_dfm_8) | mul_loop_mul_if_land_8_lpi_1_dfm_9) &
      or_4390_cse);
  assign mux_283_nl = MUX_s_1_2_2((or_480_nl), (mux_282_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_69_cse = core_wen & (~ and_dcpl_50)
      & (~ (mux_283_nl));
  assign FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_24_cse = MUX_s_1_2_2(or_2742_cse,
      FpMul_8U_23U_lor_25_lpi_1_dfm_st, and_dcpl_104);
  assign nor_1445_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_9_lpi_1_dfm_st_6);
  assign nor_1446_nl = ~(mul_loop_mul_9_FpMul_8U_23U_oelse_1_acc_itm_9_1 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_9_lpi_1_dfm_st_6);
  assign mux_289_nl = MUX_s_1_2_2((nor_1446_nl), (nor_1445_nl), reg_FpMul_8U_23U_lor_11_lpi_1_dfm_4_cse);
  assign and_2241_nl = nor_87_cse & (mux_289_nl);
  assign nor_1447_nl = ~((~ mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_26_lpi_1_dfm_st | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_9_lpi_1_dfm_st_6);
  assign mux_290_nl = MUX_s_1_2_2((nor_1447_nl), (and_2241_nl), nor_53_cse);
  assign mux_291_nl = MUX_s_1_2_2(nor_257_cse, (mux_290_nl), or_309_cse);
  assign IsZero_8U_23U_aelse_and_40_cse = core_wen & (~ and_dcpl_50) & (mux_291_nl);
  assign mux_293_nl = MUX_s_1_2_2(or_517_cse, or_tmp_413, mul_loop_mul_9_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_294_nl = MUX_s_1_2_2((mux_293_nl), or_517_cse, reg_FpMul_8U_23U_lor_11_lpi_1_dfm_4_cse);
  assign mux_295_nl = MUX_s_1_2_2(or_tmp_413, (mux_294_nl), nor_87_cse);
  assign mux_296_nl = MUX_s_1_2_2(or_517_cse, or_tmp_413, or_2745_cse);
  assign mux_297_nl = MUX_s_1_2_2((mux_296_nl), (mux_295_nl), nor_53_cse);
  assign or_508_nl = (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_9_lpi_1_dfm_st_7
      | ((IsNaN_8U_23U_land_9_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | (~
      IsNaN_8U_23U_1_land_9_lpi_1_dfm_8) | mul_loop_mul_if_land_9_lpi_1_dfm_9) &
      or_4391_cse);
  assign mux_298_nl = MUX_s_1_2_2((or_508_nl), (mux_297_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_72_cse = core_wen & (~ and_dcpl_50)
      & (~ (mux_298_nl));
  assign or_517_cse = mul_loop_mul_if_land_9_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_23_cse = MUX_s_1_2_2(FpMul_8U_23U_lor_26_lpi_1_dfm_mx0w0,
      FpMul_8U_23U_lor_26_lpi_1_dfm_st, and_dcpl_104);
  assign nor_1441_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_10_lpi_1_dfm_st_6);
  assign nor_1442_nl = ~(mul_loop_mul_10_FpMul_8U_23U_oelse_1_acc_itm_9_1 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_10_lpi_1_dfm_st_6);
  assign mux_304_nl = MUX_s_1_2_2((nor_1442_nl), (nor_1441_nl), reg_FpMul_8U_23U_lor_12_lpi_1_dfm_4_cse);
  assign and_2240_nl = nor_91_cse & (mux_304_nl);
  assign nor_1443_nl = ~((~ mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_27_lpi_1_dfm_st | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_10_lpi_1_dfm_st_6);
  assign mux_305_nl = MUX_s_1_2_2((nor_1443_nl), (and_2240_nl), nor_53_cse);
  assign mux_306_nl = MUX_s_1_2_2(nor_273_cse, (mux_305_nl), or_309_cse);
  assign IsZero_8U_23U_aelse_and_41_cse = core_wen & (~ and_dcpl_50) & (mux_306_nl);
  assign mux_308_nl = MUX_s_1_2_2(or_2767_cse, or_tmp_442, mul_loop_mul_10_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_309_nl = MUX_s_1_2_2((mux_308_nl), or_2767_cse, reg_FpMul_8U_23U_lor_12_lpi_1_dfm_4_cse);
  assign mux_310_nl = MUX_s_1_2_2(or_tmp_442, (mux_309_nl), nor_91_cse);
  assign mux_311_nl = MUX_s_1_2_2(or_2767_cse, or_tmp_442, or_533_cse);
  assign mux_312_nl = MUX_s_1_2_2((mux_311_nl), (mux_310_nl), nor_53_cse);
  assign or_537_nl = (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_10_lpi_1_dfm_st_7
      | ((IsNaN_8U_23U_land_10_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 |
      (~ IsNaN_8U_23U_1_land_10_lpi_1_dfm_8) | mul_loop_mul_if_land_10_lpi_1_dfm_9)
      & or_2386_cse);
  assign mux_313_nl = MUX_s_1_2_2((or_537_nl), (mux_312_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_75_cse = core_wen & (~ and_dcpl_50)
      & (~ (mux_313_nl));
  assign FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_22_cse = MUX_s_1_2_2(FpMul_8U_23U_lor_27_lpi_1_dfm_mx0w0,
      FpMul_8U_23U_lor_27_lpi_1_dfm_st, and_dcpl_104);
  assign nor_1437_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_11_lpi_1_dfm_st_6);
  assign nor_1438_nl = ~(mul_loop_mul_11_FpMul_8U_23U_oelse_1_acc_itm_9_1 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_11_lpi_1_dfm_st_6);
  assign mux_319_nl = MUX_s_1_2_2((nor_1438_nl), (nor_1437_nl), reg_FpMul_8U_23U_lor_13_lpi_1_dfm_4_cse);
  assign and_2239_nl = nor_95_cse & (mux_319_nl);
  assign nor_1439_nl = ~((~ mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_28_lpi_1_dfm_st | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_11_lpi_1_dfm_st_6);
  assign mux_320_nl = MUX_s_1_2_2((nor_1439_nl), (and_2239_nl), nor_53_cse);
  assign mux_321_nl = MUX_s_1_2_2(nor_289_cse, (mux_320_nl), or_309_cse);
  assign IsZero_8U_23U_aelse_and_42_cse = core_wen & (~ and_dcpl_50) & (mux_321_nl);
  assign mux_323_nl = MUX_s_1_2_2(or_2774_cse, or_tmp_471, mul_loop_mul_11_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_324_nl = MUX_s_1_2_2((mux_323_nl), or_2774_cse, reg_FpMul_8U_23U_lor_13_lpi_1_dfm_4_cse);
  assign mux_325_nl = MUX_s_1_2_2(or_tmp_471, (mux_324_nl), nor_95_cse);
  assign mux_326_nl = MUX_s_1_2_2(or_2774_cse, or_tmp_471, or_562_cse);
  assign mux_327_nl = MUX_s_1_2_2((mux_326_nl), (mux_325_nl), nor_53_cse);
  assign or_566_nl = (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_11_lpi_1_dfm_st_7
      | ((IsNaN_8U_23U_land_11_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 |
      (~ IsNaN_8U_23U_1_land_11_lpi_1_dfm_8) | mul_loop_mul_if_land_11_lpi_1_dfm_9)
      & or_1819_cse);
  assign mux_328_nl = MUX_s_1_2_2((or_566_nl), (mux_327_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_78_cse = core_wen & (~ and_dcpl_50)
      & (~ (mux_328_nl));
  assign or_570_cse = mul_loop_mul_11_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_13_lpi_1_dfm_4_cse;
  assign FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_21_cse = MUX_s_1_2_2(or_570_cse,
      FpMul_8U_23U_lor_28_lpi_1_dfm_st, and_dcpl_104);
  assign nor_1431_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_12_lpi_1_dfm_st_6);
  assign nor_1432_nl = ~(mul_loop_mul_12_FpMul_8U_23U_oelse_1_acc_itm_9_1 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_12_lpi_1_dfm_st_6);
  assign mux_333_nl = MUX_s_1_2_2((nor_1432_nl), (nor_1431_nl), reg_FpMul_8U_23U_lor_14_lpi_1_dfm_4_cse);
  assign and_2238_nl = nor_100_cse & (mux_333_nl);
  assign nor_1433_nl = ~((~ mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_29_lpi_1_dfm_st | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_12_lpi_1_dfm_st_6);
  assign mux_334_nl = MUX_s_1_2_2((nor_1433_nl), (and_2238_nl), nor_53_cse);
  assign mux_335_nl = MUX_s_1_2_2(nor_305_cse, (mux_334_nl), or_309_cse);
  assign IsZero_8U_23U_aelse_and_43_cse = core_wen & (~ and_dcpl_50) & (mux_335_nl);
  assign mux_337_nl = MUX_s_1_2_2(or_2787_cse, or_tmp_494, mul_loop_mul_12_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_338_nl = MUX_s_1_2_2((mux_337_nl), or_2787_cse, reg_FpMul_8U_23U_lor_14_lpi_1_dfm_4_cse);
  assign mux_339_nl = MUX_s_1_2_2(or_tmp_494, (mux_338_nl), nor_100_cse);
  assign mux_340_nl = MUX_s_1_2_2(or_2787_cse, or_tmp_494, or_585_cse);
  assign mux_341_nl = MUX_s_1_2_2((mux_340_nl), (mux_339_nl), nor_53_cse);
  assign or_589_nl = (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_12_lpi_1_dfm_st_7
      | ((IsNaN_8U_23U_land_12_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 |
      (~ IsNaN_8U_23U_1_land_12_lpi_1_dfm_8) | mul_loop_mul_if_land_12_lpi_1_dfm_9)
      & or_1898_cse);
  assign mux_342_nl = MUX_s_1_2_2((or_589_nl), (mux_341_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_81_cse = core_wen & (~ and_dcpl_50)
      & (~ (mux_342_nl));
  assign or_593_cse = mul_loop_mul_12_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_14_lpi_1_dfm_4_cse;
  assign FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_20_cse = MUX_s_1_2_2(or_593_cse,
      FpMul_8U_23U_lor_29_lpi_1_dfm_st, and_dcpl_104);
  assign nor_1425_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_13_lpi_1_dfm_st_6);
  assign nor_1426_nl = ~(mul_loop_mul_13_FpMul_8U_23U_oelse_1_acc_itm_9_1 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_13_lpi_1_dfm_st_6);
  assign mux_347_nl = MUX_s_1_2_2((nor_1426_nl), (nor_1425_nl), reg_FpMul_8U_23U_lor_15_lpi_1_dfm_4_cse);
  assign and_2237_nl = nor_105_cse & (mux_347_nl);
  assign nor_1427_nl = ~((~ mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_30_lpi_1_dfm_st | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_13_lpi_1_dfm_st_6);
  assign mux_348_nl = MUX_s_1_2_2((nor_1427_nl), (and_2237_nl), nor_53_cse);
  assign mux_349_nl = MUX_s_1_2_2(nor_321_cse, (mux_348_nl), or_309_cse);
  assign IsZero_8U_23U_aelse_and_44_cse = core_wen & (~ and_dcpl_50) & (mux_349_nl);
  assign mux_351_nl = MUX_s_1_2_2(or_2797_cse, or_tmp_517, mul_loop_mul_13_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_352_nl = MUX_s_1_2_2((mux_351_nl), or_2797_cse, reg_FpMul_8U_23U_lor_15_lpi_1_dfm_4_cse);
  assign mux_353_nl = MUX_s_1_2_2(or_tmp_517, (mux_352_nl), nor_105_cse);
  assign mux_354_nl = MUX_s_1_2_2(or_2797_cse, or_tmp_517, or_2798_cse);
  assign mux_355_nl = MUX_s_1_2_2((mux_354_nl), (mux_353_nl), nor_53_cse);
  assign or_612_nl = (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_13_lpi_1_dfm_st_7
      | ((IsNaN_8U_23U_land_13_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 |
      (~ IsNaN_8U_23U_1_land_13_lpi_1_dfm_8) | mul_loop_mul_if_land_13_lpi_1_dfm_9)
      & or_1981_cse);
  assign mux_356_nl = MUX_s_1_2_2((or_612_nl), (mux_355_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_84_cse = core_wen & (~ and_dcpl_50)
      & (~ (mux_356_nl));
  assign or_616_cse = mul_loop_mul_13_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_15_lpi_1_dfm_4_cse;
  assign FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_19_cse = MUX_s_1_2_2(or_616_cse,
      FpMul_8U_23U_lor_30_lpi_1_dfm_st, and_dcpl_104);
  assign nor_1419_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_14_lpi_1_dfm_st_6);
  assign nor_1420_nl = ~(mul_loop_mul_14_FpMul_8U_23U_oelse_1_acc_itm_9_1 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_14_lpi_1_dfm_st_6);
  assign mux_361_nl = MUX_s_1_2_2((nor_1420_nl), (nor_1419_nl), reg_FpMul_8U_23U_lor_16_lpi_1_dfm_4_cse);
  assign and_2236_nl = nor_110_cse & (mux_361_nl);
  assign nor_1421_nl = ~((~ mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_31_lpi_1_dfm_st | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_14_lpi_1_dfm_st_6);
  assign mux_362_nl = MUX_s_1_2_2((nor_1421_nl), (and_2236_nl), nor_53_cse);
  assign mux_363_nl = MUX_s_1_2_2(nor_336_cse, (mux_362_nl), or_309_cse);
  assign IsZero_8U_23U_aelse_and_45_cse = core_wen & (~ and_dcpl_50) & (mux_363_nl);
  assign mux_365_nl = MUX_s_1_2_2(or_2823_cse, or_tmp_540, mul_loop_mul_14_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_366_nl = MUX_s_1_2_2((mux_365_nl), or_2823_cse, reg_FpMul_8U_23U_lor_16_lpi_1_dfm_4_cse);
  assign mux_367_nl = MUX_s_1_2_2(or_tmp_540, (mux_366_nl), nor_110_cse);
  assign mux_368_nl = MUX_s_1_2_2(or_2823_cse, or_tmp_540, or_631_cse);
  assign mux_369_nl = MUX_s_1_2_2((mux_368_nl), (mux_367_nl), nor_53_cse);
  assign or_635_nl = (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_14_lpi_1_dfm_st_7
      | ((IsNaN_8U_23U_land_14_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 |
      (~ IsNaN_8U_23U_1_land_14_lpi_1_dfm_8) | mul_loop_mul_if_land_14_lpi_1_dfm_9)
      & or_4398_cse);
  assign mux_370_nl = MUX_s_1_2_2((or_635_nl), (mux_369_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_87_cse = core_wen & (~ and_dcpl_50)
      & (~ (mux_370_nl));
  assign or_639_cse = mul_loop_mul_14_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_16_lpi_1_dfm_4_cse;
  assign FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_18_cse = MUX_s_1_2_2(or_639_cse,
      FpMul_8U_23U_lor_31_lpi_1_dfm_st, and_dcpl_104);
  assign nor_1413_cse = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_15_lpi_1_dfm_st_6);
  assign nor_1414_nl = ~(mul_loop_mul_15_FpMul_8U_23U_oelse_1_acc_itm_9_1 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_15_lpi_1_dfm_st_6);
  assign mux_375_nl = MUX_s_1_2_2((nor_1414_nl), nor_1413_cse, reg_FpMul_8U_23U_lor_17_lpi_1_dfm_4_cse);
  assign and_2235_nl = nor_115_cse & (mux_375_nl);
  assign nor_1415_nl = ~((~ mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_32_lpi_1_dfm_st | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_15_lpi_1_dfm_st_6);
  assign mux_376_nl = MUX_s_1_2_2((nor_1415_nl), (and_2235_nl), nor_53_cse);
  assign mux_377_nl = MUX_s_1_2_2(nor_352_cse, (mux_376_nl), or_309_cse);
  assign IsZero_8U_23U_aelse_and_46_cse = core_wen & (~ and_dcpl_50) & (mux_377_nl);
  assign mux_379_nl = MUX_s_1_2_2(or_2833_cse, or_tmp_563, mul_loop_mul_15_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_380_nl = MUX_s_1_2_2((mux_379_nl), or_2833_cse, reg_FpMul_8U_23U_lor_17_lpi_1_dfm_4_cse);
  assign mux_381_nl = MUX_s_1_2_2(or_tmp_563, (mux_380_nl), nor_115_cse);
  assign mux_382_nl = MUX_s_1_2_2(or_2833_cse, or_tmp_563, or_2834_cse);
  assign mux_383_nl = MUX_s_1_2_2((mux_382_nl), (mux_381_nl), nor_53_cse);
  assign or_658_nl = (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_15_lpi_1_dfm_st_7
      | ((IsNaN_8U_23U_land_15_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 |
      (~ IsNaN_8U_23U_1_land_15_lpi_1_dfm_8) | mul_loop_mul_if_land_15_lpi_1_dfm_9)
      & or_4399_cse);
  assign mux_384_nl = MUX_s_1_2_2((or_658_nl), (mux_383_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_90_cse = core_wen & (~ and_dcpl_50)
      & (~ (mux_384_nl));
  assign or_662_cse = mul_loop_mul_15_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_17_lpi_1_dfm_4_cse;
  assign FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_17_cse = MUX_s_1_2_2(or_662_cse,
      FpMul_8U_23U_lor_32_lpi_1_dfm_st, and_dcpl_104);
  assign nor_1407_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_lpi_1_dfm_st_6);
  assign nor_1408_nl = ~(mul_loop_mul_16_FpMul_8U_23U_oelse_1_acc_itm_9_1 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_lpi_1_dfm_st_6);
  assign mux_389_nl = MUX_s_1_2_2((nor_1408_nl), (nor_1407_nl), reg_FpMul_8U_23U_lor_lpi_1_dfm_4_cse);
  assign and_2234_nl = nor_120_cse & (mux_389_nl);
  assign nor_1409_nl = ~((~ mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_1_lpi_1_dfm_st | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_lpi_1_dfm_st_6);
  assign mux_390_nl = MUX_s_1_2_2((nor_1409_nl), (and_2234_nl), nor_53_cse);
  assign mux_391_nl = MUX_s_1_2_2(nor_368_cse, (mux_390_nl), or_309_cse);
  assign IsZero_8U_23U_aelse_and_47_cse = core_wen & (~ and_dcpl_50) & (mux_391_nl);
  assign mux_393_nl = MUX_s_1_2_2(or_2864_cse, or_tmp_586, mul_loop_mul_16_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_394_nl = MUX_s_1_2_2((mux_393_nl), or_2864_cse, reg_FpMul_8U_23U_lor_lpi_1_dfm_4_cse);
  assign mux_395_nl = MUX_s_1_2_2(or_tmp_586, (mux_394_nl), nor_120_cse);
  assign mux_396_nl = MUX_s_1_2_2(or_2864_cse, or_tmp_586, or_2865_cse);
  assign mux_397_nl = MUX_s_1_2_2((mux_396_nl), (mux_395_nl), nor_53_cse);
  assign or_681_nl = (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_lpi_1_dfm_st_7
      | ((IsNaN_8U_23U_land_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | (~
      IsNaN_8U_23U_1_land_lpi_1_dfm_8) | mul_loop_mul_if_land_lpi_1_dfm_9) & or_4400_cse);
  assign mux_398_nl = MUX_s_1_2_2((or_681_nl), (mux_397_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_93_cse = core_wen & (~ and_dcpl_50)
      & (~ (mux_398_nl));
  assign FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_16_cse = MUX_s_1_2_2(or_2885_cse,
      FpMul_8U_23U_lor_1_lpi_1_dfm_st, and_dcpl_104);
  assign mux_404_nl = MUX_s_1_2_2(or_tmp_608, or_tmp_204, or_309_cse);
  assign mul_loop_mul_if_aelse_and_48_cse = core_wen & (~ and_dcpl_50) & (~ (mux_404_nl));
  assign mux_405_nl = MUX_s_1_2_2(main_stage_v_4, main_stage_v_3, or_309_cse);
  assign MulIn_data_and_2_cse = core_wen & (~ and_dcpl_50) & (mux_405_nl);
  assign and_718_nl = and_dcpl_172 & and_dcpl_85;
  assign and_719_nl = and_dcpl_172 & or_90_cse;
  assign mux_1616_nl = MUX_s_1_2_2(IsNaN_8U_23U_1_land_1_lpi_1_dfm_9, IsNaN_8U_23U_1_land_1_lpi_1_dfm_8,
      or_309_cse);
  assign FpMul_8U_23U_p_expo_mux1h_1_itm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_1_sva_1_mx0w0,
      FpMul_8U_23U_p_expo_1_sva_1, ({4'b0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_10}),
      {(and_718_nl) , (and_719_nl) , (mux_1616_nl)});
  assign or_cse = (~ (mul_loop_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) | mul_loop_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  assign or_4735_nl = (or_cse & mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2)
      | FpMul_8U_23U_lor_18_lpi_1_dfm_6;
  assign and_2512_nl = FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_2
      & mul_loop_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
      & or_tmp_893;
  assign mux_1689_nl = MUX_s_1_2_2((and_2512_nl), or_tmp_893, FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm);
  assign mux_1690_cse = MUX_s_1_2_2((mux_1689_nl), (or_4735_nl), nor_53_cse);
  assign nor_129_cse = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_1_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_18_lpi_1_dfm_st_3
      | (~ mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1387_nl = ~(IsNaN_8U_23U_land_1_lpi_1_dfm_st_7 | (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_1_lpi_1_dfm_10 | mul_loop_mul_if_land_1_lpi_1_dfm_st_7
      | mul_loop_mul_if_land_1_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign nor_1388_nl = ~((~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_9) | IsNaN_8U_23U_land_1_lpi_1_dfm_st_8
      | IsNaN_8U_23U_land_1_lpi_1_dfm_11 | mul_loop_mul_if_land_1_lpi_1_dfm_st_8
      | mul_loop_mul_if_land_1_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4));
  assign mux_516_nl = MUX_s_1_2_2((nor_1388_nl), (nor_1387_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_96_cse = core_wen & (~ and_dcpl_50)
      & (mux_516_nl);
  assign nor_133_cse = ~(FpMul_8U_23U_lor_18_lpi_1_dfm_st_3 | (~ mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1383_cse = ~((~ (mul_loop_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7);
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_31_cse = MUX_s_1_2_2(mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs_mx0w0,
      mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs, and_dcpl_104);
  assign nor_1379_nl = ~((~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_8) | IsNaN_8U_23U_land_1_lpi_1_dfm_10
      | mul_loop_mul_if_land_1_lpi_1_dfm_st_7 | mul_loop_mul_if_land_1_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3));
  assign nor_1380_nl = ~((~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_9) | IsNaN_8U_23U_land_1_lpi_1_dfm_11
      | mul_loop_mul_if_land_1_lpi_1_dfm_st_8 | mul_loop_mul_if_land_1_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4));
  assign mux_521_nl = MUX_s_1_2_2((nor_1380_nl), (nor_1379_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_96_cse = core_wen & (~ and_dcpl_50)
      & (mux_521_nl);
  assign IsNaN_8U_23U_aelse_and_48_cse = core_wen & (~ and_dcpl_50) & (~ mux_522_itm);
  assign nor_1373_nl = ~(nor_1383_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_1_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_1_lpi_1_dfm_10
      | FpMul_8U_23U_lor_18_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8
      | mul_loop_mul_if_land_1_lpi_1_dfm_9);
  assign nor_1375_nl = ~((FpMul_8U_23U_p_mant_p1_1_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_1_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_1_lpi_1_dfm_10 | FpMul_8U_23U_lor_18_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 | mul_loop_mul_if_land_1_lpi_1_dfm_9);
  assign mux_524_nl = MUX_s_1_2_2((nor_1375_nl), (nor_1373_nl), nor_133_cse);
  assign and_2228_nl = mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_524_nl);
  assign nor_1376_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_1_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_1_lpi_1_dfm_10 | FpMul_8U_23U_lor_18_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 | mul_loop_mul_if_land_1_lpi_1_dfm_9);
  assign mux_525_nl = MUX_s_1_2_2((nor_1376_nl), (and_2228_nl), nor_53_cse);
  assign nor_1377_nl = ~((~((~ mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs_2) |
      mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs_st_2)) | (~ main_stage_v_4) |
      IsNaN_8U_23U_land_1_lpi_1_dfm_11 | mul_loop_mul_if_land_1_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_1_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_1_lpi_1_dfm_9 | FpMul_8U_23U_lor_18_lpi_1_dfm_7 | (~
      FpMul_8U_23U_FpMul_8U_23U_and_itm_2));
  assign mux_526_nl = MUX_s_1_2_2((nor_1377_nl), (mux_525_nl), or_309_cse);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_cse = core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse
      & (mux_526_nl);
  assign and_723_nl = and_dcpl_177 & and_dcpl_85;
  assign and_724_nl = and_dcpl_177 & or_90_cse;
  assign mux_1617_nl = MUX_s_1_2_2(IsNaN_8U_23U_1_land_2_lpi_1_dfm_9, IsNaN_8U_23U_1_land_2_lpi_1_dfm_8,
      or_309_cse);
  assign FpMul_8U_23U_p_expo_mux1h_3_itm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_2_sva_1_mx0w0,
      FpMul_8U_23U_p_expo_2_sva_1, ({4'b0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_10}),
      {(and_723_nl) , (and_724_nl) , (mux_1617_nl)});
  assign or_4962_cse = (~ (mul_loop_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) |
      mul_loop_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  assign or_4747_nl = (or_4962_cse & mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2)
      | FpMul_8U_23U_lor_19_lpi_1_dfm_6;
  assign and_2534_nl = FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_2
      & mul_loop_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
      & or_tmp_975;
  assign mux_1694_nl = MUX_s_1_2_2((and_2534_nl), or_tmp_975, FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm);
  assign mux_1695_cse = MUX_s_1_2_2((mux_1694_nl), (or_4747_nl), nor_53_cse);
  assign nor_145_cse = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_2_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_19_lpi_1_dfm_st_3
      | (~ mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1355_nl = ~(IsNaN_8U_23U_land_2_lpi_1_dfm_st_7 | (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_2_lpi_1_dfm_10 | mul_loop_mul_if_land_2_lpi_1_dfm_st_7
      | mul_loop_mul_if_land_2_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign nor_1356_nl = ~((~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_9) | IsNaN_8U_23U_land_2_lpi_1_dfm_st_8
      | IsNaN_8U_23U_land_2_lpi_1_dfm_11 | mul_loop_mul_if_land_2_lpi_1_dfm_st_8
      | mul_loop_mul_if_land_2_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4));
  assign mux_540_nl = MUX_s_1_2_2((nor_1356_nl), (nor_1355_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_98_cse = core_wen & (~ and_dcpl_50)
      & (mux_540_nl);
  assign nor_149_cse = ~(FpMul_8U_23U_lor_19_lpi_1_dfm_st_3 | (~ mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1351_cse = ~((~ (mul_loop_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7);
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_29_cse = MUX_s_1_2_2(mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs_mx0w0,
      mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs, and_dcpl_104);
  assign nor_1347_nl = ~((~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_8) | IsNaN_8U_23U_land_2_lpi_1_dfm_10
      | mul_loop_mul_if_land_2_lpi_1_dfm_st_7 | mul_loop_mul_if_land_2_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3));
  assign nor_1348_nl = ~((~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_9) | IsNaN_8U_23U_land_2_lpi_1_dfm_11
      | mul_loop_mul_if_land_2_lpi_1_dfm_st_8 | mul_loop_mul_if_land_2_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4));
  assign mux_545_nl = MUX_s_1_2_2((nor_1348_nl), (nor_1347_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_99_cse = core_wen & (~ and_dcpl_50)
      & (mux_545_nl);
  assign IsNaN_8U_23U_aelse_and_50_cse = core_wen & (~ and_dcpl_50) & (~ mux_546_itm);
  assign nor_1341_nl = ~(nor_1351_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_2_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_2_lpi_1_dfm_10
      | FpMul_8U_23U_lor_19_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_2_lpi_1_dfm_8
      | mul_loop_mul_if_land_2_lpi_1_dfm_9);
  assign nor_1343_nl = ~((FpMul_8U_23U_p_mant_p1_2_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_2_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_2_lpi_1_dfm_10 | FpMul_8U_23U_lor_19_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 | mul_loop_mul_if_land_2_lpi_1_dfm_9);
  assign mux_548_nl = MUX_s_1_2_2((nor_1343_nl), (nor_1341_nl), nor_149_cse);
  assign and_2222_nl = mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_548_nl);
  assign nor_1344_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_64_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_2_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_2_lpi_1_dfm_10 | FpMul_8U_23U_lor_19_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 | mul_loop_mul_if_land_2_lpi_1_dfm_9);
  assign mux_549_nl = MUX_s_1_2_2((nor_1344_nl), (and_2222_nl), nor_53_cse);
  assign nor_1345_nl = ~((~((~ mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs_2) |
      mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs_st_2)) | (~ main_stage_v_4) |
      io_read_cfg_mul_bypass_rsc_svs_8 | IsNaN_8U_23U_land_2_lpi_1_dfm_11 | mul_loop_mul_if_land_2_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_2_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_2_lpi_1_dfm_9 | FpMul_8U_23U_lor_19_lpi_1_dfm_7 | (~
      FpMul_8U_23U_FpMul_8U_23U_and_64_itm_2));
  assign mux_550_nl = MUX_s_1_2_2((nor_1345_nl), (mux_549_nl), or_309_cse);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_1_cse = core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse
      & (mux_550_nl);
  assign and_728_nl = and_dcpl_182 & and_dcpl_85;
  assign and_729_nl = and_dcpl_182 & or_90_cse;
  assign mux_1618_nl = MUX_s_1_2_2(IsNaN_8U_23U_1_land_3_lpi_1_dfm_9, IsNaN_8U_23U_1_land_3_lpi_1_dfm_8,
      or_309_cse);
  assign FpMul_8U_23U_p_expo_mux1h_5_itm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_3_sva_1_mx0w0,
      FpMul_8U_23U_p_expo_3_sva_1, ({4'b0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_10}),
      {(and_728_nl) , (and_729_nl) , (mux_1618_nl)});
  assign or_4959_cse = (~ (mul_loop_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) |
      mul_loop_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  assign or_4759_nl = (or_4959_cse & mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2)
      | FpMul_8U_23U_lor_20_lpi_1_dfm_6;
  assign and_2556_nl = FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_2
      & mul_loop_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
      & or_tmp_1055;
  assign mux_1699_nl = MUX_s_1_2_2((and_2556_nl), or_tmp_1055, FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm);
  assign mux_1700_cse = MUX_s_1_2_2((mux_1699_nl), (or_4759_nl), nor_53_cse);
  assign nor_161_cse = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_3_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_20_lpi_1_dfm_st_3
      | (~ mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1321_nl = ~(IsNaN_8U_23U_land_3_lpi_1_dfm_st_7 | (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_3_lpi_1_dfm_10 | mul_loop_mul_if_land_3_lpi_1_dfm_st_7
      | mul_loop_mul_if_land_3_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign nor_1322_nl = ~(IsNaN_8U_23U_land_3_lpi_1_dfm_st_8 | (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_9)
      | IsNaN_8U_23U_land_3_lpi_1_dfm_11 | mul_loop_mul_if_land_3_lpi_1_dfm_st_8
      | mul_loop_mul_if_land_3_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4));
  assign mux_564_nl = MUX_s_1_2_2((nor_1322_nl), (nor_1321_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_100_cse = core_wen & (~ and_dcpl_50)
      & (mux_564_nl);
  assign nor_165_cse = ~(FpMul_8U_23U_lor_20_lpi_1_dfm_st_3 | (~ mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1317_cse = ~((~ (mul_loop_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7);
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_27_cse = MUX_s_1_2_2(mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs_mx0w0,
      mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs, and_dcpl_104);
  assign nor_1313_nl = ~((~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_8) | IsNaN_8U_23U_land_3_lpi_1_dfm_10
      | mul_loop_mul_if_land_3_lpi_1_dfm_st_7 | mul_loop_mul_if_land_3_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3));
  assign nor_1314_nl = ~((~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_9) | IsNaN_8U_23U_land_3_lpi_1_dfm_11
      | mul_loop_mul_if_land_3_lpi_1_dfm_st_8 | mul_loop_mul_if_land_3_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4));
  assign mux_569_nl = MUX_s_1_2_2((nor_1314_nl), (nor_1313_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_102_cse = core_wen & (~ and_dcpl_50)
      & (mux_569_nl);
  assign IsNaN_8U_23U_aelse_and_52_cse = core_wen & (~ and_dcpl_50) & (~ mux_570_itm);
  assign nor_1307_nl = ~(nor_1317_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_3_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_3_lpi_1_dfm_10
      | FpMul_8U_23U_lor_20_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_3_lpi_1_dfm_8
      | mul_loop_mul_if_land_3_lpi_1_dfm_9);
  assign nor_1309_nl = ~((FpMul_8U_23U_p_mant_p1_3_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_3_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_3_lpi_1_dfm_10 | FpMul_8U_23U_lor_20_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 | mul_loop_mul_if_land_3_lpi_1_dfm_9);
  assign mux_572_nl = MUX_s_1_2_2((nor_1309_nl), (nor_1307_nl), nor_165_cse);
  assign and_2216_nl = mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_572_nl);
  assign nor_1310_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_65_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_3_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_3_lpi_1_dfm_10 | FpMul_8U_23U_lor_20_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 | mul_loop_mul_if_land_3_lpi_1_dfm_9);
  assign mux_573_nl = MUX_s_1_2_2((nor_1310_nl), (and_2216_nl), nor_53_cse);
  assign nor_1311_nl = ~((~((~ mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs_2) |
      mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs_st_2)) | (~ main_stage_v_4) |
      io_read_cfg_mul_bypass_rsc_svs_8 | IsNaN_8U_23U_land_3_lpi_1_dfm_11 | mul_loop_mul_if_land_3_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_3_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_3_lpi_1_dfm_9 | FpMul_8U_23U_lor_20_lpi_1_dfm_7 | (~
      FpMul_8U_23U_FpMul_8U_23U_and_65_itm_2));
  assign mux_574_nl = MUX_s_1_2_2((nor_1311_nl), (mux_573_nl), or_309_cse);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_2_cse = core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse
      & (mux_574_nl);
  assign and_733_nl = and_dcpl_187 & and_dcpl_85;
  assign and_734_nl = and_dcpl_187 & or_90_cse;
  assign mux_1619_nl = MUX_s_1_2_2(IsNaN_8U_23U_1_land_4_lpi_1_dfm_9, IsNaN_8U_23U_1_land_4_lpi_1_dfm_8,
      or_309_cse);
  assign FpMul_8U_23U_p_expo_mux1h_7_itm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_4_sva_1_mx0w0,
      FpMul_8U_23U_p_expo_4_sva_1, ({4'b0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_10}),
      {(and_733_nl) , (and_734_nl) , (mux_1619_nl)});
  assign or_4956_cse = (~ (mul_loop_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) |
      mul_loop_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  assign or_4771_nl = (or_4956_cse & mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2)
      | FpMul_8U_23U_lor_21_lpi_1_dfm_6;
  assign and_2578_nl = FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_4_sva_st_2
      & mul_loop_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
      & or_tmp_1137;
  assign mux_1704_nl = MUX_s_1_2_2((and_2578_nl), or_tmp_1137, FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm);
  assign mux_1705_cse = MUX_s_1_2_2((mux_1704_nl), (or_4771_nl), nor_53_cse);
  assign nor_177_cse = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_4_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_21_lpi_1_dfm_st_3
      | (~ mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign or_1253_cse = (~ mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_21_lpi_1_dfm_st_3;
  assign nor_1291_nl = ~(IsNaN_8U_23U_land_4_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_4_lpi_1_dfm_10
      | (~ IsNaN_8U_23U_1_land_4_lpi_1_dfm_8) | mul_loop_mul_if_land_4_lpi_1_dfm_st_7
      | mul_loop_mul_if_land_4_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign nor_1292_nl = ~((~ IsNaN_8U_23U_1_land_4_lpi_1_dfm_9) | IsNaN_8U_23U_land_4_lpi_1_dfm_st_8
      | IsNaN_8U_23U_land_4_lpi_1_dfm_11 | mul_loop_mul_if_land_4_lpi_1_dfm_st_8
      | mul_loop_mul_if_land_4_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4));
  assign mux_590_nl = MUX_s_1_2_2((nor_1292_nl), (nor_1291_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_102_cse = core_wen & (~ and_dcpl_50)
      & (mux_590_nl);
  assign nor_181_cse = ~(FpMul_8U_23U_lor_21_lpi_1_dfm_st_3 | (~ mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1287_cse = ~((~ (mul_loop_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7);
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_25_cse = MUX_s_1_2_2(mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs_mx0w0,
      mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs, and_dcpl_104);
  assign nor_1283_nl = ~(IsNaN_8U_23U_land_4_lpi_1_dfm_10 | (~ IsNaN_8U_23U_1_land_4_lpi_1_dfm_8)
      | mul_loop_mul_if_land_4_lpi_1_dfm_st_7 | mul_loop_mul_if_land_4_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3));
  assign nor_1284_nl = ~((~ IsNaN_8U_23U_1_land_4_lpi_1_dfm_9) | IsNaN_8U_23U_land_4_lpi_1_dfm_11
      | mul_loop_mul_if_land_4_lpi_1_dfm_st_8 | mul_loop_mul_if_land_4_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4));
  assign mux_595_nl = MUX_s_1_2_2((nor_1284_nl), (nor_1283_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_105_cse = core_wen & (~ and_dcpl_50)
      & (mux_595_nl);
  assign IsNaN_8U_23U_aelse_and_54_cse = core_wen & (~ and_dcpl_50) & (~ mux_596_itm);
  assign nor_1277_nl = ~(nor_1287_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_4_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_4_lpi_1_dfm_10
      | FpMul_8U_23U_lor_21_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_4_lpi_1_dfm_8
      | mul_loop_mul_if_land_4_lpi_1_dfm_9);
  assign nor_1279_nl = ~((FpMul_8U_23U_p_mant_p1_4_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_4_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_4_lpi_1_dfm_10 | FpMul_8U_23U_lor_21_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_4_lpi_1_dfm_8 | mul_loop_mul_if_land_4_lpi_1_dfm_9);
  assign mux_598_nl = MUX_s_1_2_2((nor_1279_nl), (nor_1277_nl), nor_181_cse);
  assign and_2210_nl = mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_598_nl);
  assign nor_1280_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_66_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_4_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_4_lpi_1_dfm_10 | FpMul_8U_23U_lor_21_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_4_lpi_1_dfm_8 | mul_loop_mul_if_land_4_lpi_1_dfm_9);
  assign mux_599_nl = MUX_s_1_2_2((nor_1280_nl), (and_2210_nl), nor_53_cse);
  assign nor_1281_nl = ~((~((~ mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs_2) |
      mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs_st_2)) | (~ main_stage_v_4) |
      io_read_cfg_mul_bypass_rsc_svs_8 | IsNaN_8U_23U_land_4_lpi_1_dfm_11 | mul_loop_mul_if_land_4_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_4_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_4_lpi_1_dfm_9 | FpMul_8U_23U_lor_21_lpi_1_dfm_7 | (~
      FpMul_8U_23U_FpMul_8U_23U_and_66_itm_2));
  assign mux_600_nl = MUX_s_1_2_2((nor_1281_nl), (mux_599_nl), or_309_cse);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_3_cse = core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse
      & (mux_600_nl);
  assign and_738_nl = and_dcpl_192 & and_dcpl_85;
  assign and_739_nl = and_dcpl_192 & or_90_cse;
  assign mux_1620_nl = MUX_s_1_2_2(IsNaN_8U_23U_1_land_5_lpi_1_dfm_9, IsNaN_8U_23U_1_land_5_lpi_1_dfm_8,
      or_309_cse);
  assign FpMul_8U_23U_p_expo_mux1h_9_itm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_5_sva_1_mx0w0,
      FpMul_8U_23U_p_expo_5_sva_1, ({4'b0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_10}),
      {(and_738_nl) , (and_739_nl) , (mux_1620_nl)});
  assign or_4953_cse = (~ (mul_loop_mul_5_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) |
      mul_loop_mul_5_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  assign or_4783_nl = (or_4953_cse & mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2)
      | FpMul_8U_23U_lor_22_lpi_1_dfm_6;
  assign and_2600_nl = FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_5_sva_st_2
      & mul_loop_mul_5_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
      & or_tmp_1220;
  assign mux_1709_nl = MUX_s_1_2_2((and_2600_nl), or_tmp_1220, FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_4_itm);
  assign mux_1710_cse = MUX_s_1_2_2((mux_1709_nl), (or_4783_nl), nor_53_cse);
  assign nor_193_cse = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_5_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_22_lpi_1_dfm_st_3
      | (~ mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1259_nl = ~(IsNaN_8U_23U_land_5_lpi_1_dfm_st_7 | (~ IsNaN_8U_23U_1_land_5_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_5_lpi_1_dfm_10 | mul_loop_mul_if_land_5_lpi_1_dfm_st_7
      | mul_loop_mul_if_land_5_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign nor_1260_nl = ~(IsNaN_8U_23U_land_5_lpi_1_dfm_st_8 | IsNaN_8U_23U_land_5_lpi_1_dfm_11
      | (~ IsNaN_8U_23U_1_land_5_lpi_1_dfm_9) | mul_loop_mul_if_land_5_lpi_1_dfm_st_8
      | mul_loop_mul_if_land_5_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4));
  assign mux_614_nl = MUX_s_1_2_2((nor_1260_nl), (nor_1259_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_104_cse = core_wen & (~ and_dcpl_50)
      & (mux_614_nl);
  assign nor_197_cse = ~(FpMul_8U_23U_lor_22_lpi_1_dfm_st_3 | (~ mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1255_cse = ~((~ (mul_loop_mul_5_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_5_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7);
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_23_cse = MUX_s_1_2_2(mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs_mx0w0,
      mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs, and_dcpl_104);
  assign nor_1251_nl = ~((~ IsNaN_8U_23U_1_land_5_lpi_1_dfm_8) | IsNaN_8U_23U_land_5_lpi_1_dfm_10
      | mul_loop_mul_if_land_5_lpi_1_dfm_st_7 | mul_loop_mul_if_land_5_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3));
  assign nor_1252_nl = ~(IsNaN_8U_23U_land_5_lpi_1_dfm_11 | (~ IsNaN_8U_23U_1_land_5_lpi_1_dfm_9)
      | mul_loop_mul_if_land_5_lpi_1_dfm_st_8 | mul_loop_mul_if_land_5_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4));
  assign mux_619_nl = MUX_s_1_2_2((nor_1252_nl), (nor_1251_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_108_cse = core_wen & (~ and_dcpl_50)
      & (mux_619_nl);
  assign IsNaN_8U_23U_aelse_and_56_cse = core_wen & (~ and_dcpl_50) & (~ mux_620_itm);
  assign nor_1245_nl = ~(nor_1255_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_5_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_5_lpi_1_dfm_10
      | FpMul_8U_23U_lor_22_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_5_lpi_1_dfm_8
      | mul_loop_mul_if_land_5_lpi_1_dfm_9);
  assign nor_1247_nl = ~((FpMul_8U_23U_p_mant_p1_5_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_5_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_5_lpi_1_dfm_10 | FpMul_8U_23U_lor_22_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_5_lpi_1_dfm_8 | mul_loop_mul_if_land_5_lpi_1_dfm_9);
  assign mux_622_nl = MUX_s_1_2_2((nor_1247_nl), (nor_1245_nl), nor_197_cse);
  assign and_2204_nl = mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_622_nl);
  assign nor_1248_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_67_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_5_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_5_lpi_1_dfm_10 | FpMul_8U_23U_lor_22_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_5_lpi_1_dfm_8 | mul_loop_mul_if_land_5_lpi_1_dfm_9);
  assign mux_623_nl = MUX_s_1_2_2((nor_1248_nl), (and_2204_nl), nor_53_cse);
  assign nor_1249_nl = ~((~((~ mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs_2) |
      mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs_st_2)) | (~ main_stage_v_4) |
      io_read_cfg_mul_bypass_rsc_svs_8 | IsNaN_8U_23U_land_5_lpi_1_dfm_11 | mul_loop_mul_if_land_5_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_5_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_5_lpi_1_dfm_9 | FpMul_8U_23U_lor_22_lpi_1_dfm_7 | (~
      FpMul_8U_23U_FpMul_8U_23U_and_67_itm_2));
  assign mux_624_nl = MUX_s_1_2_2((nor_1249_nl), (mux_623_nl), or_309_cse);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_4_cse = core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse
      & (mux_624_nl);
  assign and_743_nl = and_dcpl_197 & and_dcpl_85;
  assign and_744_nl = and_dcpl_197 & or_90_cse;
  assign mux_1621_nl = MUX_s_1_2_2(IsNaN_8U_23U_1_land_6_lpi_1_dfm_9, IsNaN_8U_23U_1_land_6_lpi_1_dfm_8,
      or_309_cse);
  assign FpMul_8U_23U_p_expo_mux1h_11_itm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_6_sva_1_mx0w0,
      FpMul_8U_23U_p_expo_6_sva_1, ({4'b0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_10}),
      {(and_743_nl) , (and_744_nl) , (mux_1621_nl)});
  assign and_2876_cse = ((~ (mul_loop_mul_6_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_6_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7) & mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign or_4795_nl = and_2876_cse | FpMul_8U_23U_lor_23_lpi_1_dfm_6;
  assign and_2622_nl = FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_6_sva_st_2
      & mul_loop_mul_6_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
      & or_tmp_1300;
  assign mux_1714_nl = MUX_s_1_2_2((and_2622_nl), or_tmp_1300, FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_5_itm);
  assign mux_1715_cse = MUX_s_1_2_2((mux_1714_nl), (or_4795_nl), nor_53_cse);
  assign nor_209_cse = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_6_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_23_lpi_1_dfm_st_3
      | (~ mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1225_nl = ~(IsNaN_8U_23U_land_6_lpi_1_dfm_st_7 | (~ IsNaN_8U_23U_1_land_6_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_6_lpi_1_dfm_10 | mul_loop_mul_if_land_6_lpi_1_dfm_st_7
      | mul_loop_mul_if_land_6_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign nor_1226_nl = ~((~ IsNaN_8U_23U_1_land_6_lpi_1_dfm_9) | IsNaN_8U_23U_land_6_lpi_1_dfm_st_8
      | IsNaN_8U_23U_land_6_lpi_1_dfm_11 | mul_loop_mul_if_land_6_lpi_1_dfm_st_8
      | mul_loop_mul_if_land_6_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4));
  assign mux_638_nl = MUX_s_1_2_2((nor_1226_nl), (nor_1225_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_106_cse = core_wen & (~ and_dcpl_50)
      & (mux_638_nl);
  assign nor_1221_cse = ~((~ (mul_loop_mul_6_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_6_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7);
  assign nor_213_cse = ~(FpMul_8U_23U_lor_23_lpi_1_dfm_st_3 | (~ mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_21_cse = MUX_s_1_2_2(mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs_mx0w0,
      mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs, and_dcpl_104);
  assign nor_1217_nl = ~((~ IsNaN_8U_23U_1_land_6_lpi_1_dfm_8) | IsNaN_8U_23U_land_6_lpi_1_dfm_10
      | mul_loop_mul_if_land_6_lpi_1_dfm_st_7 | mul_loop_mul_if_land_6_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3));
  assign nor_1218_nl = ~((~ IsNaN_8U_23U_1_land_6_lpi_1_dfm_9) | IsNaN_8U_23U_land_6_lpi_1_dfm_11
      | mul_loop_mul_if_land_6_lpi_1_dfm_st_8 | mul_loop_mul_if_land_6_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4));
  assign mux_643_nl = MUX_s_1_2_2((nor_1218_nl), (nor_1217_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_111_cse = core_wen & (~ and_dcpl_50)
      & (mux_643_nl);
  assign IsNaN_8U_23U_aelse_and_58_cse = core_wen & (~ and_dcpl_50) & (~ mux_644_itm);
  assign nor_1211_nl = ~(nor_1221_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_6_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_6_lpi_1_dfm_10
      | FpMul_8U_23U_lor_23_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_6_lpi_1_dfm_8
      | mul_loop_mul_if_land_6_lpi_1_dfm_9);
  assign nor_1213_nl = ~((FpMul_8U_23U_p_mant_p1_6_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_6_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_6_lpi_1_dfm_10 | FpMul_8U_23U_lor_23_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_6_lpi_1_dfm_8 | mul_loop_mul_if_land_6_lpi_1_dfm_9);
  assign mux_646_nl = MUX_s_1_2_2((nor_1213_nl), (nor_1211_nl), nor_213_cse);
  assign and_2198_nl = mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_646_nl);
  assign nor_1214_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_68_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_6_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_6_lpi_1_dfm_10 | FpMul_8U_23U_lor_23_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_6_lpi_1_dfm_8 | mul_loop_mul_if_land_6_lpi_1_dfm_9);
  assign mux_647_nl = MUX_s_1_2_2((nor_1214_nl), (and_2198_nl), nor_53_cse);
  assign nor_1215_nl = ~((~((~ mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs_2) |
      mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs_st_2)) | (~ main_stage_v_4) |
      io_read_cfg_mul_bypass_rsc_svs_8 | IsNaN_8U_23U_land_6_lpi_1_dfm_11 | mul_loop_mul_if_land_6_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_6_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_6_lpi_1_dfm_9 | FpMul_8U_23U_lor_23_lpi_1_dfm_7 | (~
      FpMul_8U_23U_FpMul_8U_23U_and_68_itm_2));
  assign mux_648_nl = MUX_s_1_2_2((nor_1215_nl), (mux_647_nl), or_309_cse);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_5_cse = core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse
      & (mux_648_nl);
  assign and_748_nl = and_dcpl_202 & and_dcpl_85;
  assign and_749_nl = and_dcpl_202 & or_90_cse;
  assign mux_1622_nl = MUX_s_1_2_2(IsNaN_8U_23U_1_land_7_lpi_1_dfm_9, IsNaN_8U_23U_1_land_7_lpi_1_dfm_8,
      or_309_cse);
  assign FpMul_8U_23U_p_expo_mux1h_13_itm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_7_sva_1_mx0w0,
      FpMul_8U_23U_p_expo_7_sva_1, ({4'b0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_10}),
      {(and_748_nl) , (and_749_nl) , (mux_1622_nl)});
  assign or_4947_cse = (~ (mul_loop_mul_7_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) |
      mul_loop_mul_7_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  assign or_4807_nl = (or_4947_cse & mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2)
      | FpMul_8U_23U_lor_24_lpi_1_dfm_6;
  assign and_2644_nl = FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_7_sva_st_2
      & mul_loop_mul_7_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
      & or_tmp_1382;
  assign mux_1719_nl = MUX_s_1_2_2((and_2644_nl), or_tmp_1382, FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_6_itm);
  assign mux_1720_cse = MUX_s_1_2_2((mux_1719_nl), (or_4807_nl), nor_53_cse);
  assign nor_225_cse = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_7_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_24_lpi_1_dfm_st_3
      | (~ mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1191_nl = ~(IsNaN_8U_23U_land_7_lpi_1_dfm_st_7 | (~ IsNaN_8U_23U_1_land_7_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_7_lpi_1_dfm_10 | mul_loop_mul_if_land_7_lpi_1_dfm_st_7
      | mul_loop_mul_if_land_7_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign nor_1192_nl = ~(IsNaN_8U_23U_land_7_lpi_1_dfm_st_8 | (~ IsNaN_8U_23U_1_land_7_lpi_1_dfm_9)
      | IsNaN_8U_23U_land_7_lpi_1_dfm_11 | mul_loop_mul_if_land_7_lpi_1_dfm_st_8
      | mul_loop_mul_if_land_7_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4));
  assign mux_662_nl = MUX_s_1_2_2((nor_1192_nl), (nor_1191_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_108_cse = core_wen & (~ and_dcpl_50)
      & (mux_662_nl);
  assign nor_229_cse = ~(FpMul_8U_23U_lor_24_lpi_1_dfm_st_3 | (~ mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1187_cse = ~((~ (mul_loop_mul_7_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_7_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7);
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_19_cse = MUX_s_1_2_2(mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs_mx0w0,
      mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs, and_dcpl_104);
  assign nor_1183_nl = ~((~ IsNaN_8U_23U_1_land_7_lpi_1_dfm_8) | IsNaN_8U_23U_land_7_lpi_1_dfm_10
      | mul_loop_mul_if_land_7_lpi_1_dfm_st_7 | mul_loop_mul_if_land_7_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3));
  assign nor_1184_nl = ~((~ IsNaN_8U_23U_1_land_7_lpi_1_dfm_9) | IsNaN_8U_23U_land_7_lpi_1_dfm_11
      | mul_loop_mul_if_land_7_lpi_1_dfm_st_8 | mul_loop_mul_if_land_7_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4));
  assign mux_667_nl = MUX_s_1_2_2((nor_1184_nl), (nor_1183_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_114_cse = core_wen & (~ and_dcpl_50)
      & (mux_667_nl);
  assign IsNaN_8U_23U_aelse_and_60_cse = core_wen & (~ and_dcpl_50) & (~ mux_668_itm);
  assign nor_1177_nl = ~(nor_1187_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_7_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_7_lpi_1_dfm_10
      | FpMul_8U_23U_lor_24_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_7_lpi_1_dfm_8
      | mul_loop_mul_if_land_7_lpi_1_dfm_9);
  assign nor_1179_nl = ~((FpMul_8U_23U_p_mant_p1_7_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_7_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_7_lpi_1_dfm_10 | FpMul_8U_23U_lor_24_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_7_lpi_1_dfm_8 | mul_loop_mul_if_land_7_lpi_1_dfm_9);
  assign mux_670_nl = MUX_s_1_2_2((nor_1179_nl), (nor_1177_nl), nor_229_cse);
  assign and_2192_nl = mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_670_nl);
  assign nor_1180_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_69_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_7_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_7_lpi_1_dfm_10 | FpMul_8U_23U_lor_24_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_7_lpi_1_dfm_8 | mul_loop_mul_if_land_7_lpi_1_dfm_9);
  assign mux_671_nl = MUX_s_1_2_2((nor_1180_nl), (and_2192_nl), nor_53_cse);
  assign nor_1181_nl = ~((~((~ mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs_2) |
      mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs_st_2)) | (~ main_stage_v_4) |
      io_read_cfg_mul_bypass_rsc_svs_8 | IsNaN_8U_23U_land_7_lpi_1_dfm_11 | mul_loop_mul_if_land_7_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_7_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_7_lpi_1_dfm_9 | FpMul_8U_23U_lor_24_lpi_1_dfm_7 | (~
      FpMul_8U_23U_FpMul_8U_23U_and_69_itm_2));
  assign mux_672_nl = MUX_s_1_2_2((nor_1181_nl), (mux_671_nl), or_309_cse);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_6_cse = core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse
      & (mux_672_nl);
  assign and_753_nl = and_dcpl_207 & and_dcpl_85;
  assign and_754_nl = and_dcpl_207 & or_90_cse;
  assign mux_1623_nl = MUX_s_1_2_2(IsNaN_8U_23U_1_land_8_lpi_1_dfm_9, IsNaN_8U_23U_1_land_8_lpi_1_dfm_8,
      or_309_cse);
  assign FpMul_8U_23U_p_expo_mux1h_15_itm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_8_sva_1_mx0w0,
      FpMul_8U_23U_p_expo_8_sva_1, ({4'b0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_10}),
      {(and_753_nl) , (and_754_nl) , (mux_1623_nl)});
  assign or_4944_cse = (~ (mul_loop_mul_8_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) |
      mul_loop_mul_8_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  assign or_4819_nl = (or_4944_cse & mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2)
      | FpMul_8U_23U_lor_25_lpi_1_dfm_6;
  assign and_2666_nl = FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_8_sva_st_2
      & mul_loop_mul_8_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
      & or_tmp_1464;
  assign mux_1724_nl = MUX_s_1_2_2((and_2666_nl), or_tmp_1464, FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_7_itm);
  assign mux_1725_cse = MUX_s_1_2_2((mux_1724_nl), (or_4819_nl), nor_53_cse);
  assign nor_241_cse = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_8_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_25_lpi_1_dfm_st_3
      | (~ mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1159_nl = ~(IsNaN_8U_23U_land_8_lpi_1_dfm_st_7 | (~ IsNaN_8U_23U_1_land_8_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_8_lpi_1_dfm_10 | mul_loop_mul_if_land_8_lpi_1_dfm_st_7
      | mul_loop_mul_if_land_8_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign nor_1160_nl = ~((~ IsNaN_8U_23U_1_land_8_lpi_1_dfm_9) | IsNaN_8U_23U_land_8_lpi_1_dfm_st_8
      | IsNaN_8U_23U_land_8_lpi_1_dfm_11 | mul_loop_mul_if_land_8_lpi_1_dfm_st_8
      | mul_loop_mul_if_land_8_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4));
  assign mux_686_nl = MUX_s_1_2_2((nor_1160_nl), (nor_1159_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_110_cse = core_wen & (~ and_dcpl_50)
      & (mux_686_nl);
  assign nor_245_cse = ~(FpMul_8U_23U_lor_25_lpi_1_dfm_st_3 | (~ mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1155_cse = ~((~ (mul_loop_mul_8_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_8_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7);
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_17_cse = MUX_s_1_2_2(mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs_mx0w0,
      mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs, and_dcpl_104);
  assign nor_1151_nl = ~((~ IsNaN_8U_23U_1_land_8_lpi_1_dfm_8) | IsNaN_8U_23U_land_8_lpi_1_dfm_10
      | mul_loop_mul_if_land_8_lpi_1_dfm_st_7 | mul_loop_mul_if_land_8_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3));
  assign nor_1152_nl = ~((~ IsNaN_8U_23U_1_land_8_lpi_1_dfm_9) | IsNaN_8U_23U_land_8_lpi_1_dfm_11
      | mul_loop_mul_if_land_8_lpi_1_dfm_st_8 | mul_loop_mul_if_land_8_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4));
  assign mux_691_nl = MUX_s_1_2_2((nor_1152_nl), (nor_1151_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_117_cse = core_wen & (~ and_dcpl_50)
      & (mux_691_nl);
  assign IsNaN_8U_23U_aelse_and_62_cse = core_wen & (~ and_dcpl_50) & (~ mux_692_itm);
  assign nor_1145_nl = ~(nor_1155_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_8_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_8_lpi_1_dfm_10
      | FpMul_8U_23U_lor_25_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_8_lpi_1_dfm_8
      | mul_loop_mul_if_land_8_lpi_1_dfm_9);
  assign nor_1147_nl = ~((FpMul_8U_23U_p_mant_p1_8_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_8_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_8_lpi_1_dfm_10 | FpMul_8U_23U_lor_25_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_8_lpi_1_dfm_8 | mul_loop_mul_if_land_8_lpi_1_dfm_9);
  assign mux_694_nl = MUX_s_1_2_2((nor_1147_nl), (nor_1145_nl), nor_245_cse);
  assign and_2186_nl = mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_694_nl);
  assign nor_1148_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_70_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_8_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_8_lpi_1_dfm_10 | FpMul_8U_23U_lor_25_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_8_lpi_1_dfm_8 | mul_loop_mul_if_land_8_lpi_1_dfm_9);
  assign mux_695_nl = MUX_s_1_2_2((nor_1148_nl), (and_2186_nl), nor_53_cse);
  assign nor_1149_nl = ~((~((~ mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs_2) |
      mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs_st_2)) | (~ main_stage_v_4) |
      io_read_cfg_mul_bypass_rsc_svs_8 | IsNaN_8U_23U_land_8_lpi_1_dfm_11 | mul_loop_mul_if_land_8_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_8_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_8_lpi_1_dfm_9 | FpMul_8U_23U_lor_25_lpi_1_dfm_7 | (~
      FpMul_8U_23U_FpMul_8U_23U_and_70_itm_2));
  assign mux_696_nl = MUX_s_1_2_2((nor_1149_nl), (mux_695_nl), or_309_cse);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_7_cse = core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse
      & (mux_696_nl);
  assign and_758_nl = and_dcpl_212 & and_dcpl_85;
  assign and_759_nl = and_dcpl_212 & or_90_cse;
  assign mux_1624_nl = MUX_s_1_2_2(IsNaN_8U_23U_1_land_9_lpi_1_dfm_9, IsNaN_8U_23U_1_land_9_lpi_1_dfm_8,
      or_309_cse);
  assign FpMul_8U_23U_p_expo_mux1h_17_itm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_9_sva_1_mx0w0,
      FpMul_8U_23U_p_expo_9_sva_1, ({4'b0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_10}),
      {(and_758_nl) , (and_759_nl) , (mux_1624_nl)});
  assign or_4941_cse = (~ (mul_loop_mul_9_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) |
      mul_loop_mul_9_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  assign or_4831_nl = (or_4941_cse & mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2)
      | FpMul_8U_23U_lor_26_lpi_1_dfm_6;
  assign and_2688_nl = FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_9_sva_st_2
      & mul_loop_mul_9_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
      & or_tmp_1544;
  assign mux_1729_nl = MUX_s_1_2_2((and_2688_nl), or_tmp_1544, FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_8_itm);
  assign mux_1730_cse = MUX_s_1_2_2((mux_1729_nl), (or_4831_nl), nor_53_cse);
  assign nor_257_cse = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_9_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_26_lpi_1_dfm_st_3
      | (~ mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1127_nl = ~(IsNaN_8U_23U_land_9_lpi_1_dfm_st_7 | (~ IsNaN_8U_23U_1_land_9_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_9_lpi_1_dfm_10 | mul_loop_mul_if_land_9_lpi_1_dfm_st_7
      | mul_loop_mul_if_land_9_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign nor_1128_nl = ~((~ IsNaN_8U_23U_1_land_9_lpi_1_dfm_9) | IsNaN_8U_23U_land_9_lpi_1_dfm_st_8
      | IsNaN_8U_23U_land_9_lpi_1_dfm_11 | mul_loop_mul_if_land_9_lpi_1_dfm_st_8
      | mul_loop_mul_if_land_9_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4));
  assign mux_710_nl = MUX_s_1_2_2((nor_1128_nl), (nor_1127_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_112_cse = core_wen & (~ and_dcpl_50)
      & (mux_710_nl);
  assign nor_261_cse = ~(FpMul_8U_23U_lor_26_lpi_1_dfm_st_3 | (~ mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1123_cse = ~((~ (mul_loop_mul_9_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_9_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7);
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_15_cse = MUX_s_1_2_2(mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs_mx0w0,
      mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs, and_dcpl_104);
  assign nor_1119_nl = ~((~ IsNaN_8U_23U_1_land_9_lpi_1_dfm_8) | IsNaN_8U_23U_land_9_lpi_1_dfm_10
      | mul_loop_mul_if_land_9_lpi_1_dfm_st_7 | mul_loop_mul_if_land_9_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3));
  assign nor_1120_nl = ~((~ IsNaN_8U_23U_1_land_9_lpi_1_dfm_9) | IsNaN_8U_23U_land_9_lpi_1_dfm_11
      | mul_loop_mul_if_land_9_lpi_1_dfm_st_8 | mul_loop_mul_if_land_9_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4));
  assign mux_715_nl = MUX_s_1_2_2((nor_1120_nl), (nor_1119_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_120_cse = core_wen & (~ and_dcpl_50)
      & (mux_715_nl);
  assign IsNaN_8U_23U_aelse_and_64_cse = core_wen & (~ and_dcpl_50) & (~ mux_716_itm);
  assign nor_1113_nl = ~(nor_1123_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_9_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_9_lpi_1_dfm_10
      | FpMul_8U_23U_lor_26_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_9_lpi_1_dfm_8
      | mul_loop_mul_if_land_9_lpi_1_dfm_9);
  assign nor_1115_nl = ~((FpMul_8U_23U_p_mant_p1_9_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_9_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_9_lpi_1_dfm_10 | FpMul_8U_23U_lor_26_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_9_lpi_1_dfm_8 | mul_loop_mul_if_land_9_lpi_1_dfm_9);
  assign mux_718_nl = MUX_s_1_2_2((nor_1115_nl), (nor_1113_nl), nor_261_cse);
  assign and_2180_nl = mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_718_nl);
  assign nor_1116_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_71_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_9_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_9_lpi_1_dfm_10 | FpMul_8U_23U_lor_26_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_9_lpi_1_dfm_8 | mul_loop_mul_if_land_9_lpi_1_dfm_9);
  assign mux_719_nl = MUX_s_1_2_2((nor_1116_nl), (and_2180_nl), nor_53_cse);
  assign nor_1117_nl = ~((~((~ mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs_2) |
      mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs_st_2)) | (~ main_stage_v_4) |
      io_read_cfg_mul_bypass_rsc_svs_8 | IsNaN_8U_23U_land_9_lpi_1_dfm_11 | mul_loop_mul_if_land_9_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_9_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_9_lpi_1_dfm_9 | FpMul_8U_23U_lor_26_lpi_1_dfm_7 | (~
      FpMul_8U_23U_FpMul_8U_23U_and_71_itm_2));
  assign mux_720_nl = MUX_s_1_2_2((nor_1117_nl), (mux_719_nl), or_309_cse);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_8_cse = core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse
      & (mux_720_nl);
  assign and_763_nl = and_dcpl_217 & and_dcpl_85;
  assign and_764_nl = and_dcpl_217 & or_90_cse;
  assign mux_1625_nl = MUX_s_1_2_2(IsNaN_8U_23U_1_land_10_lpi_1_dfm_9, IsNaN_8U_23U_1_land_10_lpi_1_dfm_8,
      or_309_cse);
  assign FpMul_8U_23U_p_expo_mux1h_19_itm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_10_sva_1_mx0w0,
      FpMul_8U_23U_p_expo_10_sva_1, ({4'b0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_10}),
      {(and_763_nl) , (and_764_nl) , (mux_1625_nl)});
  assign and_2868_cse = ((~ (mul_loop_mul_10_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_10_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7) & mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign or_4843_nl = and_2868_cse | FpMul_8U_23U_lor_27_lpi_1_dfm_6;
  assign and_2710_nl = FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_10_sva_st_2
      & mul_loop_mul_10_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
      & or_tmp_1624;
  assign mux_1734_nl = MUX_s_1_2_2((and_2710_nl), or_tmp_1624, FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_9_itm);
  assign mux_1735_cse = MUX_s_1_2_2((mux_1734_nl), (or_4843_nl), nor_53_cse);
  assign nor_273_cse = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_10_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_27_lpi_1_dfm_st_3
      | (~ mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1103_cse = ~((~ mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs_2) |
      mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs_st_2);
  assign nor_1094_nl = ~(IsNaN_8U_23U_land_10_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_10_lpi_1_dfm_10
      | (~ IsNaN_8U_23U_1_land_10_lpi_1_dfm_8) | mul_loop_mul_if_land_10_lpi_1_dfm_st_7
      | mul_loop_mul_if_land_10_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7 |
      io_read_cfg_mul_bypass_rsc_svs_st_6 | (~ main_stage_v_3));
  assign nor_1095_nl = ~(IsNaN_8U_23U_land_10_lpi_1_dfm_st_8 | (~ IsNaN_8U_23U_1_land_10_lpi_1_dfm_9)
      | IsNaN_8U_23U_land_10_lpi_1_dfm_11 | mul_loop_mul_if_land_10_lpi_1_dfm_st_8
      | mul_loop_mul_if_land_10_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4));
  assign mux_734_nl = MUX_s_1_2_2((nor_1095_nl), (nor_1094_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_114_cse = core_wen & (~ and_dcpl_50)
      & (mux_734_nl);
  assign nor_1090_cse = ~((~ (mul_loop_mul_10_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_10_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7);
  assign nor_277_cse = ~(FpMul_8U_23U_lor_27_lpi_1_dfm_st_3 | (~ mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_13_cse = MUX_s_1_2_2(mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs_mx0w0,
      mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs, and_dcpl_104);
  assign nor_1086_nl = ~(IsNaN_8U_23U_land_10_lpi_1_dfm_10 | (~ IsNaN_8U_23U_1_land_10_lpi_1_dfm_8)
      | mul_loop_mul_if_land_10_lpi_1_dfm_st_7 | mul_loop_mul_if_land_10_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3));
  assign nor_1087_nl = ~((~ IsNaN_8U_23U_1_land_10_lpi_1_dfm_9) | IsNaN_8U_23U_land_10_lpi_1_dfm_11
      | mul_loop_mul_if_land_10_lpi_1_dfm_st_8 | mul_loop_mul_if_land_10_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4));
  assign mux_739_nl = MUX_s_1_2_2((nor_1087_nl), (nor_1086_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_123_cse = core_wen & (~ and_dcpl_50)
      & (mux_739_nl);
  assign IsNaN_8U_23U_aelse_and_66_cse = core_wen & (~ and_dcpl_50) & (~ mux_740_itm);
  assign nor_1080_nl = ~(nor_1090_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_10_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_10_lpi_1_dfm_10
      | FpMul_8U_23U_lor_27_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_10_lpi_1_dfm_8
      | mul_loop_mul_if_land_10_lpi_1_dfm_9);
  assign nor_1082_nl = ~((FpMul_8U_23U_p_mant_p1_10_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_10_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_10_lpi_1_dfm_10 | FpMul_8U_23U_lor_27_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_10_lpi_1_dfm_8 | mul_loop_mul_if_land_10_lpi_1_dfm_9);
  assign mux_742_nl = MUX_s_1_2_2((nor_1082_nl), (nor_1080_nl), nor_277_cse);
  assign and_2173_nl = mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_742_nl);
  assign nor_1083_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_72_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_10_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_10_lpi_1_dfm_10 | FpMul_8U_23U_lor_27_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_10_lpi_1_dfm_8 | mul_loop_mul_if_land_10_lpi_1_dfm_9);
  assign mux_743_nl = MUX_s_1_2_2((nor_1083_nl), (and_2173_nl), nor_53_cse);
  assign nor_1084_nl = ~(nor_1103_cse | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_10_lpi_1_dfm_11 | mul_loop_mul_if_land_10_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_10_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_10_lpi_1_dfm_9 | FpMul_8U_23U_lor_27_lpi_1_dfm_7 | (~
      FpMul_8U_23U_FpMul_8U_23U_and_72_itm_2));
  assign mux_744_nl = MUX_s_1_2_2((nor_1084_nl), (mux_743_nl), or_309_cse);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_9_cse = core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse
      & (mux_744_nl);
  assign nor_283_cse = ~(FpMul_8U_23U_lor_28_lpi_1_dfm_st_3 | (~ mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign and_768_nl = and_dcpl_222 & and_dcpl_85;
  assign and_769_nl = and_dcpl_222 & or_90_cse;
  assign mux_1626_nl = MUX_s_1_2_2(IsNaN_8U_23U_1_land_11_lpi_1_dfm_9, IsNaN_8U_23U_1_land_11_lpi_1_dfm_8,
      or_309_cse);
  assign FpMul_8U_23U_p_expo_mux1h_21_itm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_11_sva_1_mx0w0,
      FpMul_8U_23U_p_expo_11_sva_1, ({4'b0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_10}),
      {(and_768_nl) , (and_769_nl) , (mux_1626_nl)});
  assign or_4854_nl = (~ (mul_loop_mul_11_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) |
      mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 | FpMul_8U_23U_lor_28_lpi_1_dfm_6;
  assign mux_1739_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_28_lpi_1_dfm_6, (or_4854_nl),
      mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign and_2732_nl = mul_loop_mul_11_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
      & FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_11_sva_st_2
      & or_tmp_1703;
  assign mux_1740_nl = MUX_s_1_2_2((and_2732_nl), or_tmp_1703, FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_10_itm);
  assign mux_1741_cse = MUX_s_1_2_2((mux_1740_nl), (mux_1739_nl), nor_53_cse);
  assign nor_289_cse = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_11_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_28_lpi_1_dfm_st_3
      | (~ mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1070_cse = ~((~ mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs_2) |
      mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs_st_2);
  assign or_1819_cse = (~ mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_28_lpi_1_dfm_st_3;
  assign nor_1063_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_11_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_11_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_11_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | (~
      IsNaN_8U_23U_1_land_11_lpi_1_dfm_8) | mul_loop_mul_if_land_11_lpi_1_dfm_9);
  assign nor_1064_nl = ~((~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8 |
      IsNaN_8U_23U_land_11_lpi_1_dfm_11 | mul_loop_mul_if_land_11_lpi_1_dfm_10 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_11_lpi_1_dfm_st_8
      | (~ IsNaN_8U_23U_1_land_11_lpi_1_dfm_9) | IsNaN_8U_23U_land_11_lpi_1_dfm_st_8);
  assign mux_761_nl = MUX_s_1_2_2((nor_1064_nl), (nor_1063_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_116_cse = core_wen & (~ and_dcpl_50)
      & (mux_761_nl);
  assign nor_1059_cse = ~((~ (mul_loop_mul_11_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7);
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_11_cse = MUX_s_1_2_2(mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs_mx0w0,
      mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs, and_dcpl_104);
  assign nor_1055_nl = ~((~ IsNaN_8U_23U_1_land_11_lpi_1_dfm_8) | IsNaN_8U_23U_land_11_lpi_1_dfm_10
      | mul_loop_mul_if_land_11_lpi_1_dfm_st_7 | mul_loop_mul_if_land_11_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3));
  assign nor_1056_nl = ~((~ IsNaN_8U_23U_1_land_11_lpi_1_dfm_9) | IsNaN_8U_23U_land_11_lpi_1_dfm_11
      | mul_loop_mul_if_land_11_lpi_1_dfm_st_8 | mul_loop_mul_if_land_11_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4));
  assign mux_766_nl = MUX_s_1_2_2((nor_1056_nl), (nor_1055_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_126_cse = core_wen & (~ and_dcpl_50)
      & (mux_766_nl);
  assign IsNaN_8U_23U_aelse_and_68_cse = core_wen & (~ and_dcpl_50) & (~ mux_tmp_748);
  assign nor_1049_nl = ~(nor_1059_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_11_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_11_lpi_1_dfm_10
      | FpMul_8U_23U_lor_28_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_11_lpi_1_dfm_8
      | mul_loop_mul_if_land_11_lpi_1_dfm_9);
  assign nor_1051_nl = ~((FpMul_8U_23U_p_mant_p1_11_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_11_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_11_lpi_1_dfm_10 | FpMul_8U_23U_lor_28_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_11_lpi_1_dfm_8 | mul_loop_mul_if_land_11_lpi_1_dfm_9);
  assign mux_768_nl = MUX_s_1_2_2((nor_1051_nl), (nor_1049_nl), nor_283_cse);
  assign and_2164_nl = mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_768_nl);
  assign nor_1052_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_73_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_11_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_11_lpi_1_dfm_10 | FpMul_8U_23U_lor_28_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_11_lpi_1_dfm_8 | mul_loop_mul_if_land_11_lpi_1_dfm_9);
  assign mux_769_nl = MUX_s_1_2_2((nor_1052_nl), (and_2164_nl), nor_53_cse);
  assign nor_1053_nl = ~(nor_1070_cse | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_11_lpi_1_dfm_11 | mul_loop_mul_if_land_11_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_11_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_11_lpi_1_dfm_9 | FpMul_8U_23U_lor_28_lpi_1_dfm_7 | (~
      FpMul_8U_23U_FpMul_8U_23U_and_73_itm_2));
  assign mux_770_nl = MUX_s_1_2_2((nor_1053_nl), (mux_769_nl), or_309_cse);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_10_cse = core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse
      & (mux_770_nl);
  assign and_773_nl = and_dcpl_227 & and_dcpl_85;
  assign and_774_nl = and_dcpl_227 & or_90_cse;
  assign mux_1627_nl = MUX_s_1_2_2(IsNaN_8U_23U_1_land_12_lpi_1_dfm_9, IsNaN_8U_23U_1_land_12_lpi_1_dfm_8,
      or_309_cse);
  assign FpMul_8U_23U_p_expo_mux1h_23_itm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_12_sva_1_mx0w0,
      FpMul_8U_23U_p_expo_12_sva_1, ({4'b0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_10}),
      {(and_773_nl) , (and_774_nl) , (mux_1627_nl)});
  assign or_4934_cse = (~ (mul_loop_mul_12_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) |
      mul_loop_mul_12_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  assign or_4865_nl = (or_4934_cse & mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2)
      | FpMul_8U_23U_lor_29_lpi_1_dfm_6;
  assign and_2754_nl = FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_12_sva_st_2
      & mul_loop_mul_12_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
      & or_tmp_1782;
  assign mux_1746_nl = MUX_s_1_2_2((and_2754_nl), or_tmp_1782, FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_11_itm);
  assign mux_1747_cse = MUX_s_1_2_2((mux_1746_nl), (or_4865_nl), nor_53_cse);
  assign nor_305_cse = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_12_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_29_lpi_1_dfm_st_3
      | (~ mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1037_cse = ~((~ mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs_2) |
      mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs_st_2);
  assign or_1898_cse = (~ mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_29_lpi_1_dfm_st_3;
  assign nor_1030_nl = ~(IsNaN_8U_23U_land_12_lpi_1_dfm_st_7 | (~ IsNaN_8U_23U_1_land_12_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_12_lpi_1_dfm_10 | mul_loop_mul_if_land_12_lpi_1_dfm_st_7
      | mul_loop_mul_if_land_12_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7 |
      io_read_cfg_mul_bypass_rsc_svs_st_6 | (~ main_stage_v_3));
  assign nor_1031_nl = ~((~ IsNaN_8U_23U_1_land_12_lpi_1_dfm_9) | IsNaN_8U_23U_land_12_lpi_1_dfm_st_8
      | IsNaN_8U_23U_land_12_lpi_1_dfm_11 | mul_loop_mul_if_land_12_lpi_1_dfm_st_8
      | mul_loop_mul_if_land_12_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4));
  assign mux_787_nl = MUX_s_1_2_2((nor_1031_nl), (nor_1030_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_118_cse = core_wen & (~ and_dcpl_50)
      & (mux_787_nl);
  assign nor_309_cse = ~(FpMul_8U_23U_lor_29_lpi_1_dfm_st_3 | (~ mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1026_cse = ~((~ (mul_loop_mul_12_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_12_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7);
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_9_cse = MUX_s_1_2_2(mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs_mx0w0,
      mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs, and_dcpl_104);
  assign nor_1022_nl = ~((~ IsNaN_8U_23U_1_land_12_lpi_1_dfm_8) | IsNaN_8U_23U_land_12_lpi_1_dfm_10
      | mul_loop_mul_if_land_12_lpi_1_dfm_st_7 | mul_loop_mul_if_land_12_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3));
  assign nor_1023_nl = ~((~ IsNaN_8U_23U_1_land_12_lpi_1_dfm_9) | IsNaN_8U_23U_land_12_lpi_1_dfm_11
      | mul_loop_mul_if_land_12_lpi_1_dfm_st_8 | mul_loop_mul_if_land_12_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4));
  assign mux_792_nl = MUX_s_1_2_2((nor_1023_nl), (nor_1022_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_129_cse = core_wen & (~ and_dcpl_50)
      & (mux_792_nl);
  assign IsNaN_8U_23U_aelse_and_70_cse = core_wen & (~ and_dcpl_50) & (~ mux_793_itm);
  assign nor_1016_nl = ~(nor_1026_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_12_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_12_lpi_1_dfm_10
      | FpMul_8U_23U_lor_29_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_12_lpi_1_dfm_8
      | mul_loop_mul_if_land_12_lpi_1_dfm_9);
  assign nor_1018_nl = ~((FpMul_8U_23U_p_mant_p1_12_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_12_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_12_lpi_1_dfm_10 | FpMul_8U_23U_lor_29_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_12_lpi_1_dfm_8 | mul_loop_mul_if_land_12_lpi_1_dfm_9);
  assign mux_795_nl = MUX_s_1_2_2((nor_1018_nl), (nor_1016_nl), nor_309_cse);
  assign and_2158_nl = mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_795_nl);
  assign nor_1019_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_74_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_12_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_12_lpi_1_dfm_10 | FpMul_8U_23U_lor_29_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_12_lpi_1_dfm_8 | mul_loop_mul_if_land_12_lpi_1_dfm_9);
  assign mux_796_nl = MUX_s_1_2_2((nor_1019_nl), (and_2158_nl), nor_53_cse);
  assign nor_1020_nl = ~(nor_1037_cse | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_12_lpi_1_dfm_11 | mul_loop_mul_if_land_12_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_12_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_12_lpi_1_dfm_9 | FpMul_8U_23U_lor_29_lpi_1_dfm_7 | (~
      FpMul_8U_23U_FpMul_8U_23U_and_74_itm_2));
  assign mux_797_nl = MUX_s_1_2_2((nor_1020_nl), (mux_796_nl), or_309_cse);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_11_cse = core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse
      & (mux_797_nl);
  assign and_778_nl = and_dcpl_232 & and_dcpl_85;
  assign and_779_nl = and_dcpl_232 & or_90_cse;
  assign mux_1628_nl = MUX_s_1_2_2(IsNaN_8U_23U_1_land_13_lpi_1_dfm_9, IsNaN_8U_23U_1_land_13_lpi_1_dfm_8,
      or_309_cse);
  assign FpMul_8U_23U_p_expo_mux1h_25_itm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_13_sva_1_mx0w0,
      FpMul_8U_23U_p_expo_13_sva_1, ({4'b0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_10}),
      {(and_778_nl) , (and_779_nl) , (mux_1628_nl)});
  assign or_4931_cse = (~ (mul_loop_mul_13_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) |
      mul_loop_mul_13_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  assign or_4877_nl = (or_4931_cse & mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2)
      | FpMul_8U_23U_lor_30_lpi_1_dfm_6;
  assign and_2776_nl = FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_13_sva_st_2
      & mul_loop_mul_13_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
      & or_tmp_1865;
  assign mux_1751_nl = MUX_s_1_2_2((and_2776_nl), or_tmp_1865, FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_12_itm);
  assign mux_1752_cse = MUX_s_1_2_2((mux_1751_nl), (or_4877_nl), nor_53_cse);
  assign nor_321_cse = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_13_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_30_lpi_1_dfm_st_3
      | (~ mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_1004_cse = ~((~ mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs_2) |
      mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs_st_2);
  assign or_1981_cse = (~ mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_30_lpi_1_dfm_st_3;
  assign nor_997_nl = ~(IsNaN_8U_23U_land_13_lpi_1_dfm_st_7 | (~ IsNaN_8U_23U_1_land_13_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_13_lpi_1_dfm_10 | mul_loop_mul_if_land_13_lpi_1_dfm_st_7
      | mul_loop_mul_if_land_13_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7 |
      io_read_cfg_mul_bypass_rsc_svs_st_6 | (~ main_stage_v_3));
  assign nor_998_nl = ~((~ IsNaN_8U_23U_1_land_13_lpi_1_dfm_9) | IsNaN_8U_23U_land_13_lpi_1_dfm_st_8
      | IsNaN_8U_23U_land_13_lpi_1_dfm_11 | mul_loop_mul_if_land_13_lpi_1_dfm_st_8
      | mul_loop_mul_if_land_13_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4));
  assign mux_814_nl = MUX_s_1_2_2((nor_998_nl), (nor_997_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_120_cse = core_wen & (~ and_dcpl_50)
      & (mux_814_nl);
  assign nor_325_cse = ~(FpMul_8U_23U_lor_30_lpi_1_dfm_st_3 | (~ mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_993_cse = ~((~ (mul_loop_mul_13_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_13_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7);
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_7_cse = MUX_s_1_2_2(mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs_mx0w0,
      mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs, and_dcpl_104);
  assign nor_989_nl = ~((~ IsNaN_8U_23U_1_land_13_lpi_1_dfm_8) | IsNaN_8U_23U_land_13_lpi_1_dfm_10
      | mul_loop_mul_if_land_13_lpi_1_dfm_st_7 | mul_loop_mul_if_land_13_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3));
  assign nor_990_nl = ~((~ IsNaN_8U_23U_1_land_13_lpi_1_dfm_9) | IsNaN_8U_23U_land_13_lpi_1_dfm_11
      | mul_loop_mul_if_land_13_lpi_1_dfm_st_8 | mul_loop_mul_if_land_13_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4));
  assign mux_819_nl = MUX_s_1_2_2((nor_990_nl), (nor_989_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_132_cse = core_wen & (~ and_dcpl_50)
      & (mux_819_nl);
  assign IsNaN_8U_23U_aelse_and_72_cse = core_wen & (~ and_dcpl_50) & (~ mux_820_itm);
  assign nor_983_nl = ~(nor_993_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_13_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_13_lpi_1_dfm_10
      | FpMul_8U_23U_lor_30_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_13_lpi_1_dfm_8
      | mul_loop_mul_if_land_13_lpi_1_dfm_9);
  assign nor_985_nl = ~((FpMul_8U_23U_p_mant_p1_13_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_13_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_13_lpi_1_dfm_10 | FpMul_8U_23U_lor_30_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_13_lpi_1_dfm_8 | mul_loop_mul_if_land_13_lpi_1_dfm_9);
  assign mux_822_nl = MUX_s_1_2_2((nor_985_nl), (nor_983_nl), nor_325_cse);
  assign and_2152_nl = mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_822_nl);
  assign nor_986_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_75_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_13_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_13_lpi_1_dfm_10 | FpMul_8U_23U_lor_30_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_13_lpi_1_dfm_8 | mul_loop_mul_if_land_13_lpi_1_dfm_9);
  assign mux_823_nl = MUX_s_1_2_2((nor_986_nl), (and_2152_nl), nor_53_cse);
  assign nor_987_nl = ~(nor_1004_cse | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_13_lpi_1_dfm_11 | mul_loop_mul_if_land_13_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_13_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_13_lpi_1_dfm_9 | FpMul_8U_23U_lor_30_lpi_1_dfm_7 | (~
      FpMul_8U_23U_FpMul_8U_23U_and_75_itm_2));
  assign mux_824_nl = MUX_s_1_2_2((nor_987_nl), (mux_823_nl), or_309_cse);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_12_cse = core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse
      & (mux_824_nl);
  assign nor_332_cse = ~(mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      | (~ (mul_loop_mul_14_FpMul_8U_23U_p_mant_p1_mul_tmp[47])));
  assign and_783_nl = and_dcpl_237 & and_dcpl_85;
  assign and_784_nl = and_dcpl_237 & or_90_cse;
  assign mux_1629_nl = MUX_s_1_2_2(IsNaN_8U_23U_1_land_14_lpi_1_dfm_9, IsNaN_8U_23U_1_land_14_lpi_1_dfm_8,
      or_309_cse);
  assign FpMul_8U_23U_p_expo_mux1h_27_itm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_14_sva_1_mx0w0,
      FpMul_8U_23U_p_expo_14_sva_1, ({4'b0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_10}),
      {(and_783_nl) , (and_784_nl) , (mux_1629_nl)});
  assign or_4888_nl = mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      | (~ (mul_loop_mul_14_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) | FpMul_8U_23U_lor_31_lpi_1_dfm_6;
  assign mux_1756_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_31_lpi_1_dfm_6, (or_4888_nl),
      mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign and_2798_nl = FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_14_sva_st_2
      & mul_loop_mul_14_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
      & or_tmp_1947;
  assign mux_1757_nl = MUX_s_1_2_2((and_2798_nl), or_tmp_1947, FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_13_itm);
  assign mux_1758_cse = MUX_s_1_2_2((mux_1757_nl), (mux_1756_nl), nor_53_cse);
  assign nor_336_cse = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_14_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_31_lpi_1_dfm_st_3
      | (~ mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_972_cse = ~((~ mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs_2) | mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs_st_2);
  assign nor_961_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_14_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_14_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_14_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | (~
      IsNaN_8U_23U_1_land_14_lpi_1_dfm_8) | mul_loop_mul_if_land_14_lpi_1_dfm_9);
  assign nor_962_nl = ~((~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8 | IsNaN_8U_23U_land_14_lpi_1_dfm_11
      | mul_loop_mul_if_land_14_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | mul_loop_mul_if_land_14_lpi_1_dfm_st_8 | (~ IsNaN_8U_23U_1_land_14_lpi_1_dfm_9)
      | IsNaN_8U_23U_land_14_lpi_1_dfm_st_8);
  assign mux_839_nl = MUX_s_1_2_2((nor_962_nl), (nor_961_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_122_cse = core_wen & (~ and_dcpl_50)
      & (mux_839_nl);
  assign nor_340_cse = ~(FpMul_8U_23U_lor_31_lpi_1_dfm_st_3 | (~ mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_5_cse = MUX_s_1_2_2(mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs_mx0w0,
      mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs, and_dcpl_104);
  assign nor_953_nl = ~((~ IsNaN_8U_23U_1_land_14_lpi_1_dfm_8) | IsNaN_8U_23U_land_14_lpi_1_dfm_10
      | mul_loop_mul_if_land_14_lpi_1_dfm_st_7 | mul_loop_mul_if_land_14_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3));
  assign nor_954_nl = ~((~ IsNaN_8U_23U_1_land_14_lpi_1_dfm_9) | IsNaN_8U_23U_land_14_lpi_1_dfm_11
      | mul_loop_mul_if_land_14_lpi_1_dfm_st_8 | mul_loop_mul_if_land_14_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4));
  assign mux_844_nl = MUX_s_1_2_2((nor_954_nl), (nor_953_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_135_cse = core_wen & (~ and_dcpl_50)
      & (mux_844_nl);
  assign IsNaN_8U_23U_aelse_and_74_cse = core_wen & (~ and_dcpl_50) & (~ mux_845_itm);
  assign nor_947_nl = ~(nor_332_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_14_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_14_lpi_1_dfm_10
      | FpMul_8U_23U_lor_31_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_14_lpi_1_dfm_8
      | mul_loop_mul_if_land_14_lpi_1_dfm_9);
  assign nor_949_nl = ~((FpMul_8U_23U_p_mant_p1_14_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_14_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_14_lpi_1_dfm_10 | FpMul_8U_23U_lor_31_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_14_lpi_1_dfm_8 | mul_loop_mul_if_land_14_lpi_1_dfm_9);
  assign mux_847_nl = MUX_s_1_2_2((nor_949_nl), (nor_947_nl), nor_340_cse);
  assign and_2147_nl = mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_847_nl);
  assign nor_950_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_76_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_14_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_14_lpi_1_dfm_10 | FpMul_8U_23U_lor_31_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_14_lpi_1_dfm_8 | mul_loop_mul_if_land_14_lpi_1_dfm_9);
  assign mux_848_nl = MUX_s_1_2_2((nor_950_nl), (and_2147_nl), nor_53_cse);
  assign nor_951_nl = ~(nor_972_cse | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_14_lpi_1_dfm_11 | mul_loop_mul_if_land_14_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_14_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_14_lpi_1_dfm_9 | FpMul_8U_23U_lor_31_lpi_1_dfm_7 | (~
      FpMul_8U_23U_FpMul_8U_23U_and_76_itm_2));
  assign mux_849_nl = MUX_s_1_2_2((nor_951_nl), (mux_848_nl), or_309_cse);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_13_cse = core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse
      & (mux_849_nl);
  assign and_788_nl = and_dcpl_242 & and_dcpl_85;
  assign and_789_nl = and_dcpl_242 & or_90_cse;
  assign mux_1630_nl = MUX_s_1_2_2(IsNaN_8U_23U_1_land_15_lpi_1_dfm_9, IsNaN_8U_23U_1_land_15_lpi_1_dfm_8,
      or_309_cse);
  assign FpMul_8U_23U_p_expo_mux1h_29_itm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_15_sva_1_mx0w0,
      FpMul_8U_23U_p_expo_15_sva_1, ({4'b0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_10}),
      {(and_788_nl) , (and_789_nl) , (mux_1630_nl)});
  assign or_4927_cse = (~ (mul_loop_mul_15_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) |
      mul_loop_mul_15_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  assign or_4900_nl = (or_4927_cse & mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2)
      | FpMul_8U_23U_lor_32_lpi_1_dfm_6;
  assign and_2819_nl = FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_15_sva_st_2
      & mul_loop_mul_15_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
      & or_tmp_2032;
  assign mux_1763_nl = MUX_s_1_2_2((and_2819_nl), or_tmp_2032, FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_14_itm);
  assign mux_1764_cse = MUX_s_1_2_2((mux_1763_nl), (or_4900_nl), nor_53_cse);
  assign nor_352_cse = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_15_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_32_lpi_1_dfm_st_3
      | (~ mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_935_cse = ~((~ mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs_2) | mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs_st_2);
  assign nor_924_nl = ~(IsNaN_8U_23U_land_15_lpi_1_dfm_st_7 | (~ IsNaN_8U_23U_1_land_15_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_15_lpi_1_dfm_10 | mul_loop_mul_if_land_15_lpi_1_dfm_st_7
      | mul_loop_mul_if_land_15_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7 |
      io_read_cfg_mul_bypass_rsc_svs_st_6 | (~ main_stage_v_3));
  assign nor_925_nl = ~((~ IsNaN_8U_23U_1_land_15_lpi_1_dfm_9) | IsNaN_8U_23U_land_15_lpi_1_dfm_st_8
      | IsNaN_8U_23U_land_15_lpi_1_dfm_11 | mul_loop_mul_if_land_15_lpi_1_dfm_st_8
      | mul_loop_mul_if_land_15_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4));
  assign mux_864_nl = MUX_s_1_2_2((nor_925_nl), (nor_924_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_124_cse = core_wen & (~ and_dcpl_50)
      & (mux_864_nl);
  assign nor_356_cse = ~(FpMul_8U_23U_lor_32_lpi_1_dfm_st_3 | (~ mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_920_cse = ~((~ (mul_loop_mul_15_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_15_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7);
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_3_cse = MUX_s_1_2_2(mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs_mx0w0,
      mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs, and_dcpl_104);
  assign nor_916_nl = ~((~ IsNaN_8U_23U_1_land_15_lpi_1_dfm_8) | IsNaN_8U_23U_land_15_lpi_1_dfm_10
      | mul_loop_mul_if_land_15_lpi_1_dfm_st_7 | mul_loop_mul_if_land_15_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3));
  assign nor_917_nl = ~((~ IsNaN_8U_23U_1_land_15_lpi_1_dfm_9) | IsNaN_8U_23U_land_15_lpi_1_dfm_11
      | mul_loop_mul_if_land_15_lpi_1_dfm_st_8 | mul_loop_mul_if_land_15_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4));
  assign mux_869_nl = MUX_s_1_2_2((nor_917_nl), (nor_916_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_138_cse = core_wen & (~ and_dcpl_50)
      & (mux_869_nl);
  assign IsNaN_8U_23U_aelse_and_76_cse = core_wen & (~ and_dcpl_50) & (~ mux_870_itm);
  assign nor_910_nl = ~(nor_920_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_15_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_15_lpi_1_dfm_10
      | FpMul_8U_23U_lor_32_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_15_lpi_1_dfm_8
      | mul_loop_mul_if_land_15_lpi_1_dfm_9);
  assign nor_912_nl = ~((FpMul_8U_23U_p_mant_p1_15_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_15_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_15_lpi_1_dfm_10 | FpMul_8U_23U_lor_32_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_15_lpi_1_dfm_8 | mul_loop_mul_if_land_15_lpi_1_dfm_9);
  assign mux_872_nl = MUX_s_1_2_2((nor_912_nl), (nor_910_nl), nor_356_cse);
  assign and_2141_nl = mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_872_nl);
  assign nor_913_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_77_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_15_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_15_lpi_1_dfm_10 | FpMul_8U_23U_lor_32_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_15_lpi_1_dfm_8 | mul_loop_mul_if_land_15_lpi_1_dfm_9);
  assign mux_873_nl = MUX_s_1_2_2((nor_913_nl), (and_2141_nl), nor_53_cse);
  assign nor_914_nl = ~(nor_935_cse | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_15_lpi_1_dfm_11 | mul_loop_mul_if_land_15_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_15_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_15_lpi_1_dfm_9 | FpMul_8U_23U_lor_32_lpi_1_dfm_7 | (~
      FpMul_8U_23U_FpMul_8U_23U_and_77_itm_2));
  assign mux_874_nl = MUX_s_1_2_2((nor_914_nl), (mux_873_nl), or_309_cse);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_14_cse = core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse
      & (mux_874_nl);
  assign and_793_nl = and_dcpl_247 & and_dcpl_85;
  assign and_794_nl = and_dcpl_247 & or_90_cse;
  assign mux_1631_nl = MUX_s_1_2_2(IsNaN_8U_23U_1_land_lpi_1_dfm_9, IsNaN_8U_23U_1_land_lpi_1_dfm_8,
      or_309_cse);
  assign FpMul_8U_23U_p_expo_mux1h_31_itm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_sva_1_mx0w0,
      FpMul_8U_23U_p_expo_sva_1, ({4'b0 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_10}),
      {(and_793_nl) , (and_794_nl) , (mux_1631_nl)});
  assign or_4924_cse = (~ (mul_loop_mul_16_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) |
      mul_loop_mul_16_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  assign or_4912_nl = (or_4924_cse & mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2)
      | FpMul_8U_23U_lor_1_lpi_1_dfm_6;
  assign and_2841_nl = FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_2
      & mul_loop_mul_16_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
      & or_tmp_2114;
  assign mux_1768_nl = MUX_s_1_2_2((and_2841_nl), or_tmp_2114, FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_15_itm);
  assign mux_1769_cse = MUX_s_1_2_2((mux_1768_nl), (or_4912_nl), nor_53_cse);
  assign nor_368_cse = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 |
      (~ mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_898_cse = ~((~ mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs_2) | mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs_st_2);
  assign nor_889_nl = ~(IsNaN_8U_23U_land_lpi_1_dfm_st_7 | (~ IsNaN_8U_23U_1_land_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_lpi_1_dfm_10 | mul_loop_mul_if_land_lpi_1_dfm_st_7 | mul_loop_mul_if_land_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3));
  assign nor_890_nl = ~(IsNaN_8U_23U_land_lpi_1_dfm_st_8 | (~ IsNaN_8U_23U_1_land_lpi_1_dfm_9)
      | IsNaN_8U_23U_land_lpi_1_dfm_11 | mul_loop_mul_if_land_lpi_1_dfm_st_8 | mul_loop_mul_if_land_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4));
  assign mux_889_nl = MUX_s_1_2_2((nor_890_nl), (nor_889_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_126_cse = core_wen & (~ and_dcpl_50)
      & (mux_889_nl);
  assign nor_372_cse = ~(FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | (~ mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_885_cse = ~((~ (mul_loop_mul_16_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_16_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7);
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_1_cse = MUX_s_1_2_2(mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs_mx0w0,
      mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs, and_dcpl_104);
  assign nor_881_nl = ~((~ IsNaN_8U_23U_1_land_lpi_1_dfm_8) | IsNaN_8U_23U_land_lpi_1_dfm_10
      | mul_loop_mul_if_land_lpi_1_dfm_st_7 | mul_loop_mul_if_land_lpi_1_dfm_9 |
      io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 | (~
      main_stage_v_3));
  assign nor_882_nl = ~((~ IsNaN_8U_23U_1_land_lpi_1_dfm_9) | IsNaN_8U_23U_land_lpi_1_dfm_11
      | mul_loop_mul_if_land_lpi_1_dfm_st_8 | mul_loop_mul_if_land_lpi_1_dfm_10 |
      io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~
      main_stage_v_4));
  assign mux_894_nl = MUX_s_1_2_2((nor_882_nl), (nor_881_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_141_cse = core_wen & (~ and_dcpl_50)
      & (mux_894_nl);
  assign IsNaN_8U_23U_aelse_and_78_cse = core_wen & (~ and_dcpl_50) & (~ mux_895_itm);
  assign nor_875_nl = ~(nor_885_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_lpi_1_dfm_10 | FpMul_8U_23U_lor_1_lpi_1_dfm_6
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_lpi_1_dfm_8 | mul_loop_mul_if_land_lpi_1_dfm_9);
  assign nor_877_nl = ~((FpMul_8U_23U_p_mant_p1_sva[47]) | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_lpi_1_dfm_10 | FpMul_8U_23U_lor_1_lpi_1_dfm_6
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_lpi_1_dfm_8 | mul_loop_mul_if_land_lpi_1_dfm_9);
  assign mux_897_nl = MUX_s_1_2_2((nor_877_nl), (nor_875_nl), nor_372_cse);
  assign and_2135_nl = mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_897_nl);
  assign nor_878_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_78_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_lpi_1_dfm_10 | FpMul_8U_23U_lor_1_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_lpi_1_dfm_8 | mul_loop_mul_if_land_lpi_1_dfm_9);
  assign mux_898_nl = MUX_s_1_2_2((nor_878_nl), (and_2135_nl), nor_53_cse);
  assign nor_879_nl = ~(nor_898_cse | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_lpi_1_dfm_11 | mul_loop_mul_if_land_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | mul_loop_mul_if_land_lpi_1_dfm_st_8 | IsNaN_8U_23U_1_land_lpi_1_dfm_9 | FpMul_8U_23U_lor_1_lpi_1_dfm_7
      | (~ FpMul_8U_23U_FpMul_8U_23U_and_78_itm_2));
  assign mux_899_nl = MUX_s_1_2_2((nor_879_nl), (mux_898_nl), or_309_cse);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_15_cse = core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse
      & (mux_899_nl);
  assign or_2278_nl = io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_900_nl = MUX_s_1_2_2((or_2278_nl), or_tmp_608, or_309_cse);
  assign mul_loop_mul_if_aelse_and_64_cse = core_wen & (~ and_dcpl_50) & (~ (mux_900_nl));
  assign nor_872_cse = ~((~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt);
  assign FpMantRNE_48U_24U_else_and_cse = core_wen & (~ or_dcpl_96);
  assign FpMul_8U_23U_p_expo_and_cse = core_wen & (~ or_dcpl_92);
  assign FpMantRNE_48U_24U_else_and_2_cse = core_wen & (~ or_dcpl_103);
  assign FpMul_8U_23U_p_expo_and_1_cse = core_wen & (~ or_dcpl_100);
  assign FpMantRNE_48U_24U_else_carry_and_2_cse = core_wen & (~ or_dcpl_110);
  assign FpMul_8U_23U_p_expo_and_2_cse = core_wen & (~ or_dcpl_107);
  assign FpMantRNE_48U_24U_else_and_6_cse = core_wen & (~ or_dcpl_118);
  assign FpMul_8U_23U_p_expo_and_3_cse = core_wen & (~ or_dcpl_115);
  assign FpMantRNE_48U_24U_else_and_8_cse = core_wen & (~ or_dcpl_125);
  assign FpMul_8U_23U_p_expo_and_4_cse = core_wen & (~ or_dcpl_122);
  assign FpMantRNE_48U_24U_else_and_10_cse = core_wen & (~ or_dcpl_132);
  assign or_2342_cse = (~ mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_23_lpi_1_dfm_st_3;
  assign FpMul_8U_23U_p_expo_and_5_cse = core_wen & (~ or_dcpl_129);
  assign FpMantRNE_48U_24U_else_carry_and_6_cse = core_wen & (~ or_dcpl_139);
  assign FpMul_8U_23U_p_expo_and_6_cse = core_wen & (~ or_dcpl_136);
  assign FpMantRNE_48U_24U_else_and_14_cse = core_wen & (~ or_dcpl_146);
  assign FpMul_8U_23U_p_expo_and_7_cse = core_wen & (~ or_dcpl_143);
  assign FpMantRNE_48U_24U_else_and_16_cse = core_wen & (~ or_dcpl_153);
  assign FpMul_8U_23U_p_expo_and_8_cse = core_wen & (~ or_dcpl_150);
  assign FpMantRNE_48U_24U_else_and_18_cse = core_wen & (~ or_dcpl_160);
  assign or_2386_cse = (~ mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_27_lpi_1_dfm_st_3;
  assign FpMul_8U_23U_p_expo_and_9_cse = core_wen & (~ or_dcpl_157);
  assign FpMantRNE_48U_24U_else_and_20_cse = core_wen & (~ or_dcpl_168);
  assign FpMul_8U_23U_p_expo_and_10_cse = core_wen & (~ or_dcpl_165);
  assign FpMantRNE_48U_24U_else_and_22_cse = core_wen & (~ or_dcpl_176);
  assign FpMul_8U_23U_p_expo_and_11_cse = core_wen & (~ or_dcpl_173);
  assign FpMantRNE_48U_24U_else_and_24_cse = core_wen & (~ or_dcpl_184);
  assign FpMul_8U_23U_p_expo_and_12_cse = core_wen & (~ or_dcpl_181);
  assign FpMantRNE_48U_24U_else_and_26_cse = core_wen & (~ or_dcpl_191);
  assign FpMul_8U_23U_p_expo_and_13_cse = core_wen & (~ or_dcpl_188);
  assign FpMantRNE_48U_24U_else_and_28_cse = core_wen & (~ or_dcpl_198);
  assign FpMul_8U_23U_p_expo_and_14_cse = core_wen & (~ or_dcpl_195);
  assign FpMantRNE_48U_24U_else_carry_and_15_cse = core_wen & (~ or_dcpl_205);
  assign FpMul_8U_23U_p_expo_and_15_cse = core_wen & (~ or_dcpl_202);
  assign mux_987_nl = MUX_s_1_2_2(or_2576_cse, or_tmp_2358, mul_loop_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_988_nl = MUX_s_1_2_2((mux_987_nl), or_2576_cse, reg_FpMul_8U_23U_lor_3_lpi_1_dfm_4_cse);
  assign mux_989_nl = MUX_s_1_2_2(or_tmp_2358, (mux_988_nl), nor_50_cse);
  assign mux_990_nl = MUX_s_1_2_2(or_2576_cse, or_tmp_2358, or_2577_cse);
  assign mux_991_nl = MUX_s_1_2_2((mux_990_nl), (mux_989_nl), nor_53_cse);
  assign or_2453_nl = (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      mul_loop_mul_if_land_1_lpi_1_dfm_st_7 | ((IsNaN_8U_23U_land_1_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_1_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | (~
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_8) | mul_loop_mul_if_land_1_lpi_1_dfm_9) &
      or_4383_cse);
  assign mux_992_nl = MUX_s_1_2_2((or_2453_nl), (mux_991_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_128_cse = core_wen & (~ and_dcpl_50)
      & (~ (mux_992_nl));
  assign mux_994_nl = MUX_s_1_2_2(or_2607_cse, or_tmp_2366, mul_loop_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_995_nl = MUX_s_1_2_2((mux_994_nl), or_2607_cse, reg_FpMul_8U_23U_lor_4_lpi_1_dfm_4_cse);
  assign mux_996_nl = MUX_s_1_2_2(or_tmp_2366, (mux_995_nl), nor_55_cse);
  assign mux_997_nl = MUX_s_1_2_2(or_2607_cse, or_tmp_2366, or_2608_cse);
  assign mux_998_nl = MUX_s_1_2_2((mux_997_nl), (mux_996_nl), nor_53_cse);
  assign or_2461_nl = (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      mul_loop_mul_if_land_2_lpi_1_dfm_st_7 | ((IsNaN_8U_23U_land_2_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_2_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | (~
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_8) | mul_loop_mul_if_land_2_lpi_1_dfm_9) &
      or_4384_cse);
  assign mux_999_nl = MUX_s_1_2_2((or_2461_nl), (mux_998_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_131_cse = core_wen & (~ and_dcpl_50)
      & (~ (mux_999_nl));
  assign mux_1001_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2376, mul_loop_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_1002_nl = MUX_s_1_2_2((mux_1001_nl), (~ main_stage_v_2), reg_FpMul_8U_23U_lor_5_lpi_1_dfm_4_cse);
  assign mux_1003_nl = MUX_s_1_2_2(or_tmp_2376, (mux_1002_nl), nor_59_cse);
  assign mux_1004_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2376, or_2631_cse);
  assign mux_1005_nl = MUX_s_1_2_2((mux_1004_nl), (mux_1003_nl), nor_53_cse);
  assign mux_1006_nl = MUX_s_1_2_2((mux_1005_nl), or_tmp_2376, or_tmp_134);
  assign nor_838_nl = ~(or_tmp_1088 | (~(mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & main_stage_v_3)));
  assign or_2467_nl = io_read_cfg_mul_bypass_rsc_svs_7 | (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_8)
      | mul_loop_mul_if_land_3_lpi_1_dfm_9;
  assign mux_1007_nl = MUX_s_1_2_2(main_stage_v_3, (nor_838_nl), or_2467_nl);
  assign mux_1008_nl = MUX_s_1_2_2((mux_1007_nl), (~ (mux_1006_nl)), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_134_cse = core_wen & (~ and_dcpl_50)
      & (mux_1008_nl);
  assign mux_1010_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2384, mul_loop_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_1011_nl = MUX_s_1_2_2((mux_1010_nl), (~ main_stage_v_2), reg_FpMul_8U_23U_lor_6_lpi_1_dfm_4_cse);
  assign mux_1012_nl = MUX_s_1_2_2(or_tmp_2384, (mux_1011_nl), nor_64_cse);
  assign mux_1013_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2384, or_378_cse);
  assign mux_1014_nl = MUX_s_1_2_2((mux_1013_nl), (mux_1012_nl), nor_53_cse);
  assign mux_1015_nl = MUX_s_1_2_2((mux_1014_nl), or_tmp_2384, or_tmp_141);
  assign nor_837_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_4_lpi_1_dfm_st_7
      | FpMul_8U_23U_lor_21_lpi_1_dfm_st_3 | (~(mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & main_stage_v_3)));
  assign or_2475_nl = io_read_cfg_mul_bypass_rsc_svs_7 | (~ IsNaN_8U_23U_1_land_4_lpi_1_dfm_8)
      | mul_loop_mul_if_land_4_lpi_1_dfm_9;
  assign mux_1016_nl = MUX_s_1_2_2(main_stage_v_3, (nor_837_nl), or_2475_nl);
  assign mux_1017_nl = MUX_s_1_2_2((mux_1016_nl), (~ (mux_1015_nl)), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_137_cse = core_wen & (~ and_dcpl_50)
      & (mux_1017_nl);
  assign mux_1019_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2392, mul_loop_mul_5_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_1020_nl = MUX_s_1_2_2((mux_1019_nl), (~ main_stage_v_2), reg_FpMul_8U_23U_lor_7_lpi_1_dfm_4_cse);
  assign mux_1021_nl = MUX_s_1_2_2(or_tmp_2392, (mux_1020_nl), nor_69_cse);
  assign mux_1022_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2392, or_2675_cse);
  assign mux_1023_nl = MUX_s_1_2_2((mux_1022_nl), (mux_1021_nl), nor_53_cse);
  assign mux_1024_nl = MUX_s_1_2_2((mux_1023_nl), or_tmp_2392, or_tmp_147);
  assign nor_836_nl = ~(or_tmp_321 | (~(mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & main_stage_v_3)));
  assign or_2483_nl = io_read_cfg_mul_bypass_rsc_svs_7 | (~ IsNaN_8U_23U_1_land_5_lpi_1_dfm_8)
      | mul_loop_mul_if_land_5_lpi_1_dfm_9;
  assign mux_1025_nl = MUX_s_1_2_2(main_stage_v_3, (nor_836_nl), or_2483_nl);
  assign mux_1026_nl = MUX_s_1_2_2((mux_1025_nl), (~ (mux_1024_nl)), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_140_cse = core_wen & (~ and_dcpl_50)
      & (mux_1026_nl);
  assign mux_1028_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2400, mul_loop_mul_6_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_1029_nl = MUX_s_1_2_2((mux_1028_nl), (~ main_stage_v_2), reg_FpMul_8U_23U_lor_8_lpi_1_dfm_4_cse);
  assign mux_1030_nl = MUX_s_1_2_2(or_tmp_2400, (mux_1029_nl), nor_73_cse);
  assign mux_1031_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2400, or_430_cse);
  assign mux_1032_nl = MUX_s_1_2_2((mux_1031_nl), (mux_1030_nl), nor_53_cse);
  assign mux_1033_nl = MUX_s_1_2_2((mux_1032_nl), or_tmp_2400, or_tmp_151);
  assign nor_835_nl = ~(or_tmp_1333 | (~(mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & main_stage_v_3)));
  assign or_2491_nl = io_read_cfg_mul_bypass_rsc_svs_7 | (~ IsNaN_8U_23U_1_land_6_lpi_1_dfm_8)
      | mul_loop_mul_if_land_6_lpi_1_dfm_9;
  assign mux_1034_nl = MUX_s_1_2_2(main_stage_v_3, (nor_835_nl), or_2491_nl);
  assign mux_1035_nl = MUX_s_1_2_2((mux_1034_nl), (~ (mux_1033_nl)), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_143_cse = core_wen & (~ and_dcpl_50)
      & (mux_1035_nl);
  assign mux_1037_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2408, mul_loop_mul_7_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_1038_nl = MUX_s_1_2_2((mux_1037_nl), (~ main_stage_v_2), reg_FpMul_8U_23U_lor_9_lpi_1_dfm_4_cse);
  assign mux_1039_nl = MUX_s_1_2_2(or_tmp_2408, (mux_1038_nl), nor_78_cse);
  assign mux_1040_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2408, or_453_cse);
  assign mux_1041_nl = MUX_s_1_2_2((mux_1040_nl), (mux_1039_nl), nor_53_cse);
  assign mux_1042_nl = MUX_s_1_2_2((mux_1041_nl), or_tmp_2408, or_tmp_155);
  assign nor_834_nl = ~(or_tmp_1415 | (~(mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & main_stage_v_3)));
  assign or_2499_nl = io_read_cfg_mul_bypass_rsc_svs_7 | (~ IsNaN_8U_23U_1_land_7_lpi_1_dfm_8)
      | mul_loop_mul_if_land_7_lpi_1_dfm_9;
  assign mux_1043_nl = MUX_s_1_2_2(main_stage_v_3, (nor_834_nl), or_2499_nl);
  assign mux_1044_nl = MUX_s_1_2_2((mux_1043_nl), (~ (mux_1042_nl)), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_146_cse = core_wen & (~ and_dcpl_50)
      & (mux_1044_nl);
  assign mux_1046_nl = MUX_s_1_2_2(or_2721_cse, or_tmp_2414, mul_loop_mul_8_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_1047_nl = MUX_s_1_2_2((mux_1046_nl), or_2721_cse, reg_FpMul_8U_23U_lor_10_lpi_1_dfm_4_cse);
  assign mux_1048_nl = MUX_s_1_2_2(or_tmp_2414, (mux_1047_nl), nor_83_cse);
  assign mux_1049_nl = MUX_s_1_2_2(or_2721_cse, or_tmp_2414, or_2722_cse);
  assign mux_1050_nl = MUX_s_1_2_2((mux_1049_nl), (mux_1048_nl), nor_53_cse);
  assign or_2509_nl = (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      mul_loop_mul_if_land_8_lpi_1_dfm_st_7 | ((IsNaN_8U_23U_land_8_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_8_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | (~
      IsNaN_8U_23U_1_land_8_lpi_1_dfm_8) | mul_loop_mul_if_land_8_lpi_1_dfm_9) &
      or_4390_cse);
  assign mux_1051_nl = MUX_s_1_2_2((or_2509_nl), (mux_1050_nl), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_149_cse = core_wen & (~ and_dcpl_50)
      & (~ (mux_1051_nl));
  assign mux_1053_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2424, mul_loop_mul_9_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_1054_nl = MUX_s_1_2_2((mux_1053_nl), (~ main_stage_v_2), reg_FpMul_8U_23U_lor_11_lpi_1_dfm_4_cse);
  assign mux_1055_nl = MUX_s_1_2_2(or_tmp_2424, (mux_1054_nl), nor_87_cse);
  assign mux_1056_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2424, or_2745_cse);
  assign mux_1057_nl = MUX_s_1_2_2((mux_1056_nl), (mux_1055_nl), nor_53_cse);
  assign mux_1058_nl = MUX_s_1_2_2((mux_1057_nl), or_tmp_2424, or_tmp_167);
  assign nor_833_nl = ~(or_tmp_424 | (~(mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & main_stage_v_3)));
  assign or_2515_nl = io_read_cfg_mul_bypass_rsc_svs_7 | (~ IsNaN_8U_23U_1_land_9_lpi_1_dfm_8)
      | mul_loop_mul_if_land_9_lpi_1_dfm_9;
  assign mux_1059_nl = MUX_s_1_2_2(main_stage_v_3, (nor_833_nl), or_2515_nl);
  assign mux_1060_nl = MUX_s_1_2_2((mux_1059_nl), (~ (mux_1058_nl)), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_152_cse = core_wen & (~ and_dcpl_50)
      & (mux_1060_nl);
  assign mux_1062_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2432, mul_loop_mul_10_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_1063_nl = MUX_s_1_2_2((mux_1062_nl), (~ main_stage_v_2), reg_FpMul_8U_23U_lor_12_lpi_1_dfm_4_cse);
  assign mux_1064_nl = MUX_s_1_2_2(or_tmp_2432, (mux_1063_nl), nor_91_cse);
  assign mux_1065_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2432, or_533_cse);
  assign mux_1066_nl = MUX_s_1_2_2((mux_1065_nl), (mux_1064_nl), nor_53_cse);
  assign mux_1067_nl = MUX_s_1_2_2((mux_1066_nl), or_tmp_2432, or_tmp_171);
  assign nor_832_nl = ~(or_tmp_453 | (~(mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & main_stage_v_3)));
  assign or_2523_nl = io_read_cfg_mul_bypass_rsc_svs_7 | (~ IsNaN_8U_23U_1_land_10_lpi_1_dfm_8)
      | mul_loop_mul_if_land_10_lpi_1_dfm_9;
  assign mux_1068_nl = MUX_s_1_2_2(main_stage_v_3, (nor_832_nl), or_2523_nl);
  assign mux_1069_nl = MUX_s_1_2_2((mux_1068_nl), (~ (mux_1067_nl)), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_155_cse = core_wen & (~ and_dcpl_50)
      & (mux_1069_nl);
  assign mux_1071_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2440, mul_loop_mul_11_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_1072_nl = MUX_s_1_2_2((mux_1071_nl), (~ main_stage_v_2), reg_FpMul_8U_23U_lor_13_lpi_1_dfm_4_cse);
  assign mux_1073_nl = MUX_s_1_2_2(or_tmp_2440, (mux_1072_nl), nor_95_cse);
  assign mux_1074_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2440, or_562_cse);
  assign mux_1075_nl = MUX_s_1_2_2((mux_1074_nl), (mux_1073_nl), nor_53_cse);
  assign mux_1076_nl = MUX_s_1_2_2((mux_1075_nl), or_tmp_2440, or_tmp_175);
  assign nor_831_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_11_lpi_1_dfm_st_7
      | FpMul_8U_23U_lor_28_lpi_1_dfm_st_3 | (~(mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & main_stage_v_3)));
  assign or_2531_nl = io_read_cfg_mul_bypass_rsc_svs_7 | (~ IsNaN_8U_23U_1_land_11_lpi_1_dfm_8)
      | mul_loop_mul_if_land_11_lpi_1_dfm_9;
  assign mux_1077_nl = MUX_s_1_2_2(main_stage_v_3, (nor_831_nl), or_2531_nl);
  assign mux_1078_nl = MUX_s_1_2_2((mux_1077_nl), (~ (mux_1076_nl)), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_158_cse = core_wen & (~ and_dcpl_50)
      & (mux_1078_nl);
  assign mux_1080_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2448, mul_loop_mul_12_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_1081_nl = MUX_s_1_2_2((mux_1080_nl), (~ main_stage_v_2), reg_FpMul_8U_23U_lor_14_lpi_1_dfm_4_cse);
  assign mux_1082_nl = MUX_s_1_2_2(or_tmp_2448, (mux_1081_nl), nor_100_cse);
  assign mux_1083_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2448, or_585_cse);
  assign mux_1084_nl = MUX_s_1_2_2((mux_1083_nl), (mux_1082_nl), nor_53_cse);
  assign mux_1085_nl = MUX_s_1_2_2((mux_1084_nl), or_tmp_2448, or_tmp_179);
  assign nor_830_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_12_lpi_1_dfm_st_7
      | FpMul_8U_23U_lor_29_lpi_1_dfm_st_3 | (~(mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & main_stage_v_3)));
  assign or_2539_nl = io_read_cfg_mul_bypass_rsc_svs_7 | (~ IsNaN_8U_23U_1_land_12_lpi_1_dfm_8)
      | mul_loop_mul_if_land_12_lpi_1_dfm_9;
  assign mux_1086_nl = MUX_s_1_2_2(main_stage_v_3, (nor_830_nl), or_2539_nl);
  assign mux_1087_nl = MUX_s_1_2_2((mux_1086_nl), (~ (mux_1085_nl)), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_161_cse = core_wen & (~ and_dcpl_50)
      & (mux_1087_nl);
  assign mux_1089_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2456, mul_loop_mul_13_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_1090_nl = MUX_s_1_2_2((mux_1089_nl), (~ main_stage_v_2), reg_FpMul_8U_23U_lor_15_lpi_1_dfm_4_cse);
  assign mux_1091_nl = MUX_s_1_2_2(or_tmp_2456, (mux_1090_nl), nor_105_cse);
  assign mux_1092_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2456, or_2798_cse);
  assign mux_1093_nl = MUX_s_1_2_2((mux_1092_nl), (mux_1091_nl), nor_53_cse);
  assign mux_1094_nl = MUX_s_1_2_2((mux_1093_nl), or_tmp_2456, or_tmp_185);
  assign nor_829_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_13_lpi_1_dfm_st_7
      | FpMul_8U_23U_lor_30_lpi_1_dfm_st_3 | (~(mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & main_stage_v_3)));
  assign or_2547_nl = io_read_cfg_mul_bypass_rsc_svs_7 | (~ IsNaN_8U_23U_1_land_13_lpi_1_dfm_8)
      | mul_loop_mul_if_land_13_lpi_1_dfm_9;
  assign mux_1095_nl = MUX_s_1_2_2(main_stage_v_3, (nor_829_nl), or_2547_nl);
  assign mux_1096_nl = MUX_s_1_2_2((mux_1095_nl), (~ (mux_1094_nl)), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_164_cse = core_wen & (~ and_dcpl_50)
      & (mux_1096_nl);
  assign mux_1098_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2464, mul_loop_mul_14_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_1099_nl = MUX_s_1_2_2((mux_1098_nl), (~ main_stage_v_2), reg_FpMul_8U_23U_lor_16_lpi_1_dfm_4_cse);
  assign mux_1100_nl = MUX_s_1_2_2(or_tmp_2464, (mux_1099_nl), nor_110_cse);
  assign mux_1101_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2464, or_631_cse);
  assign mux_1102_nl = MUX_s_1_2_2((mux_1101_nl), (mux_1100_nl), nor_53_cse);
  assign mux_1103_nl = MUX_s_1_2_2((mux_1102_nl), or_tmp_2464, or_tmp_189);
  assign nor_828_nl = ~(or_tmp_1985 | (~(mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & main_stage_v_3)));
  assign or_2555_nl = io_read_cfg_mul_bypass_rsc_svs_7 | (~ IsNaN_8U_23U_1_land_14_lpi_1_dfm_8)
      | mul_loop_mul_if_land_14_lpi_1_dfm_9;
  assign mux_1104_nl = MUX_s_1_2_2(main_stage_v_3, (nor_828_nl), or_2555_nl);
  assign mux_1105_nl = MUX_s_1_2_2((mux_1104_nl), (~ (mux_1103_nl)), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_167_cse = core_wen & (~ and_dcpl_50)
      & (mux_1105_nl);
  assign mux_1107_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2472, mul_loop_mul_15_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_1108_nl = MUX_s_1_2_2((mux_1107_nl), (~ main_stage_v_2), reg_FpMul_8U_23U_lor_17_lpi_1_dfm_4_cse);
  assign mux_1109_nl = MUX_s_1_2_2(or_tmp_2472, (mux_1108_nl), nor_115_cse);
  assign mux_1110_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2472, or_2834_cse);
  assign mux_1111_nl = MUX_s_1_2_2((mux_1110_nl), (mux_1109_nl), nor_53_cse);
  assign mux_1112_nl = MUX_s_1_2_2((mux_1111_nl), or_tmp_2472, or_tmp_195);
  assign nor_827_nl = ~(or_tmp_2065 | (~(mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & main_stage_v_3)));
  assign or_2563_nl = io_read_cfg_mul_bypass_rsc_svs_7 | (~ IsNaN_8U_23U_1_land_15_lpi_1_dfm_8)
      | mul_loop_mul_if_land_15_lpi_1_dfm_9;
  assign mux_1113_nl = MUX_s_1_2_2(main_stage_v_3, (nor_827_nl), or_2563_nl);
  assign mux_1114_nl = MUX_s_1_2_2((mux_1113_nl), (~ (mux_1112_nl)), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_170_cse = core_wen & (~ and_dcpl_50)
      & (mux_1114_nl);
  assign mux_1115_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2480, or_tmp_201);
  assign or_2570_nl = mul_loop_mul_16_FpMul_8U_23U_oelse_1_acc_itm_9_1 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_lpi_1_dfm_st_6;
  assign mux_1116_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2480, or_2570_nl);
  assign mux_1117_nl = MUX_s_1_2_2((mux_1116_nl), (mux_1115_nl), reg_FpMul_8U_23U_lor_lpi_1_dfm_4_cse);
  assign mux_1118_nl = MUX_s_1_2_2(or_tmp_2480, (mux_1117_nl), nor_120_cse);
  assign or_2571_nl = (~ mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_1_lpi_1_dfm_st | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_lpi_1_dfm_st_6;
  assign mux_1119_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_2480, or_2571_nl);
  assign mux_1120_nl = MUX_s_1_2_2((mux_1119_nl), (mux_1118_nl), nor_53_cse);
  assign nor_826_nl = ~(or_tmp_597 | (~(mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & main_stage_v_3)));
  assign or_2572_nl = io_read_cfg_mul_bypass_rsc_svs_7 | (~ IsNaN_8U_23U_1_land_lpi_1_dfm_8)
      | mul_loop_mul_if_land_lpi_1_dfm_9;
  assign mux_1121_nl = MUX_s_1_2_2(main_stage_v_3, (nor_826_nl), or_2572_nl);
  assign mux_1122_nl = MUX_s_1_2_2((mux_1121_nl), (~ (mux_1120_nl)), or_309_cse);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_173_cse = core_wen & (~ and_dcpl_50)
      & (mux_1122_nl);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_144_cse = core_wen & (and_dcpl_262
      | and_dcpl_266 | and_dcpl_102) & mux_tmp_148;
  assign IsZero_8U_23U_aelse_and_cse = core_wen & (~ and_dcpl_50);
  assign nor_825_nl = ~(mul_loop_mul_1_FpMul_8U_23U_else_2_if_acc_itm_8_1 | (~ and_tmp_86));
  assign mux_1680_itm = MUX_s_1_2_2((nor_825_nl), and_tmp_86, mul_loop_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign or_2577_cse = (~ mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_18_lpi_1_dfm_st;
  assign or_2575_cse = (~ cfg_mul_src_1_sva_st_1) | chn_mul_op_rsci_bawt;
  assign and_2130_cse = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1)
      & (~ mul_loop_mul_if_land_1_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt;
  assign or_2576_cse = (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 |
      mul_loop_mul_if_land_1_lpi_1_dfm_st_6;
  assign FpMul_8U_23U_else_2_if_and_cse = core_wen & (~ (fsm_output[0]));
  assign nor_821_cse = ~(mul_loop_mul_if_land_1_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_147_cse = core_wen & (and_dcpl_277
      | and_dcpl_281 | and_dcpl_108) & mux_tmp_148;
  assign nor_818_nl = ~(mul_loop_mul_2_FpMul_8U_23U_else_2_if_acc_itm_8_1 | (~ and_tmp_90));
  assign mux_1681_itm = MUX_s_1_2_2((nor_818_nl), and_tmp_90, mul_loop_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign or_2608_cse = (~ mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_19_lpi_1_dfm_st;
  assign or_2607_cse = (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 |
      mul_loop_mul_if_land_2_lpi_1_dfm_st_6;
  assign or_2628_cse = mul_loop_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_4_lpi_1_dfm_4_cse;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_150_cse = core_wen & (and_dcpl_292
      | and_dcpl_296 | and_dcpl_112) & mux_tmp_148;
  assign nor_816_nl = ~(mul_loop_mul_3_FpMul_8U_23U_else_2_if_acc_itm_8_1 | (~ and_tmp_95));
  assign mux_1682_itm = MUX_s_1_2_2((nor_816_nl), and_tmp_95, mul_loop_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign or_2631_cse = (~ mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_20_lpi_1_dfm_st;
  assign or_2630_cse = (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 |
      mul_loop_mul_if_land_3_lpi_1_dfm_st_6;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_153_cse = core_wen & (and_dcpl_307
      | and_dcpl_311 | and_dcpl_116) & mux_tmp_148;
  assign IsZero_8U_23U_1_aelse_and_cse = core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse;
  assign or_2664_cse = mul_loop_mul_if_land_4_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_156_cse = core_wen & (and_dcpl_322
      | and_dcpl_326 | and_dcpl_120) & mux_tmp_148;
  assign nor_806_nl = ~(mul_loop_mul_5_FpMul_8U_23U_else_2_if_acc_itm_8_1 | (~ and_tmp_99));
  assign mux_1683_itm = MUX_s_1_2_2((nor_806_nl), and_tmp_99, mul_loop_mul_5_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign or_2675_cse = (~ mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_22_lpi_1_dfm_st;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_159_cse = core_wen & (and_dcpl_337
      | and_dcpl_341 | and_dcpl_124) & mux_tmp_148;
  assign or_2698_cse = mul_loop_mul_if_land_6_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_162_cse = core_wen & (and_dcpl_352
      | and_dcpl_356 | and_dcpl_128) & mux_tmp_148;
  assign or_2711_cse = mul_loop_mul_if_land_7_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_165_cse = core_wen & (and_dcpl_367
      | and_dcpl_371 | and_dcpl_132) & mux_tmp_148;
  assign nor_798_nl = ~(mul_loop_mul_8_FpMul_8U_23U_else_2_if_acc_itm_8_1 | (~ and_tmp_104));
  assign mux_1684_itm = MUX_s_1_2_2((nor_798_nl), and_tmp_104, mul_loop_mul_8_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign or_2722_cse = (~ mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_25_lpi_1_dfm_st;
  assign or_2721_cse = (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 |
      mul_loop_mul_if_land_8_lpi_1_dfm_st_6;
  assign or_2742_cse = mul_loop_mul_8_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_10_lpi_1_dfm_4_cse;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_168_cse = core_wen & (and_dcpl_382
      | and_dcpl_386 | and_dcpl_136) & mux_tmp_148;
  assign nor_796_nl = ~(mul_loop_mul_9_FpMul_8U_23U_else_2_if_acc_itm_8_1 | (~ and_tmp_109));
  assign mux_1685_itm = MUX_s_1_2_2((nor_796_nl), and_tmp_109, mul_loop_mul_9_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign or_2745_cse = (~ mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_26_lpi_1_dfm_st;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_171_cse = core_wen & (and_dcpl_397
      | and_dcpl_401 | and_dcpl_140) & mux_tmp_148;
  assign or_2767_cse = mul_loop_mul_if_land_10_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_174_cse = core_wen & (and_dcpl_412
      | and_dcpl_416 | and_dcpl_144) & mux_tmp_148;
  assign or_2774_cse = mul_loop_mul_if_land_11_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_177_cse = core_wen & (and_dcpl_427
      | and_dcpl_431 | and_dcpl_148) & mux_tmp_148;
  assign or_2787_cse = mul_loop_mul_if_land_12_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_180_cse = core_wen & (and_dcpl_442
      | and_dcpl_446 | and_dcpl_152) & mux_tmp_148;
  assign nor_788_nl = ~(mul_loop_mul_13_FpMul_8U_23U_else_2_if_acc_itm_8_1 | (~ and_tmp_114));
  assign mux_1686_itm = MUX_s_1_2_2((nor_788_nl), and_tmp_114, mul_loop_mul_13_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign or_2798_cse = (~ mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_30_lpi_1_dfm_st;
  assign or_2797_cse = (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 |
      mul_loop_mul_if_land_13_lpi_1_dfm_st_6;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_183_cse = core_wen & (and_dcpl_457
      | and_dcpl_461 | and_dcpl_156) & mux_tmp_148;
  assign or_2823_cse = mul_loop_mul_if_land_14_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_186_cse = core_wen & (and_dcpl_472
      | and_dcpl_476 | and_dcpl_160) & mux_tmp_148;
  assign nor_783_nl = ~(mul_loop_mul_15_FpMul_8U_23U_else_2_if_acc_itm_8_1 | (~ and_tmp_119));
  assign mux_1687_itm = MUX_s_1_2_2((nor_783_nl), and_tmp_119, mul_loop_mul_15_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign or_2834_cse = (~ mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_32_lpi_1_dfm_st;
  assign or_2833_cse = (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 |
      mul_loop_mul_if_land_15_lpi_1_dfm_st_6;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_189_cse = core_wen & (and_dcpl_487
      | and_dcpl_491 | and_dcpl_164) & mux_tmp_148;
  assign nor_776_nl = ~(mul_loop_mul_16_FpMul_8U_23U_else_2_if_acc_itm_8_1 | (~ and_tmp_123));
  assign mux_1688_itm = MUX_s_1_2_2((nor_776_nl), and_tmp_123, mul_loop_mul_16_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign or_2865_cse = (~ mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_1_lpi_1_dfm_st;
  assign or_2864_cse = (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 |
      mul_loop_mul_if_land_lpi_1_dfm_st_6;
  assign or_2885_cse = mul_loop_mul_16_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_lpi_1_dfm_4_cse;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_cse = core_wen & (~ or_dcpl_373);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_3_cse = core_wen & (~(or_dcpl_27
      | or_tmp_10 | mul_loop_mul_if_land_2_lpi_1_dfm_st_5 | or_dcpl_369));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_6_cse = core_wen & (~(or_dcpl_27
      | or_tmp_10 | mul_loop_mul_if_land_3_lpi_1_dfm_st_5 | or_dcpl_369));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_9_cse = core_wen & (~(or_dcpl_385
      | or_dcpl_382 | mul_loop_mul_if_land_4_lpi_1_dfm_st_5 | (cfg_precision!=2'b10)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_12_cse = core_wen & (~(or_dcpl_27
      | or_tmp_10 | mul_loop_mul_if_land_5_lpi_1_dfm_st_5 | or_dcpl_369));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_15_cse = core_wen & (~(or_dcpl_385
      | or_dcpl_382 | mul_loop_mul_if_land_6_lpi_1_dfm_st_5 | (cfg_precision!=2'b10)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_18_cse = core_wen & (~(or_dcpl_385
      | or_dcpl_382 | mul_loop_mul_if_land_7_lpi_1_dfm_st_5 | (cfg_precision!=2'b10)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_21_cse = core_wen & (~(or_dcpl_27
      | or_tmp_10 | mul_loop_mul_if_land_8_lpi_1_dfm_st_5 | or_dcpl_369));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_24_cse = core_wen & (~(or_dcpl_27
      | or_tmp_10 | mul_loop_mul_if_land_9_lpi_1_dfm_st_5 | or_dcpl_369));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_27_cse = core_wen & (~(or_dcpl_385
      | or_dcpl_382 | mul_loop_mul_if_land_10_lpi_1_dfm_st_5 | (cfg_precision!=2'b10)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_30_cse = core_wen & (~(or_dcpl_385
      | or_dcpl_382 | mul_loop_mul_if_land_11_lpi_1_dfm_st_5 | (cfg_precision!=2'b10)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_33_cse = core_wen & (~(or_dcpl_385
      | or_dcpl_382 | mul_loop_mul_if_land_12_lpi_1_dfm_st_5 | (cfg_precision!=2'b10)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_36_cse = core_wen & (~(or_dcpl_27
      | or_tmp_10 | mul_loop_mul_if_land_13_lpi_1_dfm_st_5 | or_dcpl_369));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_39_cse = core_wen & (~(or_dcpl_385
      | or_dcpl_382 | mul_loop_mul_if_land_14_lpi_1_dfm_st_5 | (cfg_precision!=2'b10)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_42_cse = core_wen & (~(or_dcpl_27
      | or_tmp_10 | mul_loop_mul_if_land_15_lpi_1_dfm_st_5 | or_dcpl_369));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_45_cse = core_wen & (~(or_dcpl_27
      | or_tmp_10 | mul_loop_mul_if_land_lpi_1_dfm_st_5 | or_dcpl_369));
  assign or_4649_cse = io_read_cfg_mul_bypass_rsc_svs_st_1 | (~ cfg_mul_src_1_sva_st_1)
      | chn_mul_op_rsci_bawt;
  assign mul_loop_mul_if_aelse_and_cse = core_wen & (~(and_dcpl_53 | and_dcpl_50
      | cfg_mul_bypass_rsci_d | or_90_cse | (~ chn_mul_in_rsci_bawt) | (fsm_output[0])));
  assign MulIn_data_and_3_cse = core_wen & (~ or_dcpl_46) & mux_tmp_1422;
  assign IsZero_8U_23U_aelse_and_48_cse = core_wen & ((and_dcpl_7 & or_70_cse & and_dcpl_494)
      | and_dcpl_497) & mux_tmp_1422;
  assign IsZero_8U_23U_aelse_and_49_cse = core_wen & ((and_dcpl_7 & or_75_cse & and_dcpl_494)
      | and_dcpl_500) & mux_tmp_1422;
  assign IsZero_8U_23U_aelse_and_50_cse = core_wen & ((and_dcpl_7 & or_76_cse & and_dcpl_494)
      | and_dcpl_503) & mux_tmp_1422;
  assign IsZero_8U_23U_aelse_and_51_cse = core_wen & ((and_dcpl_7 & or_77_cse & and_dcpl_494)
      | and_dcpl_506) & mux_tmp_1422;
  assign IsZero_8U_23U_aelse_and_52_cse = core_wen & ((and_dcpl_7 & or_78_cse & and_dcpl_494)
      | and_dcpl_509) & mux_tmp_1422;
  assign IsZero_8U_23U_aelse_and_53_cse = core_wen & ((and_dcpl_7 & or_79_cse & and_dcpl_494)
      | and_dcpl_512) & mux_tmp_1422;
  assign IsZero_8U_23U_aelse_and_54_cse = core_wen & ((and_dcpl_7 & or_80_cse & and_dcpl_494)
      | and_dcpl_515) & mux_tmp_1422;
  assign IsZero_8U_23U_aelse_and_55_cse = core_wen & ((and_dcpl_7 & or_81_cse & and_dcpl_494)
      | and_dcpl_518) & mux_tmp_1422;
  assign IsZero_8U_23U_aelse_and_56_cse = core_wen & ((and_dcpl_7 & or_82_cse & and_dcpl_494)
      | and_dcpl_521) & mux_tmp_1422;
  assign IsZero_8U_23U_aelse_and_57_cse = core_wen & ((and_dcpl_7 & or_83_cse & and_dcpl_494)
      | and_dcpl_524) & mux_tmp_1422;
  assign IsZero_8U_23U_aelse_and_58_cse = core_wen & ((and_dcpl_7 & or_84_cse & and_dcpl_494)
      | and_dcpl_527) & mux_tmp_1422;
  assign IsZero_8U_23U_aelse_and_59_cse = core_wen & ((and_dcpl_7 & or_85_cse & and_dcpl_494)
      | and_dcpl_530) & mux_tmp_1422;
  assign IsZero_8U_23U_aelse_and_60_cse = core_wen & ((and_dcpl_7 & or_86_cse & and_dcpl_494)
      | and_dcpl_533) & mux_tmp_1422;
  assign IsZero_8U_23U_aelse_and_61_cse = core_wen & ((and_dcpl_7 & or_87_cse & and_dcpl_494)
      | and_dcpl_536) & mux_tmp_1422;
  assign IsZero_8U_23U_aelse_and_62_cse = core_wen & ((and_dcpl_7 & or_88_cse & and_dcpl_494)
      | and_dcpl_539) & mux_tmp_1422;
  assign IsZero_8U_23U_aelse_and_63_cse = core_wen & ((and_dcpl_7 & or_89_cse & and_dcpl_494)
      | and_dcpl_542) & mux_tmp_1422;
  assign and_1108_rgt = and_dcpl_546 & IsNaN_8U_23U_land_lpi_1_dfm_9 & (cfg_precision==2'b10);
  assign and_1111_rgt = and_dcpl_546 & (~ IsNaN_8U_23U_land_lpi_1_dfm_9) & (cfg_precision==2'b10);
  assign and_1112_rgt = (or_tmp_201 | or_90_cse) & or_309_cse;
  assign and_1117_rgt = and_dcpl_555 & IsNaN_8U_23U_land_15_lpi_1_dfm_9 & (cfg_precision==2'b10);
  assign and_1120_rgt = and_dcpl_555 & (~ IsNaN_8U_23U_land_15_lpi_1_dfm_9) & (cfg_precision==2'b10);
  assign and_1121_rgt = (or_tmp_195 | or_90_cse) & or_309_cse;
  assign and_1126_rgt = and_dcpl_564 & IsNaN_8U_23U_land_14_lpi_1_dfm_9 & (cfg_precision==2'b10);
  assign and_1129_rgt = and_dcpl_564 & (~ IsNaN_8U_23U_land_14_lpi_1_dfm_9) & (cfg_precision==2'b10);
  assign and_1130_rgt = (or_tmp_189 | or_90_cse) & or_309_cse;
  assign and_1135_rgt = and_dcpl_573 & IsNaN_8U_23U_land_13_lpi_1_dfm_9 & (cfg_precision==2'b10);
  assign and_1138_rgt = and_dcpl_573 & (~ IsNaN_8U_23U_land_13_lpi_1_dfm_9) & (cfg_precision==2'b10);
  assign and_1139_rgt = (or_tmp_185 | or_90_cse) & or_309_cse;
  assign and_1144_rgt = and_dcpl_582 & IsNaN_8U_23U_land_12_lpi_1_dfm_9 & (cfg_precision==2'b10);
  assign and_1147_rgt = and_dcpl_582 & (~ IsNaN_8U_23U_land_12_lpi_1_dfm_9) & (cfg_precision==2'b10);
  assign and_1148_rgt = (or_tmp_179 | or_90_cse) & or_309_cse;
  assign and_1153_rgt = and_dcpl_591 & IsNaN_8U_23U_land_11_lpi_1_dfm_9 & (cfg_precision==2'b10);
  assign and_1156_rgt = and_dcpl_591 & (~ IsNaN_8U_23U_land_11_lpi_1_dfm_9) & (cfg_precision==2'b10);
  assign and_1157_rgt = (or_tmp_175 | or_90_cse) & or_309_cse;
  assign and_1162_rgt = and_dcpl_600 & IsNaN_8U_23U_land_10_lpi_1_dfm_9 & (cfg_precision==2'b10);
  assign and_1165_rgt = and_dcpl_600 & (~ IsNaN_8U_23U_land_10_lpi_1_dfm_9) & (cfg_precision==2'b10);
  assign and_1166_rgt = (or_tmp_171 | or_90_cse) & or_309_cse;
  assign and_1171_rgt = and_dcpl_609 & IsNaN_8U_23U_land_9_lpi_1_dfm_9 & (cfg_precision==2'b10);
  assign and_1174_rgt = and_dcpl_609 & (~ IsNaN_8U_23U_land_9_lpi_1_dfm_9) & (cfg_precision==2'b10);
  assign and_1175_rgt = (or_tmp_167 | or_90_cse) & or_309_cse;
  assign and_1180_rgt = and_dcpl_618 & IsNaN_8U_23U_land_8_lpi_1_dfm_9 & (cfg_precision==2'b10);
  assign and_1183_rgt = and_dcpl_618 & (~ IsNaN_8U_23U_land_8_lpi_1_dfm_9) & (cfg_precision==2'b10);
  assign and_1184_rgt = (or_tmp_161 | or_90_cse) & or_309_cse;
  assign and_1189_rgt = and_dcpl_627 & IsNaN_8U_23U_land_7_lpi_1_dfm_9 & (cfg_precision==2'b10);
  assign and_1192_rgt = and_dcpl_627 & (~ IsNaN_8U_23U_land_7_lpi_1_dfm_9) & (cfg_precision==2'b10);
  assign and_1193_rgt = (or_tmp_155 | or_90_cse) & or_309_cse;
  assign and_1198_rgt = and_dcpl_636 & IsNaN_8U_23U_land_6_lpi_1_dfm_9 & (cfg_precision==2'b10);
  assign and_1201_rgt = and_dcpl_636 & (~ IsNaN_8U_23U_land_6_lpi_1_dfm_9) & (cfg_precision==2'b10);
  assign and_1202_rgt = (or_tmp_151 | or_90_cse) & or_309_cse;
  assign and_1207_rgt = and_dcpl_645 & IsNaN_8U_23U_land_5_lpi_1_dfm_9 & (cfg_precision==2'b10);
  assign and_1210_rgt = and_dcpl_645 & (~ IsNaN_8U_23U_land_5_lpi_1_dfm_9) & (cfg_precision==2'b10);
  assign and_1211_rgt = (or_tmp_147 | or_90_cse) & or_309_cse;
  assign and_1216_rgt = and_dcpl_654 & IsNaN_8U_23U_land_4_lpi_1_dfm_9 & (cfg_precision==2'b10);
  assign and_1219_rgt = and_dcpl_654 & (~ IsNaN_8U_23U_land_4_lpi_1_dfm_9) & (cfg_precision==2'b10);
  assign and_1220_rgt = (or_tmp_141 | or_90_cse) & or_309_cse;
  assign and_1225_rgt = and_dcpl_663 & IsNaN_8U_23U_land_3_lpi_1_dfm_9 & (cfg_precision==2'b10);
  assign and_1228_rgt = and_dcpl_663 & (~ IsNaN_8U_23U_land_3_lpi_1_dfm_9) & (cfg_precision==2'b10);
  assign and_1229_rgt = (or_tmp_134 | or_90_cse) & or_309_cse;
  assign and_1234_rgt = and_dcpl_672 & IsNaN_8U_23U_land_2_lpi_1_dfm_9 & (cfg_precision==2'b10);
  assign and_1237_rgt = and_dcpl_672 & (~ IsNaN_8U_23U_land_2_lpi_1_dfm_9) & (cfg_precision==2'b10);
  assign and_1238_rgt = (or_tmp_128 | or_90_cse) & or_309_cse;
  assign and_1243_rgt = and_dcpl_681 & IsNaN_8U_23U_land_1_lpi_1_dfm_9 & (cfg_precision==2'b10);
  assign and_1246_rgt = and_dcpl_681 & (~ IsNaN_8U_23U_land_1_lpi_1_dfm_9) & (cfg_precision==2'b10);
  assign and_1247_rgt = (or_tmp_122 | or_90_cse) & or_309_cse;
  assign and_1252_rgt = (mul_loop_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_3_lpi_1_dfm_4_cse
      | (cfg_precision!=2'b10)) & or_309_cse;
  assign and_1257_rgt = (mul_loop_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_4_lpi_1_dfm_4_cse
      | (cfg_precision!=2'b10)) & or_309_cse;
  assign and_1262_rgt = (mul_loop_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_5_lpi_1_dfm_4_cse
      | (cfg_precision!=2'b10)) & or_309_cse;
  assign and_1267_rgt = (mul_loop_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_6_lpi_1_dfm_4_cse
      | (cfg_precision!=2'b10)) & or_309_cse;
  assign and_1272_rgt = (mul_loop_mul_5_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_7_lpi_1_dfm_4_cse
      | (cfg_precision!=2'b10)) & or_309_cse;
  assign and_1277_rgt = (mul_loop_mul_6_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_8_lpi_1_dfm_4_cse
      | (cfg_precision!=2'b10)) & or_309_cse;
  assign and_1282_rgt = (mul_loop_mul_7_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_9_lpi_1_dfm_4_cse
      | (cfg_precision!=2'b10)) & or_309_cse;
  assign and_1287_rgt = (mul_loop_mul_8_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_10_lpi_1_dfm_4_cse
      | (cfg_precision!=2'b10)) & or_309_cse;
  assign and_1292_rgt = (mul_loop_mul_9_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_11_lpi_1_dfm_4_cse
      | (cfg_precision!=2'b10)) & or_309_cse;
  assign and_1297_rgt = (mul_loop_mul_10_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_12_lpi_1_dfm_4_cse
      | (cfg_precision!=2'b10)) & or_309_cse;
  assign and_1302_rgt = (mul_loop_mul_11_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_13_lpi_1_dfm_4_cse
      | (cfg_precision!=2'b10)) & or_309_cse;
  assign and_1307_rgt = (mul_loop_mul_12_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_14_lpi_1_dfm_4_cse
      | (cfg_precision!=2'b10)) & or_309_cse;
  assign and_1312_rgt = (mul_loop_mul_13_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_15_lpi_1_dfm_4_cse
      | (cfg_precision!=2'b10)) & or_309_cse;
  assign and_1317_rgt = (mul_loop_mul_14_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_16_lpi_1_dfm_4_cse
      | (cfg_precision!=2'b10)) & or_309_cse;
  assign and_1322_rgt = (mul_loop_mul_15_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_17_lpi_1_dfm_4_cse
      | (cfg_precision!=2'b10)) & or_309_cse;
  assign and_1327_rgt = (mul_loop_mul_16_FpMul_8U_23U_oelse_1_acc_itm_9_1 | reg_FpMul_8U_23U_lor_lpi_1_dfm_4_cse
      | (cfg_precision!=2'b10)) & or_309_cse;
  assign and_384_cse = FpMul_8U_23U_lor_3_lpi_1_dfm_st & or_2577_cse;
  assign nor_749_cse = ~((~ cfg_mul_src_1_sva_st_1) | chn_mul_op_rsci_bawt);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_cse = core_wen & ((and_dcpl_873
      & and_dcpl_72 & or_dcpl_206 & and_dcpl_259 & and_dcpl_255 & and_dcpl_254 &
      (else_mux_2_tmp[1:0]==2'b11) & (~ IsNaN_5U_23U_nor_tmp)) | and_dcpl_879);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_3_cse = core_wen & ((and_dcpl_873
      & and_dcpl_72 & or_dcpl_218 & and_dcpl_274 & and_dcpl_270 & and_dcpl_269 &
      (else_mux_5_tmp[1:0]==2'b11) & (~ IsNaN_5U_23U_nor_1_tmp)) | and_dcpl_891);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_6_cse = core_wen & ((and_dcpl_873
      & and_dcpl_72 & or_dcpl_228 & and_dcpl_289 & and_dcpl_285 & and_dcpl_284 &
      (else_mux_8_tmp[1:0]==2'b11) & (~ IsNaN_5U_23U_nor_2_tmp)) | and_dcpl_903);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_9_cse = core_wen & ((and_dcpl_873
      & and_dcpl_72 & or_dcpl_238 & and_dcpl_304 & and_dcpl_300 & and_dcpl_299 &
      (else_mux_11_tmp[1:0]==2'b11) & (~ IsNaN_5U_23U_nor_3_tmp)) | and_dcpl_915);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_12_cse = core_wen & ((and_dcpl_873
      & and_dcpl_72 & or_dcpl_248 & and_dcpl_319 & and_dcpl_315 & and_dcpl_314 &
      (else_mux_14_tmp[1:0]==2'b11) & (~ IsNaN_5U_23U_nor_4_tmp)) | and_dcpl_927);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_15_cse = core_wen & ((and_dcpl_873
      & and_dcpl_72 & or_dcpl_258 & and_dcpl_334 & and_dcpl_330 & and_dcpl_329 &
      (else_mux_17_tmp[1:0]==2'b11) & (~ IsNaN_5U_23U_nor_5_tmp)) | and_dcpl_939);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_18_cse = core_wen & ((and_dcpl_873
      & and_dcpl_72 & or_dcpl_268 & and_dcpl_349 & (else_mux_20_tmp[2]) & and_dcpl_345
      & and_dcpl_344 & (~ IsNaN_5U_23U_nor_6_tmp) & and_dcpl_85) | and_dcpl_951);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_21_cse = core_wen & ((and_dcpl_873
      & and_dcpl_72 & or_dcpl_278 & and_dcpl_364 & (else_mux_23_tmp[4]) & and_dcpl_360
      & and_dcpl_359 & (~ IsNaN_5U_23U_nor_7_tmp) & and_dcpl_85) | and_dcpl_963);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_24_cse = core_wen & ((and_dcpl_873
      & and_dcpl_72 & or_dcpl_288 & and_dcpl_379 & (else_mux_26_tmp[4]) & and_dcpl_375
      & and_dcpl_374 & (~ IsNaN_5U_23U_nor_8_tmp) & and_dcpl_85) | and_dcpl_975);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_27_cse = core_wen & ((and_dcpl_873
      & and_dcpl_72 & or_dcpl_298 & and_dcpl_394 & and_dcpl_390 & and_dcpl_389 &
      (else_mux_29_tmp[3]) & (else_mux_29_tmp[2]) & (else_mux_29_tmp[0])) | and_dcpl_987);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_30_cse = core_wen & ((and_dcpl_873
      & and_dcpl_72 & or_dcpl_308 & and_dcpl_409 & and_dcpl_405 & and_dcpl_404 &
      (else_mux_32_tmp[1]) & (else_mux_32_tmp[0]) & (else_mux_32_tmp[4])) | and_dcpl_999);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_33_cse = core_wen & ((and_dcpl_873
      & and_dcpl_72 & or_dcpl_318 & and_dcpl_424 & and_dcpl_420 & and_dcpl_419 &
      (else_mux_35_tmp[3]) & (else_mux_35_tmp[1]) & (else_mux_35_tmp[0])) | and_dcpl_1011);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_36_cse = core_wen & ((and_dcpl_873
      & and_dcpl_72 & or_dcpl_328 & and_dcpl_439 & and_dcpl_435 & and_dcpl_434 &
      (else_mux_38_tmp[2:0]==3'b111)) | and_dcpl_1023);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_39_cse = core_wen & ((and_dcpl_873
      & and_dcpl_72 & or_dcpl_338 & and_dcpl_454 & and_dcpl_450 & and_dcpl_449 &
      (else_mux_41_tmp[3]) & (else_mux_41_tmp[2]) & (else_mux_41_tmp[0])) | and_dcpl_1035);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_42_cse = core_wen & ((and_dcpl_873
      & and_dcpl_72 & or_dcpl_348 & and_dcpl_469 & and_dcpl_465 & and_dcpl_464 &
      (else_mux_44_tmp[1]) & (else_mux_44_tmp[0]) & (else_mux_44_tmp[4])) | and_dcpl_1047);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_45_cse = core_wen & ((and_dcpl_873
      & and_dcpl_72 & or_dcpl_358 & and_dcpl_484 & and_dcpl_480 & and_dcpl_479 &
      (else_mux_47_tmp[3]) & (else_mux_47_tmp[1]) & (else_mux_47_tmp[0])) | and_dcpl_1059);
  assign IsZero_8U_23U_aelse_and_16_cse = core_wen & (~(and_dcpl_53 | and_dcpl_50
      | (cfg_mul_prelu_rsci_d & (~ (chn_mul_in_rsci_d_mxwt[31]))) | or_dcpl_665 |
      (fsm_output[0])));
  assign IsZero_8U_23U_aelse_and_17_cse = core_wen & (~(and_dcpl_53 | and_dcpl_50
      | (cfg_mul_prelu_rsci_d & (~ (chn_mul_in_rsci_d_mxwt[64]))) | or_dcpl_665 |
      (fsm_output[0])));
  assign IsZero_8U_23U_aelse_and_18_cse = core_wen & (~(and_dcpl_53 | and_dcpl_50
      | (cfg_mul_prelu_rsci_d & (~ (chn_mul_in_rsci_d_mxwt[97]))) | or_dcpl_665 |
      (fsm_output[0])));
  assign IsZero_8U_23U_aelse_and_19_cse = core_wen & (~(and_dcpl_53 | and_dcpl_50
      | (cfg_mul_prelu_rsci_d & (~ (chn_mul_in_rsci_d_mxwt[130]))) | or_dcpl_665
      | (fsm_output[0])));
  assign IsZero_8U_23U_aelse_and_20_cse = core_wen & (~(and_dcpl_53 | and_dcpl_50
      | (cfg_mul_prelu_rsci_d & (~ (chn_mul_in_rsci_d_mxwt[163]))) | or_dcpl_665
      | (fsm_output[0])));
  assign IsZero_8U_23U_aelse_and_21_cse = core_wen & (~(and_dcpl_53 | and_dcpl_50
      | (cfg_mul_prelu_rsci_d & (~ (chn_mul_in_rsci_d_mxwt[196]))) | or_dcpl_665
      | (fsm_output[0])));
  assign IsZero_8U_23U_aelse_and_22_cse = core_wen & (~(and_dcpl_53 | and_dcpl_50
      | (cfg_mul_prelu_rsci_d & (~ (chn_mul_in_rsci_d_mxwt[229]))) | or_dcpl_665
      | (fsm_output[0])));
  assign IsZero_8U_23U_aelse_and_23_cse = core_wen & (~(and_dcpl_53 | and_dcpl_50
      | (cfg_mul_prelu_rsci_d & (~ (chn_mul_in_rsci_d_mxwt[262]))) | or_dcpl_665
      | (fsm_output[0])));
  assign IsZero_8U_23U_aelse_and_24_cse = core_wen & (~(and_dcpl_53 | and_dcpl_50
      | (cfg_mul_prelu_rsci_d & (~ (chn_mul_in_rsci_d_mxwt[295]))) | or_dcpl_665
      | (fsm_output[0])));
  assign IsZero_8U_23U_aelse_and_25_cse = core_wen & (~(and_dcpl_53 | and_dcpl_50
      | (cfg_mul_prelu_rsci_d & (~ (chn_mul_in_rsci_d_mxwt[328]))) | or_dcpl_665
      | (fsm_output[0])));
  assign IsZero_8U_23U_aelse_and_26_cse = core_wen & (~(and_dcpl_53 | and_dcpl_50
      | (cfg_mul_prelu_rsci_d & (~ (chn_mul_in_rsci_d_mxwt[361]))) | or_dcpl_665
      | (fsm_output[0])));
  assign IsZero_8U_23U_aelse_and_27_cse = core_wen & (~(and_dcpl_53 | and_dcpl_50
      | (cfg_mul_prelu_rsci_d & (~ (chn_mul_in_rsci_d_mxwt[394]))) | or_dcpl_665
      | (fsm_output[0])));
  assign IsZero_8U_23U_aelse_and_28_cse = core_wen & (~(and_dcpl_53 | and_dcpl_50
      | (cfg_mul_prelu_rsci_d & (~ (chn_mul_in_rsci_d_mxwt[427]))) | or_dcpl_665
      | (fsm_output[0])));
  assign IsZero_8U_23U_aelse_and_29_cse = core_wen & (~(and_dcpl_53 | and_dcpl_50
      | (cfg_mul_prelu_rsci_d & (~ (chn_mul_in_rsci_d_mxwt[460]))) | or_dcpl_665
      | (fsm_output[0])));
  assign IsZero_8U_23U_aelse_and_30_cse = core_wen & (~(and_dcpl_53 | and_dcpl_50
      | (cfg_mul_prelu_rsci_d & (~ (chn_mul_in_rsci_d_mxwt[493]))) | or_dcpl_665
      | (fsm_output[0])));
  assign IsZero_8U_23U_aelse_and_31_cse = core_wen & (~(and_dcpl_53 | and_dcpl_50
      | (cfg_mul_prelu_rsci_d & (~ (chn_mul_in_rsci_d_mxwt[526]))) | or_dcpl_665
      | (fsm_output[0])));
  assign or_70_cse = (~ cfg_mul_prelu_rsci_d) | (chn_mul_in_rsci_d_mxwt[31]);
  assign and_552_nl = and_dcpl_7 & or_70_cse & and_dcpl_2 & (fsm_output[1]);
  assign mul_loop_mul_1_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_552_nl);
  assign or_75_cse = (~ cfg_mul_prelu_rsci_d) | (chn_mul_in_rsci_d_mxwt[64]);
  assign and_554_nl = and_dcpl_7 & or_75_cse & and_dcpl_2 & (fsm_output[1]);
  assign mul_loop_mul_2_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_554_nl);
  assign or_76_cse = (~ cfg_mul_prelu_rsci_d) | (chn_mul_in_rsci_d_mxwt[97]);
  assign and_556_nl = and_dcpl_7 & or_76_cse & and_dcpl_2 & (fsm_output[1]);
  assign mul_loop_mul_3_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_556_nl);
  assign or_77_cse = (~ cfg_mul_prelu_rsci_d) | (chn_mul_in_rsci_d_mxwt[130]);
  assign and_558_nl = and_dcpl_7 & or_77_cse & and_dcpl_2 & (fsm_output[1]);
  assign mul_loop_mul_4_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_558_nl);
  assign or_78_cse = (~ cfg_mul_prelu_rsci_d) | (chn_mul_in_rsci_d_mxwt[163]);
  assign and_560_nl = and_dcpl_7 & or_78_cse & and_dcpl_2 & (fsm_output[1]);
  assign mul_loop_mul_5_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_560_nl);
  assign or_79_cse = (~ cfg_mul_prelu_rsci_d) | (chn_mul_in_rsci_d_mxwt[196]);
  assign and_562_nl = and_dcpl_7 & or_79_cse & and_dcpl_2 & (fsm_output[1]);
  assign mul_loop_mul_6_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_562_nl);
  assign or_80_cse = (~ cfg_mul_prelu_rsci_d) | (chn_mul_in_rsci_d_mxwt[229]);
  assign and_564_nl = and_dcpl_7 & or_80_cse & and_dcpl_2 & (fsm_output[1]);
  assign mul_loop_mul_7_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_564_nl);
  assign or_81_cse = (~ cfg_mul_prelu_rsci_d) | (chn_mul_in_rsci_d_mxwt[262]);
  assign and_566_nl = and_dcpl_7 & or_81_cse & and_dcpl_2 & (fsm_output[1]);
  assign mul_loop_mul_8_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_566_nl);
  assign or_82_cse = (~ cfg_mul_prelu_rsci_d) | (chn_mul_in_rsci_d_mxwt[295]);
  assign and_568_nl = and_dcpl_7 & or_82_cse & and_dcpl_2 & (fsm_output[1]);
  assign mul_loop_mul_9_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_568_nl);
  assign or_83_cse = (~ cfg_mul_prelu_rsci_d) | (chn_mul_in_rsci_d_mxwt[328]);
  assign and_570_nl = and_dcpl_7 & or_83_cse & and_dcpl_2 & (fsm_output[1]);
  assign mul_loop_mul_10_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_570_nl);
  assign or_84_cse = (~ cfg_mul_prelu_rsci_d) | (chn_mul_in_rsci_d_mxwt[361]);
  assign and_572_nl = and_dcpl_7 & or_84_cse & and_dcpl_2 & (fsm_output[1]);
  assign mul_loop_mul_11_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_572_nl);
  assign or_85_cse = (~ cfg_mul_prelu_rsci_d) | (chn_mul_in_rsci_d_mxwt[394]);
  assign and_574_nl = and_dcpl_7 & or_85_cse & and_dcpl_2 & (fsm_output[1]);
  assign mul_loop_mul_12_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_574_nl);
  assign or_86_cse = (~ cfg_mul_prelu_rsci_d) | (chn_mul_in_rsci_d_mxwt[427]);
  assign and_576_nl = and_dcpl_7 & or_86_cse & and_dcpl_2 & (fsm_output[1]);
  assign mul_loop_mul_13_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_576_nl);
  assign or_87_cse = (~ cfg_mul_prelu_rsci_d) | (chn_mul_in_rsci_d_mxwt[460]);
  assign and_578_nl = and_dcpl_7 & or_87_cse & and_dcpl_2 & (fsm_output[1]);
  assign mul_loop_mul_14_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_578_nl);
  assign or_88_cse = (~ cfg_mul_prelu_rsci_d) | (chn_mul_in_rsci_d_mxwt[493]);
  assign and_580_nl = and_dcpl_7 & or_88_cse & and_dcpl_2 & (fsm_output[1]);
  assign mul_loop_mul_15_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_580_nl);
  assign or_89_cse = (~ cfg_mul_prelu_rsci_d) | (chn_mul_in_rsci_d_mxwt[526]);
  assign and_582_nl = and_dcpl_7 & or_89_cse & and_dcpl_2 & (fsm_output[1]);
  assign mul_loop_mul_16_X_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_582_nl);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_65_nl
      = MUX_v_2_2_2(2'b00, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_sva_1[3:2]),
      FpExpoWidthInc_5U_8U_23U_1U_1U_exs_261_0);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_178_nl = MUX_v_2_2_2(2'b1, (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_65_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_3_2_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_178_nl)
      | ({{1{IsInf_5U_23U_land_1_lpi_1_dfm}}, IsInf_5U_23U_land_1_lpi_1_dfm}) | ({{1{IsNaN_5U_23U_land_1_lpi_1_dfm}},
      IsNaN_5U_23U_land_1_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_2_nl =
      MUX_v_2_2_2(2'b00, ({{1{FpExpoWidthInc_5U_8U_23U_1U_1U_exs_261_0}}, FpExpoWidthInc_5U_8U_23U_1U_1U_exs_261_0}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_sva_1[0]));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_144_nl = MUX_v_2_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_1_sva[5:4]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_2_nl), FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_1_0_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_144_nl)
      | ({{1{IsInf_5U_23U_land_1_lpi_1_dfm}}, IsInf_5U_23U_land_1_lpi_1_dfm}) | ({{1{IsNaN_5U_23U_land_1_lpi_1_dfm}},
      IsNaN_5U_23U_land_1_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_nl =
      MUX1HOT_v_4_3_2((mul_nan_to_zero_op_expo_1_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_1_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_ssc
      , IsDenorm_5U_23U_land_1_lpi_1_dfm , IsInf_5U_23U_land_1_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_nl),
      4'b1111, IsNaN_5U_23U_land_1_lpi_1_dfm);
  assign FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_tmp = IsZero_8U_23U_1_land_1_lpi_1_dfm_mx0w0
      | IsZero_8U_23U_land_1_lpi_1_dfm_7;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_67_nl
      = MUX_v_2_2_2(2'b00, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_sva_1[3:2]),
      FpExpoWidthInc_5U_8U_23U_1U_1U_exs_267_0);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_182_nl = MUX_v_2_2_2(2'b1, (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_67_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_3_2_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_182_nl)
      | ({{1{IsInf_5U_23U_land_2_lpi_1_dfm}}, IsInf_5U_23U_land_2_lpi_1_dfm}) | ({{1{IsNaN_5U_23U_land_2_lpi_1_dfm}},
      IsNaN_5U_23U_land_2_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_6_nl =
      MUX_v_2_2_2(2'b00, ({{1{FpExpoWidthInc_5U_8U_23U_1U_1U_exs_267_0}}, FpExpoWidthInc_5U_8U_23U_1U_1U_exs_267_0}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_sva_1[0]));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_146_nl = MUX_v_2_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_2_sva[5:4]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_6_nl), FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_1_0_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_146_nl)
      | ({{1{IsInf_5U_23U_land_2_lpi_1_dfm}}, IsInf_5U_23U_land_2_lpi_1_dfm}) | ({{1{IsNaN_5U_23U_land_2_lpi_1_dfm}},
      IsNaN_5U_23U_land_2_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_1_nl
      = MUX1HOT_v_4_3_2((mul_nan_to_zero_op_expo_2_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_2_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_ssc
      , IsDenorm_5U_23U_land_2_lpi_1_dfm , IsInf_5U_23U_land_2_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_1_nl),
      4'b1111, IsNaN_5U_23U_land_2_lpi_1_dfm);
  assign FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_2_tmp = IsZero_8U_23U_1_land_2_lpi_1_dfm_mx0w0
      | IsZero_8U_23U_land_2_lpi_1_dfm_7;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_69_nl
      = MUX_v_2_2_2(2'b00, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_sva_1[3:2]),
      FpExpoWidthInc_5U_8U_23U_1U_1U_exs_273_0);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_186_nl = MUX_v_2_2_2(2'b1, (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_69_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_3_2_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_186_nl)
      | ({{1{IsInf_5U_23U_land_3_lpi_1_dfm}}, IsInf_5U_23U_land_3_lpi_1_dfm}) | ({{1{IsNaN_5U_23U_land_3_lpi_1_dfm}},
      IsNaN_5U_23U_land_3_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_10_nl
      = MUX_v_2_2_2(2'b00, ({{1{FpExpoWidthInc_5U_8U_23U_1U_1U_exs_273_0}}, FpExpoWidthInc_5U_8U_23U_1U_1U_exs_273_0}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_sva_1[0]));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_148_nl = MUX_v_2_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_3_sva[5:4]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_10_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_1_0_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_148_nl)
      | ({{1{IsInf_5U_23U_land_3_lpi_1_dfm}}, IsInf_5U_23U_land_3_lpi_1_dfm}) | ({{1{IsNaN_5U_23U_land_3_lpi_1_dfm}},
      IsNaN_5U_23U_land_3_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_2_nl
      = MUX1HOT_v_4_3_2((mul_nan_to_zero_op_expo_3_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_3_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_ssc
      , IsDenorm_5U_23U_land_3_lpi_1_dfm , IsInf_5U_23U_land_3_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_2_nl),
      4'b1111, IsNaN_5U_23U_land_3_lpi_1_dfm);
  assign FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_4_tmp = IsZero_8U_23U_1_land_3_lpi_1_dfm_mx0w0
      | IsZero_8U_23U_land_3_lpi_1_dfm_7;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_71_nl
      = MUX_v_2_2_2(2'b00, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_sva_1[3:2]),
      FpExpoWidthInc_5U_8U_23U_1U_1U_exs_279_0);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_190_nl = MUX_v_2_2_2(2'b1, (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_71_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_3_2_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_190_nl)
      | ({{1{IsInf_5U_23U_land_4_lpi_1_dfm}}, IsInf_5U_23U_land_4_lpi_1_dfm}) | ({{1{IsNaN_5U_23U_land_4_lpi_1_dfm}},
      IsNaN_5U_23U_land_4_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_14_nl
      = MUX_v_2_2_2(2'b00, ({{1{FpExpoWidthInc_5U_8U_23U_1U_1U_exs_279_0}}, FpExpoWidthInc_5U_8U_23U_1U_1U_exs_279_0}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_sva_1[0]));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_150_nl = MUX_v_2_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_4_sva[5:4]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_14_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_1_0_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_150_nl)
      | ({{1{IsInf_5U_23U_land_4_lpi_1_dfm}}, IsInf_5U_23U_land_4_lpi_1_dfm}) | ({{1{IsNaN_5U_23U_land_4_lpi_1_dfm}},
      IsNaN_5U_23U_land_4_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_3_nl
      = MUX1HOT_v_4_3_2((mul_nan_to_zero_op_expo_4_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_4_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_ssc
      , IsDenorm_5U_23U_land_4_lpi_1_dfm , IsInf_5U_23U_land_4_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_3_nl),
      4'b1111, IsNaN_5U_23U_land_4_lpi_1_dfm);
  assign FpMul_8U_23U_lor_6_lpi_1_dfm_mx0w0 = IsZero_8U_23U_1_land_4_lpi_1_dfm_mx0w0
      | IsZero_8U_23U_land_4_lpi_1_dfm_7;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_73_nl
      = MUX_v_2_2_2(2'b00, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_sva_1[3:2]),
      FpExpoWidthInc_5U_8U_23U_1U_1U_exs_285_0);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_194_nl = MUX_v_2_2_2(2'b1, (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_73_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_3_2_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_194_nl)
      | ({{1{IsInf_5U_23U_land_5_lpi_1_dfm}}, IsInf_5U_23U_land_5_lpi_1_dfm}) | ({{1{IsNaN_5U_23U_land_5_lpi_1_dfm}},
      IsNaN_5U_23U_land_5_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_18_nl
      = MUX_v_2_2_2(2'b00, ({{1{FpExpoWidthInc_5U_8U_23U_1U_1U_exs_285_0}}, FpExpoWidthInc_5U_8U_23U_1U_1U_exs_285_0}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_sva_1[0]));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_152_nl = MUX_v_2_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_5_sva[5:4]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_18_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_1_0_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_152_nl)
      | ({{1{IsInf_5U_23U_land_5_lpi_1_dfm}}, IsInf_5U_23U_land_5_lpi_1_dfm}) | ({{1{IsNaN_5U_23U_land_5_lpi_1_dfm}},
      IsNaN_5U_23U_land_5_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_4_nl
      = MUX1HOT_v_4_3_2((mul_nan_to_zero_op_expo_5_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_5_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_ssc
      , IsDenorm_5U_23U_land_5_lpi_1_dfm , IsInf_5U_23U_land_5_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_4_nl),
      4'b1111, IsNaN_5U_23U_land_5_lpi_1_dfm);
  assign FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_8_tmp = IsZero_8U_23U_1_land_5_lpi_1_dfm_mx0w0
      | IsZero_8U_23U_land_5_lpi_1_dfm_7;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_75_nl
      = MUX_v_2_2_2(2'b00, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_sva_1[3:2]),
      FpExpoWidthInc_5U_8U_23U_1U_1U_exs_291_0);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_198_nl = MUX_v_2_2_2(2'b1, (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_75_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_3_2_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_198_nl)
      | ({{1{IsInf_5U_23U_land_6_lpi_1_dfm}}, IsInf_5U_23U_land_6_lpi_1_dfm}) | ({{1{IsNaN_5U_23U_land_6_lpi_1_dfm}},
      IsNaN_5U_23U_land_6_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_22_nl
      = MUX_v_2_2_2(2'b00, ({{1{FpExpoWidthInc_5U_8U_23U_1U_1U_exs_291_0}}, FpExpoWidthInc_5U_8U_23U_1U_1U_exs_291_0}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_sva_1[0]));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_154_nl = MUX_v_2_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_6_sva[5:4]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_22_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_1_0_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_154_nl)
      | ({{1{IsInf_5U_23U_land_6_lpi_1_dfm}}, IsInf_5U_23U_land_6_lpi_1_dfm}) | ({{1{IsNaN_5U_23U_land_6_lpi_1_dfm}},
      IsNaN_5U_23U_land_6_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_5_nl
      = MUX1HOT_v_4_3_2((mul_nan_to_zero_op_expo_6_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_6_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_ssc
      , IsDenorm_5U_23U_land_6_lpi_1_dfm , IsInf_5U_23U_land_6_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_5_nl),
      4'b1111, IsNaN_5U_23U_land_6_lpi_1_dfm);
  assign FpMul_8U_23U_lor_8_lpi_1_dfm_mx0w0 = IsZero_8U_23U_1_land_6_lpi_1_dfm_mx0w0
      | IsZero_8U_23U_land_6_lpi_1_dfm_7;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_77_nl
      = MUX_v_2_2_2(2'b00, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_sva_1[3:2]),
      FpExpoWidthInc_5U_8U_23U_1U_1U_exs_297_0);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_202_nl = MUX_v_2_2_2(2'b1, (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_77_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_3_2_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_202_nl)
      | ({{1{IsInf_5U_23U_land_7_lpi_1_dfm}}, IsInf_5U_23U_land_7_lpi_1_dfm}) | ({{1{IsNaN_5U_23U_land_7_lpi_1_dfm}},
      IsNaN_5U_23U_land_7_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_26_nl
      = MUX_v_2_2_2(2'b00, ({{1{FpExpoWidthInc_5U_8U_23U_1U_1U_exs_297_0}}, FpExpoWidthInc_5U_8U_23U_1U_1U_exs_297_0}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_sva_1[0]));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_156_nl = MUX_v_2_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_7_sva[5:4]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_26_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_1_0_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_156_nl)
      | ({{1{IsInf_5U_23U_land_7_lpi_1_dfm}}, IsInf_5U_23U_land_7_lpi_1_dfm}) | ({{1{IsNaN_5U_23U_land_7_lpi_1_dfm}},
      IsNaN_5U_23U_land_7_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_6_nl
      = MUX1HOT_v_4_3_2((mul_nan_to_zero_op_expo_7_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_7_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_ssc
      , IsDenorm_5U_23U_land_7_lpi_1_dfm , IsInf_5U_23U_land_7_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_6_nl),
      4'b1111, IsNaN_5U_23U_land_7_lpi_1_dfm);
  assign FpMul_8U_23U_lor_9_lpi_1_dfm_mx0w0 = IsZero_8U_23U_1_land_7_lpi_1_dfm_mx0w0
      | IsZero_8U_23U_land_7_lpi_1_dfm_7;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_79_nl
      = MUX_v_2_2_2(2'b00, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_sva_1[3:2]),
      FpExpoWidthInc_5U_8U_23U_1U_1U_exs_303_0);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_206_nl = MUX_v_2_2_2(2'b1, (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_79_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_3_2_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_206_nl)
      | ({{1{IsInf_5U_23U_land_8_lpi_1_dfm}}, IsInf_5U_23U_land_8_lpi_1_dfm}) | ({{1{IsNaN_5U_23U_land_8_lpi_1_dfm}},
      IsNaN_5U_23U_land_8_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_30_nl
      = MUX_v_2_2_2(2'b00, ({{1{FpExpoWidthInc_5U_8U_23U_1U_1U_exs_303_0}}, FpExpoWidthInc_5U_8U_23U_1U_1U_exs_303_0}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_sva_1[0]));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_158_nl = MUX_v_2_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_8_sva[5:4]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_30_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_1_0_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_158_nl)
      | ({{1{IsInf_5U_23U_land_8_lpi_1_dfm}}, IsInf_5U_23U_land_8_lpi_1_dfm}) | ({{1{IsNaN_5U_23U_land_8_lpi_1_dfm}},
      IsNaN_5U_23U_land_8_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_7_nl
      = MUX1HOT_v_4_3_2((mul_nan_to_zero_op_expo_8_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_8_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_ssc
      , IsDenorm_5U_23U_land_8_lpi_1_dfm , IsInf_5U_23U_land_8_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_7_nl),
      4'b1111, IsNaN_5U_23U_land_8_lpi_1_dfm);
  assign FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_14_tmp = IsZero_8U_23U_1_land_8_lpi_1_dfm_mx0w0
      | IsZero_8U_23U_land_8_lpi_1_dfm_7;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_81_nl
      = MUX_v_2_2_2(2'b00, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_sva_1[3:2]),
      FpExpoWidthInc_5U_8U_23U_1U_1U_exs_309_0);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_210_nl = MUX_v_2_2_2(2'b1, (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_81_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_16_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_3_2_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_210_nl)
      | ({{1{IsInf_5U_23U_land_9_lpi_1_dfm}}, IsInf_5U_23U_land_9_lpi_1_dfm}) | ({{1{IsNaN_5U_23U_land_9_lpi_1_dfm}},
      IsNaN_5U_23U_land_9_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_34_nl
      = MUX_v_2_2_2(2'b00, ({{1{FpExpoWidthInc_5U_8U_23U_1U_1U_exs_309_0}}, FpExpoWidthInc_5U_8U_23U_1U_1U_exs_309_0}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_sva_1[0]));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_160_nl = MUX_v_2_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_9_sva[5:4]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_34_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_16_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_1_0_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_160_nl)
      | ({{1{IsInf_5U_23U_land_9_lpi_1_dfm}}, IsInf_5U_23U_land_9_lpi_1_dfm}) | ({{1{IsNaN_5U_23U_land_9_lpi_1_dfm}},
      IsNaN_5U_23U_land_9_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_8_nl
      = MUX1HOT_v_4_3_2((mul_nan_to_zero_op_expo_9_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_9_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_16_ssc
      , IsDenorm_5U_23U_land_9_lpi_1_dfm , IsInf_5U_23U_land_9_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_8_nl),
      4'b1111, IsNaN_5U_23U_land_9_lpi_1_dfm);
  assign FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_16_tmp = IsZero_8U_23U_1_land_9_lpi_1_dfm_mx0w0
      | IsZero_8U_23U_land_9_lpi_1_dfm_7;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_83_nl
      = MUX_v_2_2_2(2'b00, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_sva_1[3:2]),
      FpExpoWidthInc_5U_8U_23U_1U_1U_exs_315_0);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_214_nl = MUX_v_2_2_2(2'b1, (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_83_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_18_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_3_2_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_214_nl)
      | ({{1{IsInf_5U_23U_land_10_lpi_1_dfm}}, IsInf_5U_23U_land_10_lpi_1_dfm}) |
      ({{1{IsNaN_5U_23U_land_10_lpi_1_dfm}}, IsNaN_5U_23U_land_10_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_38_nl
      = MUX_v_2_2_2(2'b00, ({{1{FpExpoWidthInc_5U_8U_23U_1U_1U_exs_315_0}}, FpExpoWidthInc_5U_8U_23U_1U_1U_exs_315_0}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_sva_1[0]));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_162_nl = MUX_v_2_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_10_sva[5:4]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_38_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_18_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_1_0_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_162_nl)
      | ({{1{IsInf_5U_23U_land_10_lpi_1_dfm}}, IsInf_5U_23U_land_10_lpi_1_dfm}) |
      ({{1{IsNaN_5U_23U_land_10_lpi_1_dfm}}, IsNaN_5U_23U_land_10_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_9_nl
      = MUX1HOT_v_4_3_2((mul_nan_to_zero_op_expo_10_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_10_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_18_ssc
      , IsDenorm_5U_23U_land_10_lpi_1_dfm , IsInf_5U_23U_land_10_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_9_nl),
      4'b1111, IsNaN_5U_23U_land_10_lpi_1_dfm);
  assign FpMul_8U_23U_lor_12_lpi_1_dfm_mx0w0 = IsZero_8U_23U_1_land_10_lpi_1_dfm_mx0w0
      | IsZero_8U_23U_land_10_lpi_1_dfm_7;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_85_nl
      = MUX_v_2_2_2(2'b00, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_sva_1[3:2]),
      FpExpoWidthInc_5U_8U_23U_1U_1U_exs_321_0);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_218_nl = MUX_v_2_2_2(2'b1, (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_85_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_20_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_3_2_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_218_nl)
      | ({{1{IsInf_5U_23U_land_11_lpi_1_dfm}}, IsInf_5U_23U_land_11_lpi_1_dfm}) |
      ({{1{IsNaN_5U_23U_land_11_lpi_1_dfm}}, IsNaN_5U_23U_land_11_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_42_nl
      = MUX_v_2_2_2(2'b00, ({{1{FpExpoWidthInc_5U_8U_23U_1U_1U_exs_321_0}}, FpExpoWidthInc_5U_8U_23U_1U_1U_exs_321_0}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_sva_1[0]));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_164_nl = MUX_v_2_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_11_sva[5:4]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_42_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_20_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_1_0_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_164_nl)
      | ({{1{IsInf_5U_23U_land_11_lpi_1_dfm}}, IsInf_5U_23U_land_11_lpi_1_dfm}) |
      ({{1{IsNaN_5U_23U_land_11_lpi_1_dfm}}, IsNaN_5U_23U_land_11_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_10_nl
      = MUX1HOT_v_4_3_2((mul_nan_to_zero_op_expo_11_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_11_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_20_ssc
      , IsDenorm_5U_23U_land_11_lpi_1_dfm , IsInf_5U_23U_land_11_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_10_nl),
      4'b1111, IsNaN_5U_23U_land_11_lpi_1_dfm);
  assign FpMul_8U_23U_lor_13_lpi_1_dfm_mx0w0 = IsZero_8U_23U_1_land_11_lpi_1_dfm_mx0w0
      | IsZero_8U_23U_land_11_lpi_1_dfm_7;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_87_nl
      = MUX_v_2_2_2(2'b00, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_sva_1[3:2]),
      FpExpoWidthInc_5U_8U_23U_1U_1U_exs_327_0);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_222_nl = MUX_v_2_2_2(2'b1, (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_87_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_22_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_3_2_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_222_nl)
      | ({{1{IsInf_5U_23U_land_12_lpi_1_dfm}}, IsInf_5U_23U_land_12_lpi_1_dfm}) |
      ({{1{IsNaN_5U_23U_land_12_lpi_1_dfm}}, IsNaN_5U_23U_land_12_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_46_nl
      = MUX_v_2_2_2(2'b00, ({{1{FpExpoWidthInc_5U_8U_23U_1U_1U_exs_327_0}}, FpExpoWidthInc_5U_8U_23U_1U_1U_exs_327_0}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_sva_1[0]));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_166_nl = MUX_v_2_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_12_sva[5:4]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_46_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_22_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_1_0_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_166_nl)
      | ({{1{IsInf_5U_23U_land_12_lpi_1_dfm}}, IsInf_5U_23U_land_12_lpi_1_dfm}) |
      ({{1{IsNaN_5U_23U_land_12_lpi_1_dfm}}, IsNaN_5U_23U_land_12_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_11_nl
      = MUX1HOT_v_4_3_2((mul_nan_to_zero_op_expo_12_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_12_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_22_ssc
      , IsDenorm_5U_23U_land_12_lpi_1_dfm , IsInf_5U_23U_land_12_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_11_nl),
      4'b1111, IsNaN_5U_23U_land_12_lpi_1_dfm);
  assign FpMul_8U_23U_lor_14_lpi_1_dfm_mx0w0 = IsZero_8U_23U_1_land_12_lpi_1_dfm_mx0w0
      | IsZero_8U_23U_land_12_lpi_1_dfm_7;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_89_nl
      = MUX_v_2_2_2(2'b00, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_sva_1[3:2]),
      FpExpoWidthInc_5U_8U_23U_1U_1U_exs_333_0);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_226_nl = MUX_v_2_2_2(2'b1, (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_89_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_24_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_3_2_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_226_nl)
      | ({{1{IsInf_5U_23U_land_13_lpi_1_dfm}}, IsInf_5U_23U_land_13_lpi_1_dfm}) |
      ({{1{IsNaN_5U_23U_land_13_lpi_1_dfm}}, IsNaN_5U_23U_land_13_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_50_nl
      = MUX_v_2_2_2(2'b00, ({{1{FpExpoWidthInc_5U_8U_23U_1U_1U_exs_333_0}}, FpExpoWidthInc_5U_8U_23U_1U_1U_exs_333_0}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_sva_1[0]));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_168_nl = MUX_v_2_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_13_sva[5:4]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_50_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_24_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_1_0_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_168_nl)
      | ({{1{IsInf_5U_23U_land_13_lpi_1_dfm}}, IsInf_5U_23U_land_13_lpi_1_dfm}) |
      ({{1{IsNaN_5U_23U_land_13_lpi_1_dfm}}, IsNaN_5U_23U_land_13_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_12_nl
      = MUX1HOT_v_4_3_2((mul_nan_to_zero_op_expo_13_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_13_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_24_ssc
      , IsDenorm_5U_23U_land_13_lpi_1_dfm , IsInf_5U_23U_land_13_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_12_nl),
      4'b1111, IsNaN_5U_23U_land_13_lpi_1_dfm);
  assign FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_24_tmp = IsZero_8U_23U_1_land_13_lpi_1_dfm_mx0w0
      | IsZero_8U_23U_land_13_lpi_1_dfm_7;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_91_nl
      = MUX_v_2_2_2(2'b00, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_sva_1[3:2]),
      FpExpoWidthInc_5U_8U_23U_1U_1U_exs_339_0);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_230_nl = MUX_v_2_2_2(2'b1, (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_91_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_26_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_3_2_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_230_nl)
      | ({{1{IsInf_5U_23U_land_14_lpi_1_dfm}}, IsInf_5U_23U_land_14_lpi_1_dfm}) |
      ({{1{IsNaN_5U_23U_land_14_lpi_1_dfm}}, IsNaN_5U_23U_land_14_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_54_nl
      = MUX_v_2_2_2(2'b00, ({{1{FpExpoWidthInc_5U_8U_23U_1U_1U_exs_339_0}}, FpExpoWidthInc_5U_8U_23U_1U_1U_exs_339_0}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_sva_1[0]));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_170_nl = MUX_v_2_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_14_sva[5:4]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_54_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_26_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_1_0_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_170_nl)
      | ({{1{IsInf_5U_23U_land_14_lpi_1_dfm}}, IsInf_5U_23U_land_14_lpi_1_dfm}) |
      ({{1{IsNaN_5U_23U_land_14_lpi_1_dfm}}, IsNaN_5U_23U_land_14_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_13_nl
      = MUX1HOT_v_4_3_2((mul_nan_to_zero_op_expo_14_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_14_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_26_ssc
      , IsDenorm_5U_23U_land_14_lpi_1_dfm , IsInf_5U_23U_land_14_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_13_nl),
      4'b1111, IsNaN_5U_23U_land_14_lpi_1_dfm);
  assign FpMul_8U_23U_lor_16_lpi_1_dfm_mx0w0 = IsZero_8U_23U_1_land_14_lpi_1_dfm_mx0w0
      | IsZero_8U_23U_land_14_lpi_1_dfm_7;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_93_nl
      = MUX_v_2_2_2(2'b00, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_sva_1[3:2]),
      FpExpoWidthInc_5U_8U_23U_1U_1U_exs_345_0);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_234_nl = MUX_v_2_2_2(2'b1, (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_93_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_28_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_3_2_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_234_nl)
      | ({{1{IsInf_5U_23U_land_15_lpi_1_dfm}}, IsInf_5U_23U_land_15_lpi_1_dfm}) |
      ({{1{IsNaN_5U_23U_land_15_lpi_1_dfm}}, IsNaN_5U_23U_land_15_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_58_nl
      = MUX_v_2_2_2(2'b00, ({{1{FpExpoWidthInc_5U_8U_23U_1U_1U_exs_345_0}}, FpExpoWidthInc_5U_8U_23U_1U_1U_exs_345_0}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_sva_1[0]));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_172_nl = MUX_v_2_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_15_sva[5:4]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_58_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_28_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_1_0_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_172_nl)
      | ({{1{IsInf_5U_23U_land_15_lpi_1_dfm}}, IsInf_5U_23U_land_15_lpi_1_dfm}) |
      ({{1{IsNaN_5U_23U_land_15_lpi_1_dfm}}, IsNaN_5U_23U_land_15_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_14_nl
      = MUX1HOT_v_4_3_2((mul_nan_to_zero_op_expo_15_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_15_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_28_ssc
      , IsDenorm_5U_23U_land_15_lpi_1_dfm , IsInf_5U_23U_land_15_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_14_nl),
      4'b1111, IsNaN_5U_23U_land_15_lpi_1_dfm);
  assign FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_28_tmp = IsZero_8U_23U_1_land_15_lpi_1_dfm_mx0w0
      | IsZero_8U_23U_land_15_lpi_1_dfm_7;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_95_nl
      = MUX_v_2_2_2(2'b00, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_sva_1[3:2]),
      FpExpoWidthInc_5U_8U_23U_1U_1U_exs_351_0);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_238_nl = MUX_v_2_2_2(2'b1, (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_95_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_30_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_3_2_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_238_nl)
      | ({{1{IsInf_5U_23U_land_lpi_1_dfm}}, IsInf_5U_23U_land_lpi_1_dfm}) | ({{1{IsNaN_5U_23U_land_lpi_1_dfm}},
      IsNaN_5U_23U_land_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_62_nl
      = MUX_v_2_2_2(2'b00, ({{1{FpExpoWidthInc_5U_8U_23U_1U_1U_exs_351_0}}, FpExpoWidthInc_5U_8U_23U_1U_1U_exs_351_0}),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_sva_1[0]));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_174_nl = MUX_v_2_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_sva[5:4]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_62_nl),
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_30_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_1_0_mx0w0 = (FpExpoWidthInc_5U_8U_23U_1U_1U_mux_174_nl)
      | ({{1{IsInf_5U_23U_land_lpi_1_dfm}}, IsInf_5U_23U_land_lpi_1_dfm}) | ({{1{IsNaN_5U_23U_land_lpi_1_dfm}},
      IsNaN_5U_23U_land_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_15_nl
      = MUX1HOT_v_4_3_2((mul_nan_to_zero_op_expo_lpi_1_dfm[3:0]), (FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_sva[3:0]),
      4'b1110, {FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_30_ssc
      , IsDenorm_5U_23U_land_lpi_1_dfm , IsInf_5U_23U_land_lpi_1_dfm});
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_mux1h_15_nl),
      4'b1111, IsNaN_5U_23U_land_lpi_1_dfm);
  assign FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_30_tmp = IsZero_8U_23U_1_land_lpi_1_dfm_mx0w0
      | IsZero_8U_23U_land_lpi_1_dfm_7;
  assign nl_FpMul_8U_23U_else_2_else_acc_nl = ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_8_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_8_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_10})
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_nl = nl_FpMul_8U_23U_else_2_else_acc_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_1_sva_1_mx0w0 = (FpMul_8U_23U_else_2_else_acc_nl)
      + (MulIn_data_sva_535[30:23]);
  assign FpMul_8U_23U_p_expo_1_sva_1_mx0w0 = nl_FpMul_8U_23U_p_expo_1_sva_1_mx0w0[7:0];
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_mx0w0 = ~(mul_loop_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      & (mul_loop_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47]));
  assign mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs_mx0w0 = FpMantRNE_48U_24U_else_carry_1_sva_mx0w0
      & (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_1_sva_mx0w0 = (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_1_sva_mx1[0]) & (FpMul_8U_23U_p_mant_p1_1_sva_mx1[47]))
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_FpMul_8U_23U_and_itm_mx0w0 = (mul_loop_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      | (~ (FpMul_8U_23U_p_mant_p1_1_sva_mx1[47]))) & mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign nl_FpMul_8U_23U_else_2_else_acc_2_nl = ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_8_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_8_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_10})
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_2_nl = nl_FpMul_8U_23U_else_2_else_acc_2_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_2_sva_1_mx0w0 = (FpMul_8U_23U_else_2_else_acc_2_nl)
      + (MulIn_data_sva_535[63:56]);
  assign FpMul_8U_23U_p_expo_2_sva_1_mx0w0 = nl_FpMul_8U_23U_p_expo_2_sva_1_mx0w0[7:0];
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_mx0w0 = ~(mul_loop_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      & (mul_loop_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47]));
  assign mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs_mx0w0 = FpMantRNE_48U_24U_else_carry_2_sva_mx0w0
      & (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_2_sva_mx0w0 = (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_2_sva_mx1[0]) & (FpMul_8U_23U_p_mant_p1_2_sva_mx1[47]))
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_FpMul_8U_23U_and_64_itm_mx0w0 = (mul_loop_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      | (~ (FpMul_8U_23U_p_mant_p1_2_sva_mx1[47]))) & mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign nl_FpMul_8U_23U_else_2_else_acc_3_nl = ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_8_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_8_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_10})
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_3_nl = nl_FpMul_8U_23U_else_2_else_acc_3_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_3_sva_1_mx0w0 = (FpMul_8U_23U_else_2_else_acc_3_nl)
      + (MulIn_data_sva_535[96:89]);
  assign FpMul_8U_23U_p_expo_3_sva_1_mx0w0 = nl_FpMul_8U_23U_p_expo_3_sva_1_mx0w0[7:0];
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_mx0w0 = ~(mul_loop_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      & (mul_loop_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47]));
  assign mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs_mx0w0 = FpMantRNE_48U_24U_else_carry_3_sva_mx0w0
      & (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_3_sva_mx0w0 = (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_3_sva_mx1[0]) & (FpMul_8U_23U_p_mant_p1_3_sva_mx1[47]))
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_FpMul_8U_23U_and_65_itm_mx0w0 = (mul_loop_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      | (~ (FpMul_8U_23U_p_mant_p1_3_sva_mx1[47]))) & mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign nl_FpMul_8U_23U_else_2_else_acc_4_nl = ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_8_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_8_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_10})
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_4_nl = nl_FpMul_8U_23U_else_2_else_acc_4_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_4_sva_1_mx0w0 = (FpMul_8U_23U_else_2_else_acc_4_nl)
      + (MulIn_data_sva_535[129:122]);
  assign FpMul_8U_23U_p_expo_4_sva_1_mx0w0 = nl_FpMul_8U_23U_p_expo_4_sva_1_mx0w0[7:0];
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_mx0w0 = ~(mul_loop_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      & (mul_loop_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47]));
  assign mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs_mx0w0 = FpMantRNE_48U_24U_else_carry_4_sva_mx0w0
      & (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_4_sva_mx0w0 = (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_4_sva_mx1[0]) & (FpMul_8U_23U_p_mant_p1_4_sva_mx1[47]))
      | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_FpMul_8U_23U_and_66_itm_mx0w0 = (mul_loop_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      | (~ (FpMul_8U_23U_p_mant_p1_4_sva_mx1[47]))) & mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign nl_FpMul_8U_23U_else_2_else_acc_5_nl = ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_8_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_8_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_10})
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_5_nl = nl_FpMul_8U_23U_else_2_else_acc_5_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_5_sva_1_mx0w0 = (FpMul_8U_23U_else_2_else_acc_5_nl)
      + (MulIn_data_sva_535[162:155]);
  assign FpMul_8U_23U_p_expo_5_sva_1_mx0w0 = nl_FpMul_8U_23U_p_expo_5_sva_1_mx0w0[7:0];
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_4_itm_mx0w0 = ~(mul_loop_mul_5_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      & (mul_loop_mul_5_FpMul_8U_23U_p_mant_p1_mul_tmp[47]));
  assign mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs_mx0w0 = FpMantRNE_48U_24U_else_carry_5_sva_mx0w0
      & (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_5_sva_mx0w0 = (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_5_sva_mx1[0]) & (FpMul_8U_23U_p_mant_p1_5_sva_mx1[47]))
      | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_FpMul_8U_23U_and_67_itm_mx0w0 = (mul_loop_mul_5_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      | (~ (FpMul_8U_23U_p_mant_p1_5_sva_mx1[47]))) & mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign nl_FpMul_8U_23U_else_2_else_acc_6_nl = ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_8_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_8_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_10})
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_6_nl = nl_FpMul_8U_23U_else_2_else_acc_6_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_6_sva_1_mx0w0 = (FpMul_8U_23U_else_2_else_acc_6_nl)
      + (MulIn_data_sva_535[195:188]);
  assign FpMul_8U_23U_p_expo_6_sva_1_mx0w0 = nl_FpMul_8U_23U_p_expo_6_sva_1_mx0w0[7:0];
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_5_itm_mx0w0 = ~(mul_loop_mul_6_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      & (mul_loop_mul_6_FpMul_8U_23U_p_mant_p1_mul_tmp[47]));
  assign mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs_mx0w0 = FpMantRNE_48U_24U_else_carry_6_sva_mx0w0
      & (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_6_sva_mx0w0 = (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_6_sva_mx1[0]) & (FpMul_8U_23U_p_mant_p1_6_sva_mx1[47]))
      | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_FpMul_8U_23U_and_68_itm_mx0w0 = (mul_loop_mul_6_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      | (~ (FpMul_8U_23U_p_mant_p1_6_sva_mx1[47]))) & mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign nl_FpMul_8U_23U_else_2_else_acc_7_nl = ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_8_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_8_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_10})
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_7_nl = nl_FpMul_8U_23U_else_2_else_acc_7_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_7_sva_1_mx0w0 = (FpMul_8U_23U_else_2_else_acc_7_nl)
      + (MulIn_data_sva_535[228:221]);
  assign FpMul_8U_23U_p_expo_7_sva_1_mx0w0 = nl_FpMul_8U_23U_p_expo_7_sva_1_mx0w0[7:0];
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_6_itm_mx0w0 = ~(mul_loop_mul_7_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      & (mul_loop_mul_7_FpMul_8U_23U_p_mant_p1_mul_tmp[47]));
  assign mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs_mx0w0 = FpMantRNE_48U_24U_else_carry_7_sva_mx0w0
      & (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_7_sva_mx0w0 = (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_7_sva_mx1[0]) & (FpMul_8U_23U_p_mant_p1_7_sva_mx1[47]))
      | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_FpMul_8U_23U_and_69_itm_mx0w0 = (mul_loop_mul_7_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      | (~ (FpMul_8U_23U_p_mant_p1_7_sva_mx1[47]))) & mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign nl_FpMul_8U_23U_else_2_else_acc_8_nl = ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_8_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_8_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_10})
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_8_nl = nl_FpMul_8U_23U_else_2_else_acc_8_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_8_sva_1_mx0w0 = (FpMul_8U_23U_else_2_else_acc_8_nl)
      + (MulIn_data_sva_535[261:254]);
  assign FpMul_8U_23U_p_expo_8_sva_1_mx0w0 = nl_FpMul_8U_23U_p_expo_8_sva_1_mx0w0[7:0];
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_7_itm_mx0w0 = ~(mul_loop_mul_8_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      & (mul_loop_mul_8_FpMul_8U_23U_p_mant_p1_mul_tmp[47]));
  assign mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs_mx0w0 = FpMantRNE_48U_24U_else_carry_8_sva_mx0w0
      & (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_8_sva_mx0w0 = (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_8_sva_mx1[0]) & (FpMul_8U_23U_p_mant_p1_8_sva_mx1[47]))
      | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_FpMul_8U_23U_and_70_itm_mx0w0 = (mul_loop_mul_8_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      | (~ (FpMul_8U_23U_p_mant_p1_8_sva_mx1[47]))) & mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign nl_FpMul_8U_23U_else_2_else_acc_9_nl = ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_8_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_8_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_10})
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_9_nl = nl_FpMul_8U_23U_else_2_else_acc_9_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_9_sva_1_mx0w0 = (FpMul_8U_23U_else_2_else_acc_9_nl)
      + (MulIn_data_sva_535[294:287]);
  assign FpMul_8U_23U_p_expo_9_sva_1_mx0w0 = nl_FpMul_8U_23U_p_expo_9_sva_1_mx0w0[7:0];
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_8_itm_mx0w0 = ~(mul_loop_mul_9_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      & (mul_loop_mul_9_FpMul_8U_23U_p_mant_p1_mul_tmp[47]));
  assign mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs_mx0w0 = FpMantRNE_48U_24U_else_carry_9_sva_mx0w0
      & (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_9_sva_mx0w0 = (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_9_sva_mx1[0]) & (FpMul_8U_23U_p_mant_p1_9_sva_mx1[47]))
      | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_FpMul_8U_23U_and_71_itm_mx0w0 = (mul_loop_mul_9_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      | (~ (FpMul_8U_23U_p_mant_p1_9_sva_mx1[47]))) & mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign nl_FpMul_8U_23U_else_2_else_acc_10_nl = ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_8_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_8_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_10})
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_10_nl = nl_FpMul_8U_23U_else_2_else_acc_10_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_10_sva_1_mx0w0 = (FpMul_8U_23U_else_2_else_acc_10_nl)
      + (MulIn_data_sva_535[327:320]);
  assign FpMul_8U_23U_p_expo_10_sva_1_mx0w0 = nl_FpMul_8U_23U_p_expo_10_sva_1_mx0w0[7:0];
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_9_itm_mx0w0 = ~(mul_loop_mul_10_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      & (mul_loop_mul_10_FpMul_8U_23U_p_mant_p1_mul_tmp[47]));
  assign mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs_mx0w0 = FpMantRNE_48U_24U_else_carry_10_sva_mx0w0
      & (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_10_sva_mx0w0 = (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_10_sva_mx1[0]) & (FpMul_8U_23U_p_mant_p1_10_sva_mx1[47]))
      | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_FpMul_8U_23U_and_72_itm_mx0w0 = (mul_loop_mul_10_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      | (~ (FpMul_8U_23U_p_mant_p1_10_sva_mx1[47]))) & mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign nl_FpMul_8U_23U_else_2_else_acc_11_nl = ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_8_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_8_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_10})
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_11_nl = nl_FpMul_8U_23U_else_2_else_acc_11_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_11_sva_1_mx0w0 = (FpMul_8U_23U_else_2_else_acc_11_nl)
      + (MulIn_data_sva_535[360:353]);
  assign FpMul_8U_23U_p_expo_11_sva_1_mx0w0 = nl_FpMul_8U_23U_p_expo_11_sva_1_mx0w0[7:0];
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_10_itm_mx0w0 = ~(mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      & (mul_loop_mul_11_FpMul_8U_23U_p_mant_p1_mul_tmp[47]));
  assign mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs_mx0w0 = FpMantRNE_48U_24U_else_carry_11_sva_mx0w0
      & (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_11_sva_mx0w0 = (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_11_sva_mx1[0]) & (FpMul_8U_23U_p_mant_p1_11_sva_mx1[47]))
      | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_FpMul_8U_23U_and_73_itm_mx0w0 = (mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      | (~ (FpMul_8U_23U_p_mant_p1_11_sva_mx1[47]))) & mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign nl_FpMul_8U_23U_else_2_else_acc_12_nl = ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_8_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_8_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_10})
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_12_nl = nl_FpMul_8U_23U_else_2_else_acc_12_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_12_sva_1_mx0w0 = (FpMul_8U_23U_else_2_else_acc_12_nl)
      + (MulIn_data_sva_535[393:386]);
  assign FpMul_8U_23U_p_expo_12_sva_1_mx0w0 = nl_FpMul_8U_23U_p_expo_12_sva_1_mx0w0[7:0];
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_11_itm_mx0w0 = ~(mul_loop_mul_12_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      & (mul_loop_mul_12_FpMul_8U_23U_p_mant_p1_mul_tmp[47]));
  assign mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs_mx0w0 = FpMantRNE_48U_24U_else_carry_12_sva_mx0w0
      & (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_12_sva_mx0w0 = (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_12_sva_mx1[0]) & (FpMul_8U_23U_p_mant_p1_12_sva_mx1[47]))
      | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_FpMul_8U_23U_and_74_itm_mx0w0 = (mul_loop_mul_12_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      | (~ (FpMul_8U_23U_p_mant_p1_12_sva_mx1[47]))) & mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign nl_FpMul_8U_23U_else_2_else_acc_13_nl = ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_8_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_8_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_10})
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_13_nl = nl_FpMul_8U_23U_else_2_else_acc_13_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_13_sva_1_mx0w0 = (FpMul_8U_23U_else_2_else_acc_13_nl)
      + (MulIn_data_sva_535[426:419]);
  assign FpMul_8U_23U_p_expo_13_sva_1_mx0w0 = nl_FpMul_8U_23U_p_expo_13_sva_1_mx0w0[7:0];
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_12_itm_mx0w0 = ~(mul_loop_mul_13_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      & (mul_loop_mul_13_FpMul_8U_23U_p_mant_p1_mul_tmp[47]));
  assign mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs_mx0w0 = FpMantRNE_48U_24U_else_carry_13_sva_mx0w0
      & (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_13_sva_mx0w0 = (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_13_sva_mx1[0]) & (FpMul_8U_23U_p_mant_p1_13_sva_mx1[47]))
      | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_FpMul_8U_23U_and_75_itm_mx0w0 = (mul_loop_mul_13_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      | (~ (FpMul_8U_23U_p_mant_p1_13_sva_mx1[47]))) & mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign nl_FpMul_8U_23U_else_2_else_acc_14_nl = ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_8_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_8_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_10})
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_14_nl = nl_FpMul_8U_23U_else_2_else_acc_14_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_14_sva_1_mx0w0 = (FpMul_8U_23U_else_2_else_acc_14_nl)
      + (MulIn_data_sva_535[459:452]);
  assign FpMul_8U_23U_p_expo_14_sva_1_mx0w0 = nl_FpMul_8U_23U_p_expo_14_sva_1_mx0w0[7:0];
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_13_itm_mx0w0 = ~(mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      & (mul_loop_mul_14_FpMul_8U_23U_p_mant_p1_mul_tmp[47]));
  assign mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs_mx0w0 = FpMantRNE_48U_24U_else_carry_14_sva_mx0w0
      & (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_14_sva_mx0w0 = (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_14_sva_mx1[0]) & (FpMul_8U_23U_p_mant_p1_14_sva_mx1[47]))
      | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_FpMul_8U_23U_and_76_itm_mx0w0 = (mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      | (~ (FpMul_8U_23U_p_mant_p1_14_sva_mx1[47]))) & mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign nl_FpMul_8U_23U_else_2_else_acc_15_nl = ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_8_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_8_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_10})
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_15_nl = nl_FpMul_8U_23U_else_2_else_acc_15_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_15_sva_1_mx0w0 = (FpMul_8U_23U_else_2_else_acc_15_nl)
      + (MulIn_data_sva_535[492:485]);
  assign FpMul_8U_23U_p_expo_15_sva_1_mx0w0 = nl_FpMul_8U_23U_p_expo_15_sva_1_mx0w0[7:0];
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_14_itm_mx0w0 = ~(mul_loop_mul_15_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      & (mul_loop_mul_15_FpMul_8U_23U_p_mant_p1_mul_tmp[47]));
  assign mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs_mx0w0 = FpMantRNE_48U_24U_else_carry_15_sva_mx0w0
      & (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_15_sva_mx0w0 = (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_15_sva_mx1[0]) & (FpMul_8U_23U_p_mant_p1_15_sva_mx1[47]))
      | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_FpMul_8U_23U_and_77_itm_mx0w0 = (mul_loop_mul_15_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      | (~ (FpMul_8U_23U_p_mant_p1_15_sva_mx1[47]))) & mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign nl_FpMul_8U_23U_else_2_else_acc_16_nl = ({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_8_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_8_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_10})
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_16_nl = nl_FpMul_8U_23U_else_2_else_acc_16_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_sva_1_mx0w0 = (FpMul_8U_23U_else_2_else_acc_16_nl)
      + (MulIn_data_sva_535[525:518]);
  assign FpMul_8U_23U_p_expo_sva_1_mx0w0 = nl_FpMul_8U_23U_p_expo_sva_1_mx0w0[7:0];
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_15_itm_mx0w0 = ~(mul_loop_mul_16_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      & (mul_loop_mul_16_FpMul_8U_23U_p_mant_p1_mul_tmp[47]));
  assign mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs_mx0w0 = FpMantRNE_48U_24U_else_carry_sva_mx0w0
      & (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_sva_mx0w0 = (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_sva_mx1[0]) & (FpMul_8U_23U_p_mant_p1_sva_mx1[47]))
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_FpMul_8U_23U_and_78_itm_mx0w0 = (mul_loop_mul_16_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7
      | (~ (FpMul_8U_23U_p_mant_p1_sva_mx1[47]))) & mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_177_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_1_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_65_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_177_nl), 10'b1111111111,
      IsInf_5U_23U_land_1_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_239_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_1_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_64_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_239_nl), 10'b1111111111,
      IsInf_5U_23U_land_1_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_nl = MUX_v_3_2_2(3'b000,
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_sva_2[12:10]), (FpExpoWidthInc_5U_8U_23U_1U_1U_not_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_nl),
      3'b111, IsInf_5U_23U_land_1_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_nl),
      3'b111, IsNaN_5U_23U_land_1_lpi_1_dfm));
  assign IsZero_8U_23U_1_land_1_lpi_1_dfm_mx0w0 = (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_9_0_mx1!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_3_2_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_1_0_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_181_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_2_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_68_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_181_nl), 10'b1111111111,
      IsInf_5U_23U_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_145_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_2_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_67_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_145_nl), 10'b1111111111,
      IsInf_5U_23U_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_1_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_66_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_1_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_1_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_66_nl),
      3'b111, IsInf_5U_23U_land_2_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_1_nl),
      3'b111, IsNaN_5U_23U_land_2_lpi_1_dfm));
  assign IsZero_8U_23U_1_land_2_lpi_1_dfm_mx0w0 = (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_9_0_mx1!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_3_2_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_1_0_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_185_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_3_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_71_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_185_nl), 10'b1111111111,
      IsInf_5U_23U_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_147_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_3_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_70_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_147_nl), 10'b1111111111,
      IsInf_5U_23U_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_2_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_68_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_2_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_68_nl),
      3'b111, IsInf_5U_23U_land_3_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_nl),
      3'b111, IsNaN_5U_23U_land_3_lpi_1_dfm));
  assign IsZero_8U_23U_1_land_3_lpi_1_dfm_mx0w0 = (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_9_0_mx1!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_3_2_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_1_0_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_189_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_4_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_74_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_189_nl), 10'b1111111111,
      IsInf_5U_23U_land_4_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_149_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_4_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_73_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_149_nl), 10'b1111111111,
      IsInf_5U_23U_land_4_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_3_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_70_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_3_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_3_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_70_nl),
      3'b111, IsInf_5U_23U_land_4_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_3_nl),
      3'b111, IsNaN_5U_23U_land_4_lpi_1_dfm));
  assign IsZero_8U_23U_1_land_4_lpi_1_dfm_mx0w0 = (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_9_0_mx1!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_3_2_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_1_0_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_193_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_5_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_77_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_193_nl), 10'b1111111111,
      IsInf_5U_23U_land_5_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_151_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_5_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_76_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_151_nl), 10'b1111111111,
      IsInf_5U_23U_land_5_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_4_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_72_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_4_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_72_nl),
      3'b111, IsInf_5U_23U_land_5_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_nl),
      3'b111, IsNaN_5U_23U_land_5_lpi_1_dfm));
  assign IsZero_8U_23U_1_land_5_lpi_1_dfm_mx0w0 = (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_9_0_mx1!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_3_2_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_1_0_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_197_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_6_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_80_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_197_nl), 10'b1111111111,
      IsInf_5U_23U_land_6_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_153_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_6_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_79_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_153_nl), 10'b1111111111,
      IsInf_5U_23U_land_6_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_5_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_74_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_5_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_5_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_74_nl),
      3'b111, IsInf_5U_23U_land_6_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_5_nl),
      3'b111, IsNaN_5U_23U_land_6_lpi_1_dfm));
  assign IsZero_8U_23U_1_land_6_lpi_1_dfm_mx0w0 = (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_9_0_mx1!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_3_2_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_1_0_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_201_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_7_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_83_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_201_nl), 10'b1111111111,
      IsInf_5U_23U_land_7_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_155_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_7_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_82_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_155_nl), 10'b1111111111,
      IsInf_5U_23U_land_7_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_6_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_76_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_6_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_76_nl),
      3'b111, IsInf_5U_23U_land_7_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_nl),
      3'b111, IsNaN_5U_23U_land_7_lpi_1_dfm));
  assign IsZero_8U_23U_1_land_7_lpi_1_dfm_mx0w0 = (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_9_0_mx1!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_3_2_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_1_0_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_205_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_8_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_86_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_205_nl), 10'b1111111111,
      IsInf_5U_23U_land_8_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_157_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_8_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_85_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_157_nl), 10'b1111111111,
      IsInf_5U_23U_land_8_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_7_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_78_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_7_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_7_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_78_nl),
      3'b111, IsInf_5U_23U_land_8_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_7_nl),
      3'b111, IsNaN_5U_23U_land_8_lpi_1_dfm));
  assign IsZero_8U_23U_1_land_8_lpi_1_dfm_mx0w0 = (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_9_0_mx1!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_3_2_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_1_0_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_209_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_9_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_16_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_89_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_209_nl), 10'b1111111111,
      IsInf_5U_23U_land_9_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_159_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_9_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_16_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_88_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_159_nl), 10'b1111111111,
      IsInf_5U_23U_land_9_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_8_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_16_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_80_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_8_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_80_nl),
      3'b111, IsInf_5U_23U_land_9_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_nl),
      3'b111, IsNaN_5U_23U_land_9_lpi_1_dfm));
  assign IsZero_8U_23U_1_land_9_lpi_1_dfm_mx0w0 = (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_9_0_mx1!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_3_2_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_1_0_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_213_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_10_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_18_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_92_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_213_nl), 10'b1111111111,
      IsInf_5U_23U_land_10_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_161_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_10_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_18_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_91_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_161_nl), 10'b1111111111,
      IsInf_5U_23U_land_10_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_9_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_18_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_82_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_9_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_9_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_82_nl),
      3'b111, IsInf_5U_23U_land_10_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_9_nl),
      3'b111, IsNaN_5U_23U_land_10_lpi_1_dfm));
  assign IsZero_8U_23U_1_land_10_lpi_1_dfm_mx0w0 = (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_9_0_mx1!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_3_2_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_1_0_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_217_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_11_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_20_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_95_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_217_nl), 10'b1111111111,
      IsInf_5U_23U_land_11_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_163_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_11_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_20_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_94_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_163_nl), 10'b1111111111,
      IsInf_5U_23U_land_11_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_10_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_20_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_84_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_10_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_84_nl),
      3'b111, IsInf_5U_23U_land_11_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_nl),
      3'b111, IsNaN_5U_23U_land_11_lpi_1_dfm));
  assign IsZero_8U_23U_1_land_11_lpi_1_dfm_mx0w0 = (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_9_0_mx1!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_3_2_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_1_0_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_221_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_12_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_22_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_98_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_221_nl), 10'b1111111111,
      IsInf_5U_23U_land_12_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_165_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_12_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_22_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_97_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_165_nl), 10'b1111111111,
      IsInf_5U_23U_land_12_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_11_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_22_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_86_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_11_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_11_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_86_nl),
      3'b111, IsInf_5U_23U_land_12_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_11_nl),
      3'b111, IsNaN_5U_23U_land_12_lpi_1_dfm));
  assign IsZero_8U_23U_1_land_12_lpi_1_dfm_mx0w0 = (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_9_0_mx1!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_3_2_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_1_0_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_225_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_13_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_24_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_101_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_225_nl), 10'b1111111111,
      IsInf_5U_23U_land_13_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_167_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_13_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_24_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_100_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_167_nl), 10'b1111111111,
      IsInf_5U_23U_land_13_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_12_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_24_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_88_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_12_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_88_nl),
      3'b111, IsInf_5U_23U_land_13_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_nl),
      3'b111, IsNaN_5U_23U_land_13_lpi_1_dfm));
  assign IsZero_8U_23U_1_land_13_lpi_1_dfm_mx0w0 = (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_9_0_mx1!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_3_2_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_1_0_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_229_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_14_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_26_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_104_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_229_nl), 10'b1111111111,
      IsInf_5U_23U_land_14_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_169_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_14_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_26_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_103_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_169_nl), 10'b1111111111,
      IsInf_5U_23U_land_14_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_13_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_26_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_90_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_13_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_13_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_90_nl),
      3'b111, IsInf_5U_23U_land_14_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_13_nl),
      3'b111, IsNaN_5U_23U_land_14_lpi_1_dfm));
  assign IsZero_8U_23U_1_land_14_lpi_1_dfm_mx0w0 = (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_9_0_mx1!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_3_2_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_1_0_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_233_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_15_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_28_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_107_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_233_nl), 10'b1111111111,
      IsInf_5U_23U_land_15_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_171_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_15_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_28_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_106_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_171_nl), 10'b1111111111,
      IsInf_5U_23U_land_15_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_14_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_28_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_92_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_14_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_92_nl),
      3'b111, IsInf_5U_23U_land_15_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_nl),
      3'b111, IsNaN_5U_23U_land_15_lpi_1_dfm));
  assign IsZero_8U_23U_1_land_15_lpi_1_dfm_mx0w0 = (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_9_0_mx1!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_3_2_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_1_0_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_237_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_sva_2[22:13]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_30_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_110_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_237_nl), 10'b1111111111,
      IsInf_5U_23U_land_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_mux_173_nl = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_sva_2[9:0]),
      FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_lpi_1_dfm, FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_30_ssc);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_109_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_mux_173_nl), 10'b1111111111,
      IsInf_5U_23U_land_lpi_1_dfm);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_not_15_nl = ~ FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_30_ssc;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_94_nl
      = MUX_v_3_2_2(3'b000, (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_sva_2[12:10]),
      (FpExpoWidthInc_5U_8U_23U_1U_1U_not_15_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_nor_15_nl = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_and_94_nl),
      3'b111, IsInf_5U_23U_land_lpi_1_dfm));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_12_10_mx0w0 = ~(MUX_v_3_2_2((FpExpoWidthInc_5U_8U_23U_1U_1U_nor_15_nl),
      3'b111, IsNaN_5U_23U_land_lpi_1_dfm));
  assign IsZero_8U_23U_1_land_lpi_1_dfm_mx0w0 = (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_12_10_mx0w0!=3'b000) |
      (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_9_0_mx1!=10'b0000000000)))
      & (~((FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_3_2_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_1_0_mx0w0!=2'b00)
      | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign IsZero_8U_23U_land_1_lpi_1_dfm_mx0w0 = ~((chn_mul_in_rsci_d_mxwt[30:0]!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_land_2_lpi_1_dfm_mx0w0 = ~((chn_mul_in_rsci_d_mxwt[63:33]!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_land_3_lpi_1_dfm_mx0w0 = ~((chn_mul_in_rsci_d_mxwt[96:66]!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_land_4_lpi_1_dfm_mx0w0 = ~((chn_mul_in_rsci_d_mxwt[129:99]!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_land_5_lpi_1_dfm_mx0w0 = ~((chn_mul_in_rsci_d_mxwt[162:132]!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_land_6_lpi_1_dfm_mx0w0 = ~((chn_mul_in_rsci_d_mxwt[195:165]!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_land_7_lpi_1_dfm_mx0w0 = ~((chn_mul_in_rsci_d_mxwt[228:198]!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_land_8_lpi_1_dfm_mx0w0 = ~((chn_mul_in_rsci_d_mxwt[261:231]!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_land_9_lpi_1_dfm_mx0w0 = ~((chn_mul_in_rsci_d_mxwt[294:264]!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_land_10_lpi_1_dfm_mx0w0 = ~((chn_mul_in_rsci_d_mxwt[327:297]!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_land_11_lpi_1_dfm_mx0w0 = ~((chn_mul_in_rsci_d_mxwt[360:330]!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_land_12_lpi_1_dfm_mx0w0 = ~((chn_mul_in_rsci_d_mxwt[393:363]!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_land_13_lpi_1_dfm_mx0w0 = ~((chn_mul_in_rsci_d_mxwt[426:396]!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_land_14_lpi_1_dfm_mx0w0 = ~((chn_mul_in_rsci_d_mxwt[459:429]!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_land_15_lpi_1_dfm_mx0w0 = ~((chn_mul_in_rsci_d_mxwt[492:462]!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_land_lpi_1_dfm_mx0w0 = ~((chn_mul_in_rsci_d_mxwt[525:495]!=31'b0000000000000000000000000000000));
  assign mul_loop_mul_16_FpMul_8U_23U_xor_nl = (MulIn_data_sva_534[526]) ^ mul_nan_to_zero_op_sign_lpi_1_dfm_4;
  assign FpMul_8U_23U_else_5_mux_60_mx0w1 = MUX_s_1_2_2((mul_loop_mul_16_FpMul_8U_23U_xor_nl),
      mul_nan_to_zero_op_sign_lpi_1_dfm_4, IsNaN_8U_23U_1_land_lpi_1_dfm_7);
  assign mul_loop_mul_15_FpMul_8U_23U_xor_nl = (MulIn_data_sva_534[493]) ^ mul_nan_to_zero_op_sign_15_lpi_1_dfm_4;
  assign FpMul_8U_23U_else_5_mux_56_mx0w1 = MUX_s_1_2_2((mul_loop_mul_15_FpMul_8U_23U_xor_nl),
      mul_nan_to_zero_op_sign_15_lpi_1_dfm_4, IsNaN_8U_23U_1_land_15_lpi_1_dfm_7);
  assign mul_loop_mul_14_FpMul_8U_23U_xor_nl = (MulIn_data_sva_534[460]) ^ mul_nan_to_zero_op_sign_14_lpi_1_dfm_4;
  assign FpMul_8U_23U_else_5_mux_52_mx0w1 = MUX_s_1_2_2((mul_loop_mul_14_FpMul_8U_23U_xor_nl),
      mul_nan_to_zero_op_sign_14_lpi_1_dfm_4, IsNaN_8U_23U_1_land_14_lpi_1_dfm_7);
  assign mul_loop_mul_13_FpMul_8U_23U_xor_nl = (MulIn_data_sva_534[427]) ^ mul_nan_to_zero_op_sign_13_lpi_1_dfm_4;
  assign FpMul_8U_23U_else_5_mux_48_mx0w1 = MUX_s_1_2_2((mul_loop_mul_13_FpMul_8U_23U_xor_nl),
      mul_nan_to_zero_op_sign_13_lpi_1_dfm_4, IsNaN_8U_23U_1_land_13_lpi_1_dfm_7);
  assign mul_loop_mul_12_FpMul_8U_23U_xor_nl = (MulIn_data_sva_534[394]) ^ mul_nan_to_zero_op_sign_12_lpi_1_dfm_4;
  assign FpMul_8U_23U_else_5_mux_44_mx0w1 = MUX_s_1_2_2((mul_loop_mul_12_FpMul_8U_23U_xor_nl),
      mul_nan_to_zero_op_sign_12_lpi_1_dfm_4, IsNaN_8U_23U_1_land_12_lpi_1_dfm_7);
  assign mul_loop_mul_11_FpMul_8U_23U_xor_nl = (MulIn_data_sva_534[361]) ^ mul_nan_to_zero_op_sign_11_lpi_1_dfm_4;
  assign FpMul_8U_23U_else_5_mux_40_mx0w1 = MUX_s_1_2_2((mul_loop_mul_11_FpMul_8U_23U_xor_nl),
      mul_nan_to_zero_op_sign_11_lpi_1_dfm_4, IsNaN_8U_23U_1_land_11_lpi_1_dfm_7);
  assign FpMul_8U_23U_lor_27_lpi_1_dfm_mx0w0 = mul_loop_mul_10_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | reg_FpMul_8U_23U_lor_12_lpi_1_dfm_4_cse;
  assign mul_loop_mul_10_FpMul_8U_23U_xor_nl = (MulIn_data_sva_534[328]) ^ mul_nan_to_zero_op_sign_10_lpi_1_dfm_4;
  assign FpMul_8U_23U_else_5_mux_36_mx0w1 = MUX_s_1_2_2((mul_loop_mul_10_FpMul_8U_23U_xor_nl),
      mul_nan_to_zero_op_sign_10_lpi_1_dfm_4, IsNaN_8U_23U_1_land_10_lpi_1_dfm_7);
  assign FpMul_8U_23U_lor_26_lpi_1_dfm_mx0w0 = mul_loop_mul_9_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | reg_FpMul_8U_23U_lor_11_lpi_1_dfm_4_cse;
  assign mul_loop_mul_9_FpMul_8U_23U_xor_nl = (MulIn_data_sva_534[295]) ^ mul_nan_to_zero_op_sign_9_lpi_1_dfm_4;
  assign FpMul_8U_23U_else_5_mux_32_mx0w1 = MUX_s_1_2_2((mul_loop_mul_9_FpMul_8U_23U_xor_nl),
      mul_nan_to_zero_op_sign_9_lpi_1_dfm_4, IsNaN_8U_23U_1_land_9_lpi_1_dfm_7);
  assign mul_loop_mul_8_FpMul_8U_23U_xor_nl = (MulIn_data_sva_534[262]) ^ mul_nan_to_zero_op_sign_8_lpi_1_dfm_4;
  assign FpMul_8U_23U_else_5_mux_28_mx0w1 = MUX_s_1_2_2((mul_loop_mul_8_FpMul_8U_23U_xor_nl),
      mul_nan_to_zero_op_sign_8_lpi_1_dfm_4, IsNaN_8U_23U_1_land_8_lpi_1_dfm_7);
  assign mul_loop_mul_7_FpMul_8U_23U_xor_nl = (MulIn_data_sva_534[229]) ^ mul_nan_to_zero_op_sign_7_lpi_1_dfm_4;
  assign FpMul_8U_23U_else_5_mux_24_mx0w1 = MUX_s_1_2_2((mul_loop_mul_7_FpMul_8U_23U_xor_nl),
      mul_nan_to_zero_op_sign_7_lpi_1_dfm_4, IsNaN_8U_23U_1_land_7_lpi_1_dfm_7);
  assign mul_loop_mul_6_FpMul_8U_23U_xor_nl = (MulIn_data_sva_534[196]) ^ mul_nan_to_zero_op_sign_6_lpi_1_dfm_4;
  assign FpMul_8U_23U_else_5_mux_20_mx0w1 = MUX_s_1_2_2((mul_loop_mul_6_FpMul_8U_23U_xor_nl),
      mul_nan_to_zero_op_sign_6_lpi_1_dfm_4, IsNaN_8U_23U_1_land_6_lpi_1_dfm_7);
  assign FpMul_8U_23U_lor_22_lpi_1_dfm_mx0w0 = mul_loop_mul_5_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | reg_FpMul_8U_23U_lor_7_lpi_1_dfm_4_cse;
  assign mul_loop_mul_5_FpMul_8U_23U_xor_nl = (MulIn_data_sva_534[163]) ^ mul_nan_to_zero_op_sign_5_lpi_1_dfm_4;
  assign FpMul_8U_23U_else_5_mux_16_mx0w1 = MUX_s_1_2_2((mul_loop_mul_5_FpMul_8U_23U_xor_nl),
      mul_nan_to_zero_op_sign_5_lpi_1_dfm_4, IsNaN_8U_23U_1_land_5_lpi_1_dfm_7);
  assign mul_loop_mul_4_FpMul_8U_23U_xor_nl = (MulIn_data_sva_534[130]) ^ mul_nan_to_zero_op_sign_4_lpi_1_dfm_4;
  assign FpMul_8U_23U_else_5_mux_12_mx0w1 = MUX_s_1_2_2((mul_loop_mul_4_FpMul_8U_23U_xor_nl),
      mul_nan_to_zero_op_sign_4_lpi_1_dfm_4, IsNaN_8U_23U_1_land_4_lpi_1_dfm_7);
  assign mul_loop_mul_3_FpMul_8U_23U_xor_nl = (MulIn_data_sva_534[97]) ^ mul_nan_to_zero_op_sign_3_lpi_1_dfm_4;
  assign FpMul_8U_23U_else_5_mux_8_mx0w1 = MUX_s_1_2_2((mul_loop_mul_3_FpMul_8U_23U_xor_nl),
      mul_nan_to_zero_op_sign_3_lpi_1_dfm_4, IsNaN_8U_23U_1_land_3_lpi_1_dfm_7);
  assign mul_loop_mul_2_FpMul_8U_23U_xor_nl = (MulIn_data_sva_534[64]) ^ mul_nan_to_zero_op_sign_2_lpi_1_dfm_4;
  assign FpMul_8U_23U_else_5_mux_4_mx0w1 = MUX_s_1_2_2((mul_loop_mul_2_FpMul_8U_23U_xor_nl),
      mul_nan_to_zero_op_sign_2_lpi_1_dfm_4, IsNaN_8U_23U_1_land_2_lpi_1_dfm_7);
  assign mul_loop_mul_1_FpMul_8U_23U_xor_nl = (MulIn_data_sva_534[31]) ^ mul_nan_to_zero_op_sign_1_lpi_1_dfm_4;
  assign FpMul_8U_23U_else_5_mux_mx0w1 = MUX_s_1_2_2((mul_loop_mul_1_FpMul_8U_23U_xor_nl),
      mul_nan_to_zero_op_sign_1_lpi_1_dfm_4, IsNaN_8U_23U_1_land_1_lpi_1_dfm_7);
  assign FpMul_8U_23U_p_mant_p1_and_31_nl = mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & (~ FpMul_8U_23U_lor_18_lpi_1_dfm_st_3);
  assign FpMul_8U_23U_p_mant_p1_1_sva_mx1 = MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_1_sva,
      mul_loop_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp, FpMul_8U_23U_p_mant_p1_and_31_nl);
  assign mul_loop_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({(~ IsZero_8U_23U_land_1_lpi_1_dfm_8)
      , (MulIn_data_sva_535[22:0])}) * ({(~ IsZero_8U_23U_1_land_1_lpi_1_dfm_7) ,
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_22_13_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_12_10_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_9_0_1}));
  assign nl_mul_loop_mul_1_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(MulIn_data_sva_534[30:23])
      + conv_u2u_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_9});
  assign mul_loop_mul_1_FpMul_8U_23U_else_2_acc_1_nl = nl_mul_loop_mul_1_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_mul_loop_mul_1_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(readslicef_9_8_1((mul_loop_mul_1_FpMul_8U_23U_else_2_acc_1_nl)))
      + 9'b101000001;
  assign mul_loop_mul_1_FpMul_8U_23U_else_2_if_acc_nl = nl_mul_loop_mul_1_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign mul_loop_mul_1_FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((mul_loop_mul_1_FpMul_8U_23U_else_2_if_acc_nl));
  assign FpMul_8U_23U_p_mant_p1_and_30_nl = mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & (~ FpMul_8U_23U_lor_19_lpi_1_dfm_st_3);
  assign FpMul_8U_23U_p_mant_p1_2_sva_mx1 = MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_2_sva,
      mul_loop_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp, FpMul_8U_23U_p_mant_p1_and_30_nl);
  assign mul_loop_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({(~ IsZero_8U_23U_land_2_lpi_1_dfm_8)
      , (MulIn_data_sva_535[55:33])}) * ({(~ IsZero_8U_23U_1_land_2_lpi_1_dfm_7)
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_22_13_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_12_10_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_9_0_1}));
  assign nl_mul_loop_mul_2_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(MulIn_data_sva_534[63:56])
      + conv_u2u_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_9});
  assign mul_loop_mul_2_FpMul_8U_23U_else_2_acc_1_nl = nl_mul_loop_mul_2_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_mul_loop_mul_2_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(readslicef_9_8_1((mul_loop_mul_2_FpMul_8U_23U_else_2_acc_1_nl)))
      + 9'b101000001;
  assign mul_loop_mul_2_FpMul_8U_23U_else_2_if_acc_nl = nl_mul_loop_mul_2_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign mul_loop_mul_2_FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((mul_loop_mul_2_FpMul_8U_23U_else_2_if_acc_nl));
  assign FpMul_8U_23U_p_mant_p1_and_29_nl = mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & (~ FpMul_8U_23U_lor_20_lpi_1_dfm_st_3);
  assign FpMul_8U_23U_p_mant_p1_3_sva_mx1 = MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_3_sva,
      mul_loop_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp, FpMul_8U_23U_p_mant_p1_and_29_nl);
  assign mul_loop_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({(~ IsZero_8U_23U_land_3_lpi_1_dfm_8)
      , (MulIn_data_sva_535[88:66])}) * ({(~ IsZero_8U_23U_1_land_3_lpi_1_dfm_7)
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_22_13_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_12_10_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_9_0_1}));
  assign nl_mul_loop_mul_3_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(MulIn_data_sva_534[96:89])
      + conv_u2u_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_9});
  assign mul_loop_mul_3_FpMul_8U_23U_else_2_acc_1_nl = nl_mul_loop_mul_3_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_mul_loop_mul_3_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(readslicef_9_8_1((mul_loop_mul_3_FpMul_8U_23U_else_2_acc_1_nl)))
      + 9'b101000001;
  assign mul_loop_mul_3_FpMul_8U_23U_else_2_if_acc_nl = nl_mul_loop_mul_3_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign mul_loop_mul_3_FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((mul_loop_mul_3_FpMul_8U_23U_else_2_if_acc_nl));
  assign FpMul_8U_23U_p_mant_p1_and_28_nl = mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & (~ FpMul_8U_23U_lor_21_lpi_1_dfm_st_3);
  assign FpMul_8U_23U_p_mant_p1_4_sva_mx1 = MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_4_sva,
      mul_loop_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp, FpMul_8U_23U_p_mant_p1_and_28_nl);
  assign mul_loop_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({(~ IsZero_8U_23U_land_4_lpi_1_dfm_8)
      , (MulIn_data_sva_535[121:99])}) * ({(~ IsZero_8U_23U_1_land_4_lpi_1_dfm_6)
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_22_13_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_12_10_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_9_0_1}));
  assign nl_mul_loop_mul_4_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(MulIn_data_sva_534[129:122])
      + conv_u2u_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_9});
  assign mul_loop_mul_4_FpMul_8U_23U_else_2_acc_1_nl = nl_mul_loop_mul_4_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_mul_loop_mul_4_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(readslicef_9_8_1((mul_loop_mul_4_FpMul_8U_23U_else_2_acc_1_nl)))
      + 9'b101000001;
  assign mul_loop_mul_4_FpMul_8U_23U_else_2_if_acc_nl = nl_mul_loop_mul_4_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign mul_loop_mul_4_FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((mul_loop_mul_4_FpMul_8U_23U_else_2_if_acc_nl));
  assign FpMul_8U_23U_p_mant_p1_and_27_nl = mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & (~ FpMul_8U_23U_lor_22_lpi_1_dfm_st_3);
  assign FpMul_8U_23U_p_mant_p1_5_sva_mx1 = MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_5_sva,
      mul_loop_mul_5_FpMul_8U_23U_p_mant_p1_mul_tmp, FpMul_8U_23U_p_mant_p1_and_27_nl);
  assign mul_loop_mul_5_FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({(~ IsZero_8U_23U_land_5_lpi_1_dfm_8)
      , (MulIn_data_sva_535[154:132])}) * ({(~ IsZero_8U_23U_1_land_5_lpi_1_dfm_7)
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_22_13_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_12_10_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_9_0_1}));
  assign nl_mul_loop_mul_5_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(MulIn_data_sva_534[162:155])
      + conv_u2u_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_9});
  assign mul_loop_mul_5_FpMul_8U_23U_else_2_acc_1_nl = nl_mul_loop_mul_5_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_mul_loop_mul_5_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(readslicef_9_8_1((mul_loop_mul_5_FpMul_8U_23U_else_2_acc_1_nl)))
      + 9'b101000001;
  assign mul_loop_mul_5_FpMul_8U_23U_else_2_if_acc_nl = nl_mul_loop_mul_5_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign mul_loop_mul_5_FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((mul_loop_mul_5_FpMul_8U_23U_else_2_if_acc_nl));
  assign FpMul_8U_23U_p_mant_p1_and_26_nl = mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & (~ FpMul_8U_23U_lor_23_lpi_1_dfm_st_3);
  assign FpMul_8U_23U_p_mant_p1_6_sva_mx1 = MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_6_sva,
      mul_loop_mul_6_FpMul_8U_23U_p_mant_p1_mul_tmp, FpMul_8U_23U_p_mant_p1_and_26_nl);
  assign mul_loop_mul_6_FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({(~ IsZero_8U_23U_land_6_lpi_1_dfm_8)
      , (MulIn_data_sva_535[187:165])}) * ({(~ IsZero_8U_23U_1_land_6_lpi_1_dfm_6)
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_22_13_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_12_10_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_9_0_1}));
  assign nl_mul_loop_mul_6_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(MulIn_data_sva_534[195:188])
      + conv_u2u_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_9});
  assign mul_loop_mul_6_FpMul_8U_23U_else_2_acc_1_nl = nl_mul_loop_mul_6_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_mul_loop_mul_6_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(readslicef_9_8_1((mul_loop_mul_6_FpMul_8U_23U_else_2_acc_1_nl)))
      + 9'b101000001;
  assign mul_loop_mul_6_FpMul_8U_23U_else_2_if_acc_nl = nl_mul_loop_mul_6_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign mul_loop_mul_6_FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((mul_loop_mul_6_FpMul_8U_23U_else_2_if_acc_nl));
  assign FpMul_8U_23U_p_mant_p1_and_25_nl = mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & (~ FpMul_8U_23U_lor_24_lpi_1_dfm_st_3);
  assign FpMul_8U_23U_p_mant_p1_7_sva_mx1 = MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_7_sva,
      mul_loop_mul_7_FpMul_8U_23U_p_mant_p1_mul_tmp, FpMul_8U_23U_p_mant_p1_and_25_nl);
  assign mul_loop_mul_7_FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({(~ IsZero_8U_23U_land_7_lpi_1_dfm_8)
      , (MulIn_data_sva_535[220:198])}) * ({(~ IsZero_8U_23U_1_land_7_lpi_1_dfm_6)
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_22_13_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_12_10_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_9_0_1}));
  assign nl_mul_loop_mul_7_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(MulIn_data_sva_534[228:221])
      + conv_u2u_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_9});
  assign mul_loop_mul_7_FpMul_8U_23U_else_2_acc_1_nl = nl_mul_loop_mul_7_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_mul_loop_mul_7_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(readslicef_9_8_1((mul_loop_mul_7_FpMul_8U_23U_else_2_acc_1_nl)))
      + 9'b101000001;
  assign mul_loop_mul_7_FpMul_8U_23U_else_2_if_acc_nl = nl_mul_loop_mul_7_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign mul_loop_mul_7_FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((mul_loop_mul_7_FpMul_8U_23U_else_2_if_acc_nl));
  assign FpMul_8U_23U_p_mant_p1_and_24_nl = mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & (~ FpMul_8U_23U_lor_25_lpi_1_dfm_st_3);
  assign FpMul_8U_23U_p_mant_p1_8_sva_mx1 = MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_8_sva,
      mul_loop_mul_8_FpMul_8U_23U_p_mant_p1_mul_tmp, FpMul_8U_23U_p_mant_p1_and_24_nl);
  assign mul_loop_mul_8_FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({(~ IsZero_8U_23U_land_8_lpi_1_dfm_8)
      , (MulIn_data_sva_535[253:231])}) * ({(~ IsZero_8U_23U_1_land_8_lpi_1_dfm_7)
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_22_13_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_12_10_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_9_0_1}));
  assign nl_mul_loop_mul_8_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(MulIn_data_sva_534[261:254])
      + conv_u2u_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_9});
  assign mul_loop_mul_8_FpMul_8U_23U_else_2_acc_1_nl = nl_mul_loop_mul_8_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_mul_loop_mul_8_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(readslicef_9_8_1((mul_loop_mul_8_FpMul_8U_23U_else_2_acc_1_nl)))
      + 9'b101000001;
  assign mul_loop_mul_8_FpMul_8U_23U_else_2_if_acc_nl = nl_mul_loop_mul_8_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign mul_loop_mul_8_FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((mul_loop_mul_8_FpMul_8U_23U_else_2_if_acc_nl));
  assign FpMul_8U_23U_p_mant_p1_and_23_nl = mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & (~ FpMul_8U_23U_lor_26_lpi_1_dfm_st_3);
  assign FpMul_8U_23U_p_mant_p1_9_sva_mx1 = MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_9_sva,
      mul_loop_mul_9_FpMul_8U_23U_p_mant_p1_mul_tmp, FpMul_8U_23U_p_mant_p1_and_23_nl);
  assign mul_loop_mul_9_FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({(~ IsZero_8U_23U_land_9_lpi_1_dfm_8)
      , (MulIn_data_sva_535[286:264])}) * ({(~ IsZero_8U_23U_1_land_9_lpi_1_dfm_7)
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_22_13_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_12_10_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_9_0_1}));
  assign nl_mul_loop_mul_9_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(MulIn_data_sva_534[294:287])
      + conv_u2u_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_9});
  assign mul_loop_mul_9_FpMul_8U_23U_else_2_acc_1_nl = nl_mul_loop_mul_9_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_mul_loop_mul_9_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(readslicef_9_8_1((mul_loop_mul_9_FpMul_8U_23U_else_2_acc_1_nl)))
      + 9'b101000001;
  assign mul_loop_mul_9_FpMul_8U_23U_else_2_if_acc_nl = nl_mul_loop_mul_9_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign mul_loop_mul_9_FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((mul_loop_mul_9_FpMul_8U_23U_else_2_if_acc_nl));
  assign FpMul_8U_23U_p_mant_p1_and_22_nl = mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & (~ FpMul_8U_23U_lor_27_lpi_1_dfm_st_3);
  assign FpMul_8U_23U_p_mant_p1_10_sva_mx1 = MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_10_sva,
      mul_loop_mul_10_FpMul_8U_23U_p_mant_p1_mul_tmp, FpMul_8U_23U_p_mant_p1_and_22_nl);
  assign mul_loop_mul_10_FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({(~ IsZero_8U_23U_land_10_lpi_1_dfm_8)
      , (MulIn_data_sva_535[319:297])}) * ({(~ IsZero_8U_23U_1_land_10_lpi_1_dfm_6)
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_22_13_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_12_10_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_9_0_1}));
  assign nl_mul_loop_mul_10_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(MulIn_data_sva_534[327:320])
      + conv_u2u_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_9});
  assign mul_loop_mul_10_FpMul_8U_23U_else_2_acc_1_nl = nl_mul_loop_mul_10_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_mul_loop_mul_10_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(readslicef_9_8_1((mul_loop_mul_10_FpMul_8U_23U_else_2_acc_1_nl)))
      + 9'b101000001;
  assign mul_loop_mul_10_FpMul_8U_23U_else_2_if_acc_nl = nl_mul_loop_mul_10_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign mul_loop_mul_10_FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((mul_loop_mul_10_FpMul_8U_23U_else_2_if_acc_nl));
  assign FpMul_8U_23U_p_mant_p1_and_21_nl = mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & (~ FpMul_8U_23U_lor_28_lpi_1_dfm_st_3);
  assign FpMul_8U_23U_p_mant_p1_11_sva_mx1 = MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_11_sva,
      mul_loop_mul_11_FpMul_8U_23U_p_mant_p1_mul_tmp, FpMul_8U_23U_p_mant_p1_and_21_nl);
  assign mul_loop_mul_11_FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({(~ IsZero_8U_23U_land_11_lpi_1_dfm_8)
      , (MulIn_data_sva_535[352:330])}) * ({(~ IsZero_8U_23U_1_land_11_lpi_1_dfm_6)
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_22_13_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_12_10_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_9_0_1}));
  assign nl_mul_loop_mul_11_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(MulIn_data_sva_534[360:353])
      + conv_u2u_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_9});
  assign mul_loop_mul_11_FpMul_8U_23U_else_2_acc_1_nl = nl_mul_loop_mul_11_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_mul_loop_mul_11_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(readslicef_9_8_1((mul_loop_mul_11_FpMul_8U_23U_else_2_acc_1_nl)))
      + 9'b101000001;
  assign mul_loop_mul_11_FpMul_8U_23U_else_2_if_acc_nl = nl_mul_loop_mul_11_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign mul_loop_mul_11_FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((mul_loop_mul_11_FpMul_8U_23U_else_2_if_acc_nl));
  assign FpMul_8U_23U_p_mant_p1_and_20_nl = mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & (~ FpMul_8U_23U_lor_29_lpi_1_dfm_st_3);
  assign FpMul_8U_23U_p_mant_p1_12_sva_mx1 = MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_12_sva,
      mul_loop_mul_12_FpMul_8U_23U_p_mant_p1_mul_tmp, FpMul_8U_23U_p_mant_p1_and_20_nl);
  assign mul_loop_mul_12_FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({(~ IsZero_8U_23U_land_12_lpi_1_dfm_8)
      , (MulIn_data_sva_535[385:363])}) * ({(~ IsZero_8U_23U_1_land_12_lpi_1_dfm_6)
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_22_13_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_12_10_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_9_0_1}));
  assign nl_mul_loop_mul_12_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(MulIn_data_sva_534[393:386])
      + conv_u2u_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_9});
  assign mul_loop_mul_12_FpMul_8U_23U_else_2_acc_1_nl = nl_mul_loop_mul_12_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_mul_loop_mul_12_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(readslicef_9_8_1((mul_loop_mul_12_FpMul_8U_23U_else_2_acc_1_nl)))
      + 9'b101000001;
  assign mul_loop_mul_12_FpMul_8U_23U_else_2_if_acc_nl = nl_mul_loop_mul_12_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign mul_loop_mul_12_FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((mul_loop_mul_12_FpMul_8U_23U_else_2_if_acc_nl));
  assign FpMul_8U_23U_p_mant_p1_and_19_nl = mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & (~ FpMul_8U_23U_lor_30_lpi_1_dfm_st_3);
  assign FpMul_8U_23U_p_mant_p1_13_sva_mx1 = MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_13_sva,
      mul_loop_mul_13_FpMul_8U_23U_p_mant_p1_mul_tmp, FpMul_8U_23U_p_mant_p1_and_19_nl);
  assign mul_loop_mul_13_FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({(~ IsZero_8U_23U_land_13_lpi_1_dfm_8)
      , (MulIn_data_sva_535[418:396])}) * ({(~ IsZero_8U_23U_1_land_13_lpi_1_dfm_7)
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_22_13_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_12_10_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_9_0_1}));
  assign nl_mul_loop_mul_13_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(MulIn_data_sva_534[426:419])
      + conv_u2u_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_9});
  assign mul_loop_mul_13_FpMul_8U_23U_else_2_acc_1_nl = nl_mul_loop_mul_13_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_mul_loop_mul_13_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(readslicef_9_8_1((mul_loop_mul_13_FpMul_8U_23U_else_2_acc_1_nl)))
      + 9'b101000001;
  assign mul_loop_mul_13_FpMul_8U_23U_else_2_if_acc_nl = nl_mul_loop_mul_13_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign mul_loop_mul_13_FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((mul_loop_mul_13_FpMul_8U_23U_else_2_if_acc_nl));
  assign FpMul_8U_23U_p_mant_p1_and_18_nl = mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & (~ FpMul_8U_23U_lor_31_lpi_1_dfm_st_3);
  assign FpMul_8U_23U_p_mant_p1_14_sva_mx1 = MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_14_sva,
      mul_loop_mul_14_FpMul_8U_23U_p_mant_p1_mul_tmp, FpMul_8U_23U_p_mant_p1_and_18_nl);
  assign mul_loop_mul_14_FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({(~ IsZero_8U_23U_land_14_lpi_1_dfm_8)
      , (MulIn_data_sva_535[451:429])}) * ({(~ IsZero_8U_23U_1_land_14_lpi_1_dfm_6)
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_22_13_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_12_10_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_9_0_1}));
  assign nl_mul_loop_mul_14_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(MulIn_data_sva_534[459:452])
      + conv_u2u_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_9});
  assign mul_loop_mul_14_FpMul_8U_23U_else_2_acc_1_nl = nl_mul_loop_mul_14_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_mul_loop_mul_14_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(readslicef_9_8_1((mul_loop_mul_14_FpMul_8U_23U_else_2_acc_1_nl)))
      + 9'b101000001;
  assign mul_loop_mul_14_FpMul_8U_23U_else_2_if_acc_nl = nl_mul_loop_mul_14_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign mul_loop_mul_14_FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((mul_loop_mul_14_FpMul_8U_23U_else_2_if_acc_nl));
  assign FpMul_8U_23U_p_mant_p1_and_17_nl = mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & (~ FpMul_8U_23U_lor_32_lpi_1_dfm_st_3);
  assign FpMul_8U_23U_p_mant_p1_15_sva_mx1 = MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_15_sva,
      mul_loop_mul_15_FpMul_8U_23U_p_mant_p1_mul_tmp, FpMul_8U_23U_p_mant_p1_and_17_nl);
  assign mul_loop_mul_15_FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({(~ IsZero_8U_23U_land_15_lpi_1_dfm_8)
      , (MulIn_data_sva_535[484:462])}) * ({(~ IsZero_8U_23U_1_land_15_lpi_1_dfm_7)
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_22_13_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_12_10_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_9_0_1}));
  assign nl_mul_loop_mul_15_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(MulIn_data_sva_534[492:485])
      + conv_u2u_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_9});
  assign mul_loop_mul_15_FpMul_8U_23U_else_2_acc_1_nl = nl_mul_loop_mul_15_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_mul_loop_mul_15_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(readslicef_9_8_1((mul_loop_mul_15_FpMul_8U_23U_else_2_acc_1_nl)))
      + 9'b101000001;
  assign mul_loop_mul_15_FpMul_8U_23U_else_2_if_acc_nl = nl_mul_loop_mul_15_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign mul_loop_mul_15_FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((mul_loop_mul_15_FpMul_8U_23U_else_2_if_acc_nl));
  assign FpMul_8U_23U_p_mant_p1_and_16_nl = mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & (~ FpMul_8U_23U_lor_1_lpi_1_dfm_st_3);
  assign FpMul_8U_23U_p_mant_p1_sva_mx1 = MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_sva,
      mul_loop_mul_16_FpMul_8U_23U_p_mant_p1_mul_tmp, FpMul_8U_23U_p_mant_p1_and_16_nl);
  assign mul_loop_mul_16_FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({(~ IsZero_8U_23U_land_lpi_1_dfm_8)
      , (MulIn_data_sva_535[517:495])}) * ({(~ IsZero_8U_23U_1_land_lpi_1_dfm_7)
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_22_13_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_12_10_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_9_0_1}));
  assign nl_mul_loop_mul_16_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(MulIn_data_sva_534[525:518])
      + conv_u2u_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_9});
  assign mul_loop_mul_16_FpMul_8U_23U_else_2_acc_1_nl = nl_mul_loop_mul_16_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_mul_loop_mul_16_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(readslicef_9_8_1((mul_loop_mul_16_FpMul_8U_23U_else_2_acc_1_nl)))
      + 9'b101000001;
  assign mul_loop_mul_16_FpMul_8U_23U_else_2_if_acc_nl = nl_mul_loop_mul_16_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign mul_loop_mul_16_FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((mul_loop_mul_16_FpMul_8U_23U_else_2_if_acc_nl));
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_22_13_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_1_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_65_mx0w1,
      or_dcpl_212);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_9_0_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_1_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_64_mx0w1,
      or_dcpl_212);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_22_13_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_2_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_68_mx0w1,
      or_dcpl_224);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_9_0_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_2_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_67_mx0w1,
      or_dcpl_224);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_22_13_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_3_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_71_mx0w1,
      or_dcpl_234);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_9_0_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_3_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_70_mx0w1,
      or_dcpl_234);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_22_13_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_4_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_74_mx0w1,
      or_dcpl_244);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_9_0_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_4_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_73_mx0w1,
      or_dcpl_244);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_22_13_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_5_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_77_mx0w1,
      or_dcpl_254);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_9_0_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_5_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_76_mx0w1,
      or_dcpl_254);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_22_13_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_6_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_80_mx0w1,
      or_dcpl_264);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_9_0_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_6_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_79_mx0w1,
      or_dcpl_264);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_22_13_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_7_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_83_mx0w1,
      or_dcpl_274);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_9_0_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_7_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_82_mx0w1,
      or_dcpl_274);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_22_13_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_8_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_86_mx0w1,
      or_dcpl_284);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_9_0_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_8_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_85_mx0w1,
      or_dcpl_284);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_22_13_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_9_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_89_mx0w1,
      or_dcpl_294);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_9_0_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_9_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_88_mx0w1,
      or_dcpl_294);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_22_13_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_10_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_92_mx0w1,
      or_dcpl_304);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_9_0_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_10_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_91_mx0w1,
      or_dcpl_304);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_22_13_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_11_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_95_mx0w1,
      or_dcpl_314);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_9_0_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_11_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_94_mx0w1,
      or_dcpl_314);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_22_13_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_12_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_98_mx0w1,
      or_dcpl_324);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_9_0_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_12_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_97_mx0w1,
      or_dcpl_324);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_22_13_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_13_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_101_mx0w1,
      or_dcpl_334);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_9_0_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_13_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_100_mx0w1,
      or_dcpl_334);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_22_13_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_14_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_104_mx0w1,
      or_dcpl_344);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_9_0_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_14_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_103_mx0w1,
      or_dcpl_344);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_22_13_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_15_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_107_mx0w1,
      or_dcpl_354);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_9_0_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_15_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_106_mx0w1,
      or_dcpl_354);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_22_13_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_110_mx0w1,
      or_dcpl_364);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_9_0_mx1 = MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_lpi_1_dfm,
      FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_109_mx0w1,
      or_dcpl_364);
  assign IsNaN_8U_23U_land_1_lpi_1_dfm_mx0w0 = ~((~((chn_mul_in_rsci_d_mxwt[22:0]!=23'b00000000000000000000000)))
      | (chn_mul_in_rsci_d_mxwt[30:23]!=8'b11111111));
  assign IsNaN_8U_23U_land_2_lpi_1_dfm_mx0w0 = ~((~((chn_mul_in_rsci_d_mxwt[55:33]!=23'b00000000000000000000000)))
      | (chn_mul_in_rsci_d_mxwt[63:56]!=8'b11111111));
  assign IsNaN_8U_23U_land_3_lpi_1_dfm_mx0w0 = ~((~((chn_mul_in_rsci_d_mxwt[88:66]!=23'b00000000000000000000000)))
      | (chn_mul_in_rsci_d_mxwt[96:89]!=8'b11111111));
  assign IsNaN_8U_23U_land_4_lpi_1_dfm_mx0w0 = ~((~((chn_mul_in_rsci_d_mxwt[121:99]!=23'b00000000000000000000000)))
      | (chn_mul_in_rsci_d_mxwt[129:122]!=8'b11111111));
  assign IsNaN_8U_23U_land_5_lpi_1_dfm_mx0w0 = ~((~((chn_mul_in_rsci_d_mxwt[154:132]!=23'b00000000000000000000000)))
      | (chn_mul_in_rsci_d_mxwt[162:155]!=8'b11111111));
  assign IsNaN_8U_23U_land_6_lpi_1_dfm_mx0w0 = ~((~((chn_mul_in_rsci_d_mxwt[187:165]!=23'b00000000000000000000000)))
      | (chn_mul_in_rsci_d_mxwt[195:188]!=8'b11111111));
  assign IsNaN_8U_23U_land_7_lpi_1_dfm_mx0w0 = ~((~((chn_mul_in_rsci_d_mxwt[220:198]!=23'b00000000000000000000000)))
      | (chn_mul_in_rsci_d_mxwt[228:221]!=8'b11111111));
  assign IsNaN_8U_23U_land_8_lpi_1_dfm_mx0w0 = ~((~((chn_mul_in_rsci_d_mxwt[253:231]!=23'b00000000000000000000000)))
      | (chn_mul_in_rsci_d_mxwt[261:254]!=8'b11111111));
  assign IsNaN_8U_23U_land_9_lpi_1_dfm_mx0w0 = ~((~((chn_mul_in_rsci_d_mxwt[286:264]!=23'b00000000000000000000000)))
      | (chn_mul_in_rsci_d_mxwt[294:287]!=8'b11111111));
  assign IsNaN_8U_23U_land_10_lpi_1_dfm_mx0w0 = ~((~((chn_mul_in_rsci_d_mxwt[319:297]!=23'b00000000000000000000000)))
      | (chn_mul_in_rsci_d_mxwt[327:320]!=8'b11111111));
  assign IsNaN_8U_23U_land_11_lpi_1_dfm_mx0w0 = ~((~((chn_mul_in_rsci_d_mxwt[352:330]!=23'b00000000000000000000000)))
      | (chn_mul_in_rsci_d_mxwt[360:353]!=8'b11111111));
  assign IsNaN_8U_23U_land_12_lpi_1_dfm_mx0w0 = ~((~((chn_mul_in_rsci_d_mxwt[385:363]!=23'b00000000000000000000000)))
      | (chn_mul_in_rsci_d_mxwt[393:386]!=8'b11111111));
  assign IsNaN_8U_23U_land_13_lpi_1_dfm_mx0w0 = ~((~((chn_mul_in_rsci_d_mxwt[418:396]!=23'b00000000000000000000000)))
      | (chn_mul_in_rsci_d_mxwt[426:419]!=8'b11111111));
  assign IsNaN_8U_23U_land_14_lpi_1_dfm_mx0w0 = ~((~((chn_mul_in_rsci_d_mxwt[451:429]!=23'b00000000000000000000000)))
      | (chn_mul_in_rsci_d_mxwt[459:452]!=8'b11111111));
  assign IsNaN_8U_23U_land_15_lpi_1_dfm_mx0w0 = ~((~((chn_mul_in_rsci_d_mxwt[484:462]!=23'b00000000000000000000000)))
      | (chn_mul_in_rsci_d_mxwt[492:485]!=8'b11111111));
  assign IsNaN_8U_23U_land_lpi_1_dfm_mx0w0 = ~((~((chn_mul_in_rsci_d_mxwt[517:495]!=23'b00000000000000000000000)))
      | (chn_mul_in_rsci_d_mxwt[525:518]!=8'b11111111));
  assign IsDenorm_5U_23U_land_1_lpi_1_dfm = ((mul_nan_to_zero_op_mant_1_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_1_sva;
  assign mul_nan_to_zero_aelse_not_110_nl = ~ mul_nan_to_zero_land_1_lpi_1_dfm;
  assign mul_nan_to_zero_op_mant_1_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_MulOp_data_0_9_0_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_110_nl));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_1_sva = ~((mul_nan_to_zero_op_expo_1_lpi_1_dfm!=5'b00000));
  assign mul_nan_to_zero_aelse_not_48_nl = ~ mul_nan_to_zero_land_1_lpi_1_dfm;
  assign mul_nan_to_zero_op_expo_1_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_MulOp_data_0_14_10_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_48_nl));
  assign else_MulOp_data_0_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_mul_op_1_sva_1[9:0]),
      (chn_mul_op_rsci_d_mxwt[9:0]), cfg_mul_src_1_sva_1);
  assign IsNaN_5U_10U_nor_tmp = ~((else_MulOp_data_0_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign mul_nan_to_zero_land_1_lpi_1_dfm = (~(IsNaN_5U_10U_nor_tmp | (else_MulOp_data_0_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_MulOp_data_0_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]),
      (chn_mul_op_rsci_d_mxwt[14:10]), cfg_mul_src_1_sva_1);
  assign IsDenorm_5U_23U_land_2_lpi_1_dfm = ((mul_nan_to_zero_op_mant_2_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_2_sva;
  assign mul_nan_to_zero_aelse_not_108_nl = ~ mul_nan_to_zero_land_2_lpi_1_dfm;
  assign mul_nan_to_zero_op_mant_2_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_MulOp_data_1_9_0_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_108_nl));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_2_sva = ~((mul_nan_to_zero_op_expo_2_lpi_1_dfm!=5'b00000));
  assign mul_nan_to_zero_aelse_not_50_nl = ~ mul_nan_to_zero_land_2_lpi_1_dfm;
  assign mul_nan_to_zero_op_expo_2_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_MulOp_data_1_14_10_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_50_nl));
  assign else_MulOp_data_1_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_mul_op_1_sva_1[9:0]),
      (chn_mul_op_rsci_d_mxwt[25:16]), cfg_mul_src_1_sva_1);
  assign IsNaN_5U_10U_nor_1_tmp = ~((else_MulOp_data_1_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign mul_nan_to_zero_land_2_lpi_1_dfm = (~(IsNaN_5U_10U_nor_1_tmp | (else_MulOp_data_1_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_MulOp_data_1_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]),
      (chn_mul_op_rsci_d_mxwt[30:26]), cfg_mul_src_1_sva_1);
  assign IsDenorm_5U_23U_land_3_lpi_1_dfm = ((mul_nan_to_zero_op_mant_3_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_3_sva;
  assign mul_nan_to_zero_aelse_not_106_nl = ~ mul_nan_to_zero_land_3_lpi_1_dfm;
  assign mul_nan_to_zero_op_mant_3_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_MulOp_data_2_9_0_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_106_nl));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_3_sva = ~((mul_nan_to_zero_op_expo_3_lpi_1_dfm!=5'b00000));
  assign mul_nan_to_zero_aelse_not_52_nl = ~ mul_nan_to_zero_land_3_lpi_1_dfm;
  assign mul_nan_to_zero_op_expo_3_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_MulOp_data_2_14_10_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_52_nl));
  assign else_MulOp_data_2_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_mul_op_1_sva_1[9:0]),
      (chn_mul_op_rsci_d_mxwt[41:32]), cfg_mul_src_1_sva_1);
  assign IsNaN_5U_10U_nor_2_tmp = ~((else_MulOp_data_2_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign mul_nan_to_zero_land_3_lpi_1_dfm = (~(IsNaN_5U_10U_nor_2_tmp | (else_MulOp_data_2_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_MulOp_data_2_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]),
      (chn_mul_op_rsci_d_mxwt[46:42]), cfg_mul_src_1_sva_1);
  assign IsDenorm_5U_23U_land_4_lpi_1_dfm = ((mul_nan_to_zero_op_mant_4_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_4_sva;
  assign mul_nan_to_zero_aelse_not_104_nl = ~ mul_nan_to_zero_land_4_lpi_1_dfm;
  assign mul_nan_to_zero_op_mant_4_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_MulOp_data_3_9_0_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_104_nl));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_4_sva = ~((mul_nan_to_zero_op_expo_4_lpi_1_dfm!=5'b00000));
  assign mul_nan_to_zero_aelse_not_54_nl = ~ mul_nan_to_zero_land_4_lpi_1_dfm;
  assign mul_nan_to_zero_op_expo_4_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_MulOp_data_3_14_10_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_54_nl));
  assign else_MulOp_data_3_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_mul_op_1_sva_1[9:0]),
      (chn_mul_op_rsci_d_mxwt[57:48]), cfg_mul_src_1_sva_1);
  assign IsNaN_5U_10U_nor_3_tmp = ~((else_MulOp_data_3_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign mul_nan_to_zero_land_4_lpi_1_dfm = (~(IsNaN_5U_10U_nor_3_tmp | (else_MulOp_data_3_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_MulOp_data_3_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]),
      (chn_mul_op_rsci_d_mxwt[62:58]), cfg_mul_src_1_sva_1);
  assign IsDenorm_5U_23U_land_5_lpi_1_dfm = ((mul_nan_to_zero_op_mant_5_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_5_sva;
  assign mul_nan_to_zero_aelse_not_102_nl = ~ mul_nan_to_zero_land_5_lpi_1_dfm;
  assign mul_nan_to_zero_op_mant_5_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_MulOp_data_4_9_0_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_102_nl));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_5_sva = ~((mul_nan_to_zero_op_expo_5_lpi_1_dfm!=5'b00000));
  assign mul_nan_to_zero_aelse_not_56_nl = ~ mul_nan_to_zero_land_5_lpi_1_dfm;
  assign mul_nan_to_zero_op_expo_5_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_MulOp_data_4_14_10_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_56_nl));
  assign else_MulOp_data_4_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_mul_op_1_sva_1[9:0]),
      (chn_mul_op_rsci_d_mxwt[73:64]), cfg_mul_src_1_sva_1);
  assign IsNaN_5U_10U_nor_4_tmp = ~((else_MulOp_data_4_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign mul_nan_to_zero_land_5_lpi_1_dfm = (~(IsNaN_5U_10U_nor_4_tmp | (else_MulOp_data_4_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_MulOp_data_4_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]),
      (chn_mul_op_rsci_d_mxwt[78:74]), cfg_mul_src_1_sva_1);
  assign IsDenorm_5U_23U_land_6_lpi_1_dfm = ((mul_nan_to_zero_op_mant_6_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_6_sva;
  assign mul_nan_to_zero_aelse_not_100_nl = ~ mul_nan_to_zero_land_6_lpi_1_dfm;
  assign mul_nan_to_zero_op_mant_6_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_MulOp_data_5_9_0_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_100_nl));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_6_sva = ~((mul_nan_to_zero_op_expo_6_lpi_1_dfm!=5'b00000));
  assign mul_nan_to_zero_aelse_not_58_nl = ~ mul_nan_to_zero_land_6_lpi_1_dfm;
  assign mul_nan_to_zero_op_expo_6_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_MulOp_data_5_14_10_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_58_nl));
  assign else_MulOp_data_5_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_mul_op_1_sva_1[9:0]),
      (chn_mul_op_rsci_d_mxwt[89:80]), cfg_mul_src_1_sva_1);
  assign IsNaN_5U_10U_nor_5_tmp = ~((else_MulOp_data_5_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign mul_nan_to_zero_land_6_lpi_1_dfm = (~(IsNaN_5U_10U_nor_5_tmp | (else_MulOp_data_5_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_MulOp_data_5_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]),
      (chn_mul_op_rsci_d_mxwt[94:90]), cfg_mul_src_1_sva_1);
  assign IsDenorm_5U_23U_land_7_lpi_1_dfm = ((mul_nan_to_zero_op_mant_7_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_7_sva;
  assign mul_nan_to_zero_aelse_not_98_nl = ~ mul_nan_to_zero_land_7_lpi_1_dfm;
  assign mul_nan_to_zero_op_mant_7_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_MulOp_data_6_9_0_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_98_nl));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_7_sva = ~((mul_nan_to_zero_op_expo_7_lpi_1_dfm!=5'b00000));
  assign mul_nan_to_zero_aelse_not_60_nl = ~ mul_nan_to_zero_land_7_lpi_1_dfm;
  assign mul_nan_to_zero_op_expo_7_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_MulOp_data_6_14_10_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_60_nl));
  assign else_MulOp_data_6_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_mul_op_1_sva_1[9:0]),
      (chn_mul_op_rsci_d_mxwt[105:96]), cfg_mul_src_1_sva_1);
  assign IsNaN_5U_10U_nor_6_tmp = ~((else_MulOp_data_6_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign mul_nan_to_zero_land_7_lpi_1_dfm = (~(IsNaN_5U_10U_nor_6_tmp | (else_MulOp_data_6_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_MulOp_data_6_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]),
      (chn_mul_op_rsci_d_mxwt[110:106]), cfg_mul_src_1_sva_1);
  assign IsDenorm_5U_23U_land_8_lpi_1_dfm = ((mul_nan_to_zero_op_mant_8_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_8_sva;
  assign mul_nan_to_zero_aelse_not_96_nl = ~ mul_nan_to_zero_land_8_lpi_1_dfm;
  assign mul_nan_to_zero_op_mant_8_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_MulOp_data_7_9_0_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_96_nl));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_8_sva = ~((mul_nan_to_zero_op_expo_8_lpi_1_dfm!=5'b00000));
  assign mul_nan_to_zero_aelse_not_62_nl = ~ mul_nan_to_zero_land_8_lpi_1_dfm;
  assign mul_nan_to_zero_op_expo_8_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_MulOp_data_7_14_10_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_62_nl));
  assign else_MulOp_data_7_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_mul_op_1_sva_1[9:0]),
      (chn_mul_op_rsci_d_mxwt[121:112]), cfg_mul_src_1_sva_1);
  assign IsNaN_5U_10U_nor_7_tmp = ~((else_MulOp_data_7_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign mul_nan_to_zero_land_8_lpi_1_dfm = (~(IsNaN_5U_10U_nor_7_tmp | (else_MulOp_data_7_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_MulOp_data_7_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]),
      (chn_mul_op_rsci_d_mxwt[126:122]), cfg_mul_src_1_sva_1);
  assign IsDenorm_5U_23U_land_9_lpi_1_dfm = ((mul_nan_to_zero_op_mant_9_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_9_sva;
  assign mul_nan_to_zero_aelse_not_94_nl = ~ mul_nan_to_zero_land_9_lpi_1_dfm;
  assign mul_nan_to_zero_op_mant_9_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_MulOp_data_8_9_0_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_94_nl));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_9_sva = ~((mul_nan_to_zero_op_expo_9_lpi_1_dfm!=5'b00000));
  assign mul_nan_to_zero_aelse_not_64_nl = ~ mul_nan_to_zero_land_9_lpi_1_dfm;
  assign mul_nan_to_zero_op_expo_9_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_MulOp_data_8_14_10_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_64_nl));
  assign else_MulOp_data_8_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_mul_op_1_sva_1[9:0]),
      (chn_mul_op_rsci_d_mxwt[137:128]), cfg_mul_src_1_sva_1);
  assign IsNaN_5U_10U_nor_8_tmp = ~((else_MulOp_data_8_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign mul_nan_to_zero_land_9_lpi_1_dfm = (~(IsNaN_5U_10U_nor_8_tmp | (else_MulOp_data_8_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_MulOp_data_8_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]),
      (chn_mul_op_rsci_d_mxwt[142:138]), cfg_mul_src_1_sva_1);
  assign IsDenorm_5U_23U_land_10_lpi_1_dfm = ((mul_nan_to_zero_op_mant_10_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_10_sva;
  assign mul_nan_to_zero_aelse_not_92_nl = ~ mul_nan_to_zero_land_10_lpi_1_dfm;
  assign mul_nan_to_zero_op_mant_10_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_MulOp_data_9_9_0_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_92_nl));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_10_sva = ~((mul_nan_to_zero_op_expo_10_lpi_1_dfm!=5'b00000));
  assign mul_nan_to_zero_aelse_not_66_nl = ~ mul_nan_to_zero_land_10_lpi_1_dfm;
  assign mul_nan_to_zero_op_expo_10_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_MulOp_data_9_14_10_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_66_nl));
  assign else_MulOp_data_9_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_mul_op_1_sva_1[9:0]),
      (chn_mul_op_rsci_d_mxwt[153:144]), cfg_mul_src_1_sva_1);
  assign IsNaN_5U_10U_nor_9_tmp = ~((else_MulOp_data_9_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign mul_nan_to_zero_land_10_lpi_1_dfm = (~(IsNaN_5U_10U_nor_9_tmp | (else_MulOp_data_9_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_MulOp_data_9_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]),
      (chn_mul_op_rsci_d_mxwt[158:154]), cfg_mul_src_1_sva_1);
  assign IsDenorm_5U_23U_land_11_lpi_1_dfm = ((mul_nan_to_zero_op_mant_11_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_11_sva;
  assign mul_nan_to_zero_aelse_not_90_nl = ~ mul_nan_to_zero_land_11_lpi_1_dfm;
  assign mul_nan_to_zero_op_mant_11_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_MulOp_data_10_9_0_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_90_nl));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_11_sva = ~((mul_nan_to_zero_op_expo_11_lpi_1_dfm!=5'b00000));
  assign mul_nan_to_zero_aelse_not_68_nl = ~ mul_nan_to_zero_land_11_lpi_1_dfm;
  assign mul_nan_to_zero_op_expo_11_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_MulOp_data_10_14_10_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_68_nl));
  assign else_MulOp_data_10_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_mul_op_1_sva_1[9:0]),
      (chn_mul_op_rsci_d_mxwt[169:160]), cfg_mul_src_1_sva_1);
  assign IsNaN_5U_10U_nor_10_tmp = ~((else_MulOp_data_10_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign mul_nan_to_zero_land_11_lpi_1_dfm = (~(IsNaN_5U_10U_nor_10_tmp | (else_MulOp_data_10_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_MulOp_data_10_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]),
      (chn_mul_op_rsci_d_mxwt[174:170]), cfg_mul_src_1_sva_1);
  assign IsDenorm_5U_23U_land_12_lpi_1_dfm = ((mul_nan_to_zero_op_mant_12_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_12_sva;
  assign mul_nan_to_zero_aelse_not_88_nl = ~ mul_nan_to_zero_land_12_lpi_1_dfm;
  assign mul_nan_to_zero_op_mant_12_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_MulOp_data_11_9_0_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_88_nl));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_12_sva = ~((mul_nan_to_zero_op_expo_12_lpi_1_dfm!=5'b00000));
  assign mul_nan_to_zero_aelse_not_70_nl = ~ mul_nan_to_zero_land_12_lpi_1_dfm;
  assign mul_nan_to_zero_op_expo_12_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_MulOp_data_11_14_10_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_70_nl));
  assign else_MulOp_data_11_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_mul_op_1_sva_1[9:0]),
      (chn_mul_op_rsci_d_mxwt[185:176]), cfg_mul_src_1_sva_1);
  assign IsNaN_5U_10U_nor_11_tmp = ~((else_MulOp_data_11_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign mul_nan_to_zero_land_12_lpi_1_dfm = (~(IsNaN_5U_10U_nor_11_tmp | (else_MulOp_data_11_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_MulOp_data_11_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]),
      (chn_mul_op_rsci_d_mxwt[190:186]), cfg_mul_src_1_sva_1);
  assign IsDenorm_5U_23U_land_13_lpi_1_dfm = ((mul_nan_to_zero_op_mant_13_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_13_sva;
  assign mul_nan_to_zero_aelse_not_86_nl = ~ mul_nan_to_zero_land_13_lpi_1_dfm;
  assign mul_nan_to_zero_op_mant_13_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_MulOp_data_12_9_0_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_86_nl));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_13_sva = ~((mul_nan_to_zero_op_expo_13_lpi_1_dfm!=5'b00000));
  assign mul_nan_to_zero_aelse_not_72_nl = ~ mul_nan_to_zero_land_13_lpi_1_dfm;
  assign mul_nan_to_zero_op_expo_13_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_MulOp_data_12_14_10_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_72_nl));
  assign else_MulOp_data_12_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_mul_op_1_sva_1[9:0]),
      (chn_mul_op_rsci_d_mxwt[201:192]), cfg_mul_src_1_sva_1);
  assign IsNaN_5U_10U_nor_12_tmp = ~((else_MulOp_data_12_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign mul_nan_to_zero_land_13_lpi_1_dfm = (~(IsNaN_5U_10U_nor_12_tmp | (else_MulOp_data_12_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_MulOp_data_12_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]),
      (chn_mul_op_rsci_d_mxwt[206:202]), cfg_mul_src_1_sva_1);
  assign IsDenorm_5U_23U_land_14_lpi_1_dfm = ((mul_nan_to_zero_op_mant_14_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_14_sva;
  assign mul_nan_to_zero_aelse_not_84_nl = ~ mul_nan_to_zero_land_14_lpi_1_dfm;
  assign mul_nan_to_zero_op_mant_14_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_MulOp_data_13_9_0_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_84_nl));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_14_sva = ~((mul_nan_to_zero_op_expo_14_lpi_1_dfm!=5'b00000));
  assign mul_nan_to_zero_aelse_not_74_nl = ~ mul_nan_to_zero_land_14_lpi_1_dfm;
  assign mul_nan_to_zero_op_expo_14_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_MulOp_data_13_14_10_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_74_nl));
  assign else_MulOp_data_13_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_mul_op_1_sva_1[9:0]),
      (chn_mul_op_rsci_d_mxwt[217:208]), cfg_mul_src_1_sva_1);
  assign IsNaN_5U_10U_nor_13_tmp = ~((else_MulOp_data_13_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign mul_nan_to_zero_land_14_lpi_1_dfm = (~(IsNaN_5U_10U_nor_13_tmp | (else_MulOp_data_13_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_MulOp_data_13_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]),
      (chn_mul_op_rsci_d_mxwt[222:218]), cfg_mul_src_1_sva_1);
  assign IsDenorm_5U_23U_land_15_lpi_1_dfm = ((mul_nan_to_zero_op_mant_15_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_15_sva;
  assign mul_nan_to_zero_aelse_not_82_nl = ~ mul_nan_to_zero_land_15_lpi_1_dfm;
  assign mul_nan_to_zero_op_mant_15_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_MulOp_data_14_9_0_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_82_nl));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_15_sva = ~((mul_nan_to_zero_op_expo_15_lpi_1_dfm!=5'b00000));
  assign mul_nan_to_zero_aelse_not_76_nl = ~ mul_nan_to_zero_land_15_lpi_1_dfm;
  assign mul_nan_to_zero_op_expo_15_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_MulOp_data_14_14_10_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_76_nl));
  assign else_MulOp_data_14_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_mul_op_1_sva_1[9:0]),
      (chn_mul_op_rsci_d_mxwt[233:224]), cfg_mul_src_1_sva_1);
  assign IsNaN_5U_10U_nor_14_tmp = ~((else_MulOp_data_14_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign mul_nan_to_zero_land_15_lpi_1_dfm = (~(IsNaN_5U_10U_nor_14_tmp | (else_MulOp_data_14_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_MulOp_data_14_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]),
      (chn_mul_op_rsci_d_mxwt[238:234]), cfg_mul_src_1_sva_1);
  assign IsDenorm_5U_23U_land_lpi_1_dfm = ((mul_nan_to_zero_op_mant_lpi_1_dfm!=10'b0000000000))
      & IsZero_5U_23U_IsZero_5U_23U_nor_cse_sva;
  assign mul_nan_to_zero_aelse_not_80_nl = ~ mul_nan_to_zero_land_lpi_1_dfm;
  assign mul_nan_to_zero_op_mant_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000, else_MulOp_data_15_9_0_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_80_nl));
  assign IsZero_5U_23U_IsZero_5U_23U_nor_cse_sva = ~((mul_nan_to_zero_op_expo_lpi_1_dfm!=5'b00000));
  assign mul_nan_to_zero_aelse_not_78_nl = ~ mul_nan_to_zero_land_lpi_1_dfm;
  assign mul_nan_to_zero_op_expo_lpi_1_dfm = MUX_v_5_2_2(5'b00000, else_MulOp_data_15_14_10_lpi_1_dfm_mx0,
      (mul_nan_to_zero_aelse_not_78_nl));
  assign else_MulOp_data_15_9_0_lpi_1_dfm_mx0 = MUX_v_10_2_2((cfg_mul_op_1_sva_1[9:0]),
      (chn_mul_op_rsci_d_mxwt[249:240]), cfg_mul_src_1_sva_1);
  assign IsNaN_5U_10U_nor_15_tmp = ~((else_MulOp_data_15_9_0_lpi_1_dfm_mx0!=10'b0000000000));
  assign mul_nan_to_zero_land_lpi_1_dfm = (~(IsNaN_5U_10U_nor_15_tmp | (else_MulOp_data_15_14_10_lpi_1_dfm_mx0!=5'b11111)))
      & cfg_nan_to_zero;
  assign else_MulOp_data_15_14_10_lpi_1_dfm_mx0 = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]),
      (chn_mul_op_rsci_d_mxwt[254:250]), cfg_mul_src_1_sva_1);
  assign nl_FpMul_8U_23U_oelse_1_acc_nl = conv_u2s_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_9})
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_nl = nl_FpMul_8U_23U_oelse_1_acc_nl[8:0];
  assign nl_mul_loop_mul_1_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_nl)
      + conv_u2s_8_10(MulIn_data_sva_534[30:23]);
  assign mul_loop_mul_1_FpMul_8U_23U_oelse_1_acc_nl = nl_mul_loop_mul_1_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign mul_loop_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((mul_loop_mul_1_FpMul_8U_23U_oelse_1_acc_nl));
  assign nl_FpMul_8U_23U_oelse_1_acc_1_nl = conv_u2s_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_9})
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_1_nl = nl_FpMul_8U_23U_oelse_1_acc_1_nl[8:0];
  assign nl_mul_loop_mul_2_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_1_nl)
      + conv_u2s_8_10(MulIn_data_sva_534[63:56]);
  assign mul_loop_mul_2_FpMul_8U_23U_oelse_1_acc_nl = nl_mul_loop_mul_2_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign mul_loop_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((mul_loop_mul_2_FpMul_8U_23U_oelse_1_acc_nl));
  assign nl_FpMul_8U_23U_oelse_1_acc_2_nl = conv_u2s_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_9})
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_2_nl = nl_FpMul_8U_23U_oelse_1_acc_2_nl[8:0];
  assign nl_mul_loop_mul_3_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_2_nl)
      + conv_u2s_8_10(MulIn_data_sva_534[96:89]);
  assign mul_loop_mul_3_FpMul_8U_23U_oelse_1_acc_nl = nl_mul_loop_mul_3_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign mul_loop_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((mul_loop_mul_3_FpMul_8U_23U_oelse_1_acc_nl));
  assign nl_FpMul_8U_23U_oelse_1_acc_3_nl = conv_u2s_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_9})
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_3_nl = nl_FpMul_8U_23U_oelse_1_acc_3_nl[8:0];
  assign nl_mul_loop_mul_4_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_3_nl)
      + conv_u2s_8_10(MulIn_data_sva_534[129:122]);
  assign mul_loop_mul_4_FpMul_8U_23U_oelse_1_acc_nl = nl_mul_loop_mul_4_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign mul_loop_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((mul_loop_mul_4_FpMul_8U_23U_oelse_1_acc_nl));
  assign nl_FpMul_8U_23U_oelse_1_acc_4_nl = conv_u2s_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_9})
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_4_nl = nl_FpMul_8U_23U_oelse_1_acc_4_nl[8:0];
  assign nl_mul_loop_mul_5_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_4_nl)
      + conv_u2s_8_10(MulIn_data_sva_534[162:155]);
  assign mul_loop_mul_5_FpMul_8U_23U_oelse_1_acc_nl = nl_mul_loop_mul_5_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign mul_loop_mul_5_FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((mul_loop_mul_5_FpMul_8U_23U_oelse_1_acc_nl));
  assign nl_FpMul_8U_23U_oelse_1_acc_5_nl = conv_u2s_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_9})
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_5_nl = nl_FpMul_8U_23U_oelse_1_acc_5_nl[8:0];
  assign nl_mul_loop_mul_6_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_5_nl)
      + conv_u2s_8_10(MulIn_data_sva_534[195:188]);
  assign mul_loop_mul_6_FpMul_8U_23U_oelse_1_acc_nl = nl_mul_loop_mul_6_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign mul_loop_mul_6_FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((mul_loop_mul_6_FpMul_8U_23U_oelse_1_acc_nl));
  assign nl_FpMul_8U_23U_oelse_1_acc_6_nl = conv_u2s_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_9})
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_6_nl = nl_FpMul_8U_23U_oelse_1_acc_6_nl[8:0];
  assign nl_mul_loop_mul_7_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_6_nl)
      + conv_u2s_8_10(MulIn_data_sva_534[228:221]);
  assign mul_loop_mul_7_FpMul_8U_23U_oelse_1_acc_nl = nl_mul_loop_mul_7_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign mul_loop_mul_7_FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((mul_loop_mul_7_FpMul_8U_23U_oelse_1_acc_nl));
  assign nl_FpMul_8U_23U_oelse_1_acc_7_nl = conv_u2s_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_9})
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_7_nl = nl_FpMul_8U_23U_oelse_1_acc_7_nl[8:0];
  assign nl_mul_loop_mul_8_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_7_nl)
      + conv_u2s_8_10(MulIn_data_sva_534[261:254]);
  assign mul_loop_mul_8_FpMul_8U_23U_oelse_1_acc_nl = nl_mul_loop_mul_8_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign mul_loop_mul_8_FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((mul_loop_mul_8_FpMul_8U_23U_oelse_1_acc_nl));
  assign nl_FpMul_8U_23U_oelse_1_acc_8_nl = conv_u2s_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_9})
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_8_nl = nl_FpMul_8U_23U_oelse_1_acc_8_nl[8:0];
  assign nl_mul_loop_mul_9_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_8_nl)
      + conv_u2s_8_10(MulIn_data_sva_534[294:287]);
  assign mul_loop_mul_9_FpMul_8U_23U_oelse_1_acc_nl = nl_mul_loop_mul_9_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign mul_loop_mul_9_FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((mul_loop_mul_9_FpMul_8U_23U_oelse_1_acc_nl));
  assign nl_FpMul_8U_23U_oelse_1_acc_9_nl = conv_u2s_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_9})
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_9_nl = nl_FpMul_8U_23U_oelse_1_acc_9_nl[8:0];
  assign nl_mul_loop_mul_10_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_9_nl)
      + conv_u2s_8_10(MulIn_data_sva_534[327:320]);
  assign mul_loop_mul_10_FpMul_8U_23U_oelse_1_acc_nl = nl_mul_loop_mul_10_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign mul_loop_mul_10_FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((mul_loop_mul_10_FpMul_8U_23U_oelse_1_acc_nl));
  assign nl_FpMul_8U_23U_oelse_1_acc_10_nl = conv_u2s_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_9})
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_10_nl = nl_FpMul_8U_23U_oelse_1_acc_10_nl[8:0];
  assign nl_mul_loop_mul_11_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_10_nl)
      + conv_u2s_8_10(MulIn_data_sva_534[360:353]);
  assign mul_loop_mul_11_FpMul_8U_23U_oelse_1_acc_nl = nl_mul_loop_mul_11_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign mul_loop_mul_11_FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((mul_loop_mul_11_FpMul_8U_23U_oelse_1_acc_nl));
  assign nl_FpMul_8U_23U_oelse_1_acc_11_nl = conv_u2s_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_9})
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_11_nl = nl_FpMul_8U_23U_oelse_1_acc_11_nl[8:0];
  assign nl_mul_loop_mul_12_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_11_nl)
      + conv_u2s_8_10(MulIn_data_sva_534[393:386]);
  assign mul_loop_mul_12_FpMul_8U_23U_oelse_1_acc_nl = nl_mul_loop_mul_12_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign mul_loop_mul_12_FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((mul_loop_mul_12_FpMul_8U_23U_oelse_1_acc_nl));
  assign nl_FpMul_8U_23U_oelse_1_acc_12_nl = conv_u2s_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_9})
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_12_nl = nl_FpMul_8U_23U_oelse_1_acc_12_nl[8:0];
  assign nl_mul_loop_mul_13_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_12_nl)
      + conv_u2s_8_10(MulIn_data_sva_534[426:419]);
  assign mul_loop_mul_13_FpMul_8U_23U_oelse_1_acc_nl = nl_mul_loop_mul_13_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign mul_loop_mul_13_FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((mul_loop_mul_13_FpMul_8U_23U_oelse_1_acc_nl));
  assign nl_FpMul_8U_23U_oelse_1_acc_13_nl = conv_u2s_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_9})
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_13_nl = nl_FpMul_8U_23U_oelse_1_acc_13_nl[8:0];
  assign nl_mul_loop_mul_14_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_13_nl)
      + conv_u2s_8_10(MulIn_data_sva_534[459:452]);
  assign mul_loop_mul_14_FpMul_8U_23U_oelse_1_acc_nl = nl_mul_loop_mul_14_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign mul_loop_mul_14_FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((mul_loop_mul_14_FpMul_8U_23U_oelse_1_acc_nl));
  assign nl_FpMul_8U_23U_oelse_1_acc_14_nl = conv_u2s_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_9})
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_14_nl = nl_FpMul_8U_23U_oelse_1_acc_14_nl[8:0];
  assign nl_mul_loop_mul_15_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_14_nl)
      + conv_u2s_8_10(MulIn_data_sva_534[492:485]);
  assign mul_loop_mul_15_FpMul_8U_23U_oelse_1_acc_nl = nl_mul_loop_mul_15_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign mul_loop_mul_15_FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((mul_loop_mul_15_FpMul_8U_23U_oelse_1_acc_nl));
  assign nl_FpMul_8U_23U_oelse_1_acc_15_nl = conv_u2s_8_9({FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_7_3_2_1
      , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_7_1_0_1 , FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_9})
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_15_nl = nl_FpMul_8U_23U_oelse_1_acc_15_nl[8:0];
  assign nl_mul_loop_mul_16_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_15_nl)
      + conv_u2s_8_10(MulIn_data_sva_534[525:518]);
  assign mul_loop_mul_16_FpMul_8U_23U_oelse_1_acc_nl = nl_mul_loop_mul_16_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign mul_loop_mul_16_FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((mul_loop_mul_16_FpMul_8U_23U_oelse_1_acc_nl));
  assign else_unequal_tmp = ~((cfg_precision==2'b10));
  assign nl_mul_loop_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_nl = ({reg_FpMul_8U_23U_p_expo_1_itm
      , reg_FpMul_8U_23U_p_expo_1_2_itm}) + 8'b1;
  assign mul_loop_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_mul_loop_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign FpMul_8U_23U_p_expo_1_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((mul_loop_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_nl),
      ({reg_FpMul_8U_23U_p_expo_1_itm , reg_FpMul_8U_23U_p_expo_1_2_itm}), FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_63_nl
      = ~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_1_lpi_1_dfm = MUX_v_23_2_2(FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_1_sva,
      23'b11111111111111111111111, (FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_63_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1 = FpMul_8U_23U_p_expo_1_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1[7:0];
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_1_sva = mul_loop_mul_1_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_1_sva_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_1_sva = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_1_sva[22:0];
  assign FpMul_8U_23U_o_expo_3_0_1_lpi_1_dfm_mx1 = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_lpi_1_dfm_1[3:0]),
      or_tmp_898);
  assign FpMul_8U_23U_lor_33_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_7_4_1_lpi_1_dfm!=4'b0000)
      | (FpMul_8U_23U_o_expo_3_0_1_lpi_1_dfm_mx1!=4'b0000))) | FpMul_8U_23U_lor_18_lpi_1_dfm_7;
  assign FpMul_8U_23U_o_expo_7_4_1_lpi_1_dfm = MUX_v_4_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_lpi_1_dfm_1[7:4]),
      4'b1111, FpMul_8U_23U_is_inf_1_lpi_1_dfm_2);
  assign FpMul_8U_23U_is_inf_1_lpi_1_dfm_2 = ~(FpMul_8U_23U_FpMul_8U_23U_and_itm_2
      | FpMul_8U_23U_lor_18_lpi_1_dfm_7);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_nl = (~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp)
      & mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_1_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp
      & mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_lpi_1_dfm_1 = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_1_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1, {(~ mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs_2)
      , (FpMantWidthDec_8U_47U_23U_0U_0U_and_nl) , (FpMantWidthDec_8U_47U_23U_0U_0U_and_1_nl)});
  assign nl_mul_loop_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_nl = ({reg_FpMul_8U_23U_p_expo_2_itm
      , reg_FpMul_8U_23U_p_expo_2_2_itm}) + 8'b1;
  assign mul_loop_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_mul_loop_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign FpMul_8U_23U_p_expo_2_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((mul_loop_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_nl),
      ({reg_FpMul_8U_23U_p_expo_2_itm , reg_FpMul_8U_23U_p_expo_2_2_itm}), FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_62_nl
      = ~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_2_lpi_1_dfm = MUX_v_23_2_2(FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_2_sva,
      23'b11111111111111111111111, (FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_62_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_1 = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1 = FpMul_8U_23U_p_expo_2_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1[7:0];
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_2_sva = mul_loop_mul_2_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_2_sva_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_2_sva = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_2_sva[22:0];
  assign FpMul_8U_23U_o_expo_3_0_2_lpi_1_dfm_mx1 = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_lpi_1_dfm_1[3:0]),
      or_tmp_980);
  assign FpMul_8U_23U_lor_34_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_7_4_2_lpi_1_dfm!=4'b0000)
      | (FpMul_8U_23U_o_expo_3_0_2_lpi_1_dfm_mx1!=4'b0000))) | FpMul_8U_23U_lor_19_lpi_1_dfm_7;
  assign FpMul_8U_23U_o_expo_7_4_2_lpi_1_dfm = MUX_v_4_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_lpi_1_dfm_1[7:4]),
      4'b1111, FpMul_8U_23U_is_inf_2_lpi_1_dfm_2);
  assign FpMul_8U_23U_is_inf_2_lpi_1_dfm_2 = ~(FpMul_8U_23U_FpMul_8U_23U_and_64_itm_2
      | FpMul_8U_23U_lor_19_lpi_1_dfm_7);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_2_nl = (~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_1)
      & mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_3_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_1
      & mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_lpi_1_dfm_1 = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_2_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1, {(~ mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs_2)
      , (FpMantWidthDec_8U_47U_23U_0U_0U_and_2_nl) , (FpMantWidthDec_8U_47U_23U_0U_0U_and_3_nl)});
  assign nl_mul_loop_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_nl = ({reg_FpMul_8U_23U_p_expo_3_itm
      , reg_FpMul_8U_23U_p_expo_3_2_itm}) + 8'b1;
  assign mul_loop_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_mul_loop_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign FpMul_8U_23U_p_expo_3_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((mul_loop_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_nl),
      ({reg_FpMul_8U_23U_p_expo_3_itm , reg_FpMul_8U_23U_p_expo_3_2_itm}), FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_61_nl
      = ~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_3_lpi_1_dfm = MUX_v_23_2_2(FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_3_sva,
      23'b11111111111111111111111, (FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_61_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_2 = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1 = FpMul_8U_23U_p_expo_3_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1[7:0];
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_3_sva = mul_loop_mul_3_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_3_sva_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_3_sva = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_3_sva[22:0];
  assign FpMul_8U_23U_o_expo_3_0_3_lpi_1_dfm_mx1 = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_lpi_1_dfm_1[3:0]),
      or_tmp_1060);
  assign FpMul_8U_23U_lor_35_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_7_4_3_lpi_1_dfm!=4'b0000)
      | (FpMul_8U_23U_o_expo_3_0_3_lpi_1_dfm_mx1!=4'b0000))) | FpMul_8U_23U_lor_20_lpi_1_dfm_7;
  assign FpMul_8U_23U_o_expo_7_4_3_lpi_1_dfm = MUX_v_4_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_lpi_1_dfm_1[7:4]),
      4'b1111, FpMul_8U_23U_is_inf_3_lpi_1_dfm_2);
  assign FpMul_8U_23U_is_inf_3_lpi_1_dfm_2 = ~(FpMul_8U_23U_FpMul_8U_23U_and_65_itm_2
      | FpMul_8U_23U_lor_20_lpi_1_dfm_7);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_4_nl = (~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_2)
      & mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_5_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_2
      & mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_lpi_1_dfm_1 = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_3_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1, {(~ mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs_2)
      , (FpMantWidthDec_8U_47U_23U_0U_0U_and_4_nl) , (FpMantWidthDec_8U_47U_23U_0U_0U_and_5_nl)});
  assign nl_mul_loop_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_nl = ({reg_FpMul_8U_23U_p_expo_4_itm
      , reg_FpMul_8U_23U_p_expo_4_2_itm}) + 8'b1;
  assign mul_loop_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_mul_loop_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign FpMul_8U_23U_p_expo_4_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((mul_loop_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_nl),
      ({reg_FpMul_8U_23U_p_expo_4_itm , reg_FpMul_8U_23U_p_expo_4_2_itm}), FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_60_nl
      = ~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_3;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_4_lpi_1_dfm = MUX_v_23_2_2(FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_4_sva,
      23'b11111111111111111111111, (FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_60_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_3 = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_4_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_4_sva_1 = FpMul_8U_23U_p_expo_4_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_4_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_4_sva_1[7:0];
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_4_sva = mul_loop_mul_4_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_4_sva_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_4_sva = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_4_sva[22:0];
  assign FpMul_8U_23U_o_expo_3_0_4_lpi_1_dfm_mx1 = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_4_lpi_1_dfm_1[3:0]),
      or_tmp_1142);
  assign FpMul_8U_23U_lor_36_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_7_4_4_lpi_1_dfm!=4'b0000)
      | (FpMul_8U_23U_o_expo_3_0_4_lpi_1_dfm_mx1!=4'b0000))) | FpMul_8U_23U_lor_21_lpi_1_dfm_7;
  assign FpMul_8U_23U_o_expo_7_4_4_lpi_1_dfm = MUX_v_4_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_4_lpi_1_dfm_1[7:4]),
      4'b1111, FpMul_8U_23U_is_inf_4_lpi_1_dfm_2);
  assign FpMul_8U_23U_is_inf_4_lpi_1_dfm_2 = ~(FpMul_8U_23U_FpMul_8U_23U_and_66_itm_2
      | FpMul_8U_23U_lor_21_lpi_1_dfm_7);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_6_nl = (~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_3)
      & mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_7_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_3
      & mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_4_lpi_1_dfm_1 = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_4_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_4_sva_1, {(~ mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs_2)
      , (FpMantWidthDec_8U_47U_23U_0U_0U_and_6_nl) , (FpMantWidthDec_8U_47U_23U_0U_0U_and_7_nl)});
  assign nl_mul_loop_mul_5_FpMul_8U_23U_else_2_else_if_if_acc_nl = ({reg_FpMul_8U_23U_p_expo_5_itm
      , reg_FpMul_8U_23U_p_expo_5_2_itm}) + 8'b1;
  assign mul_loop_mul_5_FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_mul_loop_mul_5_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign FpMul_8U_23U_p_expo_5_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((mul_loop_mul_5_FpMul_8U_23U_else_2_else_if_if_acc_nl),
      ({reg_FpMul_8U_23U_p_expo_5_itm , reg_FpMul_8U_23U_p_expo_5_2_itm}), FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_4_itm_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_59_nl
      = ~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_4;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_5_lpi_1_dfm = MUX_v_23_2_2(FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_5_sva,
      23'b11111111111111111111111, (FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_59_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_4 = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_5_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_5_sva_1 = FpMul_8U_23U_p_expo_5_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_5_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_5_sva_1[7:0];
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_5_sva = mul_loop_mul_5_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_5_sva_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_5_sva = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_5_sva[22:0];
  assign FpMul_8U_23U_o_expo_3_0_5_lpi_1_dfm_mx1 = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_5_lpi_1_dfm_1[3:0]),
      or_tmp_1225);
  assign FpMul_8U_23U_lor_37_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_7_4_5_lpi_1_dfm!=4'b0000)
      | (FpMul_8U_23U_o_expo_3_0_5_lpi_1_dfm_mx1!=4'b0000))) | FpMul_8U_23U_lor_22_lpi_1_dfm_7;
  assign FpMul_8U_23U_o_expo_7_4_5_lpi_1_dfm = MUX_v_4_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_5_lpi_1_dfm_1[7:4]),
      4'b1111, FpMul_8U_23U_is_inf_5_lpi_1_dfm_2);
  assign FpMul_8U_23U_is_inf_5_lpi_1_dfm_2 = ~(FpMul_8U_23U_FpMul_8U_23U_and_67_itm_2
      | FpMul_8U_23U_lor_22_lpi_1_dfm_7);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_8_nl = (~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_4)
      & mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_9_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_4
      & mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_5_lpi_1_dfm_1 = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_5_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_5_sva_1, {(~ mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs_2)
      , (FpMantWidthDec_8U_47U_23U_0U_0U_and_8_nl) , (FpMantWidthDec_8U_47U_23U_0U_0U_and_9_nl)});
  assign nl_mul_loop_mul_6_FpMul_8U_23U_else_2_else_if_if_acc_nl = ({reg_FpMul_8U_23U_p_expo_6_itm
      , reg_FpMul_8U_23U_p_expo_6_2_itm}) + 8'b1;
  assign mul_loop_mul_6_FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_mul_loop_mul_6_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign FpMul_8U_23U_p_expo_6_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((mul_loop_mul_6_FpMul_8U_23U_else_2_else_if_if_acc_nl),
      ({reg_FpMul_8U_23U_p_expo_6_itm , reg_FpMul_8U_23U_p_expo_6_2_itm}), FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_5_itm_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_58_nl
      = ~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_5;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_6_lpi_1_dfm = MUX_v_23_2_2(FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_6_sva,
      23'b11111111111111111111111, (FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_58_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_5 = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_6_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_6_sva_1 = FpMul_8U_23U_p_expo_6_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_6_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_6_sva_1[7:0];
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_6_sva = mul_loop_mul_6_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_6_sva_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_6_sva = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_6_sva[22:0];
  assign FpMul_8U_23U_o_expo_3_0_6_lpi_1_dfm_mx1 = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_6_lpi_1_dfm_1[3:0]),
      or_tmp_1305);
  assign FpMul_8U_23U_lor_38_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_7_4_6_lpi_1_dfm!=4'b0000)
      | (FpMul_8U_23U_o_expo_3_0_6_lpi_1_dfm_mx1!=4'b0000))) | FpMul_8U_23U_lor_23_lpi_1_dfm_7;
  assign FpMul_8U_23U_o_expo_7_4_6_lpi_1_dfm = MUX_v_4_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_6_lpi_1_dfm_1[7:4]),
      4'b1111, FpMul_8U_23U_is_inf_6_lpi_1_dfm_2);
  assign FpMul_8U_23U_is_inf_6_lpi_1_dfm_2 = ~(FpMul_8U_23U_FpMul_8U_23U_and_68_itm_2
      | FpMul_8U_23U_lor_23_lpi_1_dfm_7);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_10_nl = (~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_5)
      & mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_11_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_5
      & mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_6_lpi_1_dfm_1 = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_6_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_6_sva_1, {(~ mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs_2)
      , (FpMantWidthDec_8U_47U_23U_0U_0U_and_10_nl) , (FpMantWidthDec_8U_47U_23U_0U_0U_and_11_nl)});
  assign nl_mul_loop_mul_7_FpMul_8U_23U_else_2_else_if_if_acc_nl = ({reg_FpMul_8U_23U_p_expo_7_itm
      , reg_FpMul_8U_23U_p_expo_7_2_itm}) + 8'b1;
  assign mul_loop_mul_7_FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_mul_loop_mul_7_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign FpMul_8U_23U_p_expo_7_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((mul_loop_mul_7_FpMul_8U_23U_else_2_else_if_if_acc_nl),
      ({reg_FpMul_8U_23U_p_expo_7_itm , reg_FpMul_8U_23U_p_expo_7_2_itm}), FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_6_itm_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_57_nl
      = ~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_6;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_7_lpi_1_dfm = MUX_v_23_2_2(FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_7_sva,
      23'b11111111111111111111111, (FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_57_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_6 = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_7_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_7_sva_1 = FpMul_8U_23U_p_expo_7_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_7_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_7_sva_1[7:0];
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_7_sva = mul_loop_mul_7_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_7_sva_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_7_sva = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_7_sva[22:0];
  assign FpMul_8U_23U_o_expo_3_0_7_lpi_1_dfm_mx1 = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_7_lpi_1_dfm_1[3:0]),
      or_tmp_1387);
  assign FpMul_8U_23U_lor_39_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_7_4_7_lpi_1_dfm!=4'b0000)
      | (FpMul_8U_23U_o_expo_3_0_7_lpi_1_dfm_mx1!=4'b0000))) | FpMul_8U_23U_lor_24_lpi_1_dfm_7;
  assign FpMul_8U_23U_o_expo_7_4_7_lpi_1_dfm = MUX_v_4_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_7_lpi_1_dfm_1[7:4]),
      4'b1111, FpMul_8U_23U_is_inf_7_lpi_1_dfm_2);
  assign FpMul_8U_23U_is_inf_7_lpi_1_dfm_2 = ~(FpMul_8U_23U_FpMul_8U_23U_and_69_itm_2
      | FpMul_8U_23U_lor_24_lpi_1_dfm_7);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_12_nl = (~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_6)
      & mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_13_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_6
      & mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_7_lpi_1_dfm_1 = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_7_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_7_sva_1, {(~ mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs_2)
      , (FpMantWidthDec_8U_47U_23U_0U_0U_and_12_nl) , (FpMantWidthDec_8U_47U_23U_0U_0U_and_13_nl)});
  assign nl_mul_loop_mul_8_FpMul_8U_23U_else_2_else_if_if_acc_nl = ({reg_FpMul_8U_23U_p_expo_8_itm
      , reg_FpMul_8U_23U_p_expo_8_2_itm}) + 8'b1;
  assign mul_loop_mul_8_FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_mul_loop_mul_8_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign FpMul_8U_23U_p_expo_8_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((mul_loop_mul_8_FpMul_8U_23U_else_2_else_if_if_acc_nl),
      ({reg_FpMul_8U_23U_p_expo_8_itm , reg_FpMul_8U_23U_p_expo_8_2_itm}), FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_7_itm_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_56_nl
      = ~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_7;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_8_lpi_1_dfm = MUX_v_23_2_2(FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_8_sva,
      23'b11111111111111111111111, (FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_56_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_7 = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_8_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_8_sva_1 = FpMul_8U_23U_p_expo_8_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_8_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_8_sva_1[7:0];
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_8_sva = mul_loop_mul_8_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_8_sva_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_8_sva = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_8_sva[22:0];
  assign FpMul_8U_23U_o_expo_3_0_8_lpi_1_dfm_mx1 = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_8_lpi_1_dfm_1[3:0]),
      or_tmp_1469);
  assign FpMul_8U_23U_lor_40_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_7_4_8_lpi_1_dfm!=4'b0000)
      | (FpMul_8U_23U_o_expo_3_0_8_lpi_1_dfm_mx1!=4'b0000))) | FpMul_8U_23U_lor_25_lpi_1_dfm_7;
  assign FpMul_8U_23U_o_expo_7_4_8_lpi_1_dfm = MUX_v_4_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_8_lpi_1_dfm_1[7:4]),
      4'b1111, FpMul_8U_23U_is_inf_8_lpi_1_dfm_2);
  assign FpMul_8U_23U_is_inf_8_lpi_1_dfm_2 = ~(FpMul_8U_23U_FpMul_8U_23U_and_70_itm_2
      | FpMul_8U_23U_lor_25_lpi_1_dfm_7);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_14_nl = (~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_7)
      & mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_15_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_7
      & mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_8_lpi_1_dfm_1 = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_8_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_8_sva_1, {(~ mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs_2)
      , (FpMantWidthDec_8U_47U_23U_0U_0U_and_14_nl) , (FpMantWidthDec_8U_47U_23U_0U_0U_and_15_nl)});
  assign nl_mul_loop_mul_9_FpMul_8U_23U_else_2_else_if_if_acc_nl = ({reg_FpMul_8U_23U_p_expo_9_itm
      , reg_FpMul_8U_23U_p_expo_9_2_itm}) + 8'b1;
  assign mul_loop_mul_9_FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_mul_loop_mul_9_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign FpMul_8U_23U_p_expo_9_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((mul_loop_mul_9_FpMul_8U_23U_else_2_else_if_if_acc_nl),
      ({reg_FpMul_8U_23U_p_expo_9_itm , reg_FpMul_8U_23U_p_expo_9_2_itm}), FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_8_itm_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_55_nl
      = ~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_8;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_9_lpi_1_dfm = MUX_v_23_2_2(FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_9_sva,
      23'b11111111111111111111111, (FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_55_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_8 = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_9_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_9_sva_1 = FpMul_8U_23U_p_expo_9_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_9_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_9_sva_1[7:0];
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_9_sva = mul_loop_mul_9_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_9_sva_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_9_sva = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_9_sva[22:0];
  assign FpMul_8U_23U_o_expo_3_0_9_lpi_1_dfm_mx1 = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_9_lpi_1_dfm_1[3:0]),
      or_tmp_1549);
  assign FpMul_8U_23U_lor_41_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_7_4_9_lpi_1_dfm!=4'b0000)
      | (FpMul_8U_23U_o_expo_3_0_9_lpi_1_dfm_mx1!=4'b0000))) | FpMul_8U_23U_lor_26_lpi_1_dfm_7;
  assign FpMul_8U_23U_o_expo_7_4_9_lpi_1_dfm = MUX_v_4_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_9_lpi_1_dfm_1[7:4]),
      4'b1111, FpMul_8U_23U_is_inf_9_lpi_1_dfm_2);
  assign FpMul_8U_23U_is_inf_9_lpi_1_dfm_2 = ~(FpMul_8U_23U_FpMul_8U_23U_and_71_itm_2
      | FpMul_8U_23U_lor_26_lpi_1_dfm_7);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_16_nl = (~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_8)
      & mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_17_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_8
      & mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_9_lpi_1_dfm_1 = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_9_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_9_sva_1, {(~ mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs_2)
      , (FpMantWidthDec_8U_47U_23U_0U_0U_and_16_nl) , (FpMantWidthDec_8U_47U_23U_0U_0U_and_17_nl)});
  assign nl_mul_loop_mul_10_FpMul_8U_23U_else_2_else_if_if_acc_nl = ({reg_FpMul_8U_23U_p_expo_10_itm
      , reg_FpMul_8U_23U_p_expo_10_2_itm}) + 8'b1;
  assign mul_loop_mul_10_FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_mul_loop_mul_10_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign FpMul_8U_23U_p_expo_10_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((mul_loop_mul_10_FpMul_8U_23U_else_2_else_if_if_acc_nl),
      ({reg_FpMul_8U_23U_p_expo_10_itm , reg_FpMul_8U_23U_p_expo_10_2_itm}), FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_9_itm_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_54_nl
      = ~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_9;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_10_lpi_1_dfm = MUX_v_23_2_2(FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_10_sva,
      23'b11111111111111111111111, (FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_54_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_9 = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_10_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_10_sva_1 = FpMul_8U_23U_p_expo_10_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_10_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_10_sva_1[7:0];
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_10_sva = mul_loop_mul_10_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_10_sva_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_10_sva = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_10_sva[22:0];
  assign FpMul_8U_23U_o_expo_3_0_10_lpi_1_dfm_mx1 = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_10_lpi_1_dfm_1[3:0]),
      or_tmp_1629);
  assign FpMul_8U_23U_lor_42_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_7_4_10_lpi_1_dfm!=4'b0000)
      | (FpMul_8U_23U_o_expo_3_0_10_lpi_1_dfm_mx1!=4'b0000))) | FpMul_8U_23U_lor_27_lpi_1_dfm_7;
  assign FpMul_8U_23U_o_expo_7_4_10_lpi_1_dfm = MUX_v_4_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_10_lpi_1_dfm_1[7:4]),
      4'b1111, FpMul_8U_23U_is_inf_10_lpi_1_dfm_2);
  assign FpMul_8U_23U_is_inf_10_lpi_1_dfm_2 = ~(FpMul_8U_23U_FpMul_8U_23U_and_72_itm_2
      | FpMul_8U_23U_lor_27_lpi_1_dfm_7);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_18_nl = (~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_9)
      & mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_19_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_9
      & mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_10_lpi_1_dfm_1 = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_10_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_10_sva_1, {(~ mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs_2)
      , (FpMantWidthDec_8U_47U_23U_0U_0U_and_18_nl) , (FpMantWidthDec_8U_47U_23U_0U_0U_and_19_nl)});
  assign nl_mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_nl = ({reg_FpMul_8U_23U_p_expo_11_itm
      , reg_FpMul_8U_23U_p_expo_11_2_itm}) + 8'b1;
  assign mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign FpMul_8U_23U_p_expo_11_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_nl),
      ({reg_FpMul_8U_23U_p_expo_11_itm , reg_FpMul_8U_23U_p_expo_11_2_itm}), FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_10_itm_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_53_nl
      = ~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_10;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_11_lpi_1_dfm = MUX_v_23_2_2(FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_11_sva,
      23'b11111111111111111111111, (FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_53_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_10 = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_11_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_11_sva_1 = FpMul_8U_23U_p_expo_11_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_11_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_11_sva_1[7:0];
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_11_sva = mul_loop_mul_11_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_11_sva_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_11_sva = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_11_sva[22:0];
  assign FpMul_8U_23U_o_expo_3_0_11_lpi_1_dfm_mx1 = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_11_lpi_1_dfm_1[3:0]),
      or_tmp_1709);
  assign FpMul_8U_23U_lor_43_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_7_4_11_lpi_1_dfm!=4'b0000)
      | (FpMul_8U_23U_o_expo_3_0_11_lpi_1_dfm_mx1!=4'b0000))) | FpMul_8U_23U_lor_28_lpi_1_dfm_7;
  assign FpMul_8U_23U_o_expo_7_4_11_lpi_1_dfm = MUX_v_4_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_11_lpi_1_dfm_1[7:4]),
      4'b1111, FpMul_8U_23U_is_inf_11_lpi_1_dfm_2);
  assign FpMul_8U_23U_is_inf_11_lpi_1_dfm_2 = ~(FpMul_8U_23U_FpMul_8U_23U_and_73_itm_2
      | FpMul_8U_23U_lor_28_lpi_1_dfm_7);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_20_nl = (~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_10)
      & mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_21_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_10
      & mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_11_lpi_1_dfm_1 = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_11_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_11_sva_1, {(~ mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs_2)
      , (FpMantWidthDec_8U_47U_23U_0U_0U_and_20_nl) , (FpMantWidthDec_8U_47U_23U_0U_0U_and_21_nl)});
  assign nl_mul_loop_mul_12_FpMul_8U_23U_else_2_else_if_if_acc_nl = ({reg_FpMul_8U_23U_p_expo_12_itm
      , reg_FpMul_8U_23U_p_expo_12_2_itm}) + 8'b1;
  assign mul_loop_mul_12_FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_mul_loop_mul_12_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign FpMul_8U_23U_p_expo_12_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((mul_loop_mul_12_FpMul_8U_23U_else_2_else_if_if_acc_nl),
      ({reg_FpMul_8U_23U_p_expo_12_itm , reg_FpMul_8U_23U_p_expo_12_2_itm}), FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_11_itm_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_52_nl
      = ~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_11;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_12_lpi_1_dfm = MUX_v_23_2_2(FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_12_sva,
      23'b11111111111111111111111, (FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_52_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_11 = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_12_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_12_sva_1 = FpMul_8U_23U_p_expo_12_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_12_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_12_sva_1[7:0];
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_12_sva = mul_loop_mul_12_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_12_sva_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_12_sva = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_12_sva[22:0];
  assign FpMul_8U_23U_o_expo_3_0_12_lpi_1_dfm_mx1 = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_12_lpi_1_dfm_1[3:0]),
      or_tmp_1786);
  assign FpMul_8U_23U_lor_44_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_7_4_12_lpi_1_dfm!=4'b0000)
      | (FpMul_8U_23U_o_expo_3_0_12_lpi_1_dfm_mx1!=4'b0000))) | FpMul_8U_23U_lor_29_lpi_1_dfm_7;
  assign FpMul_8U_23U_o_expo_7_4_12_lpi_1_dfm = MUX_v_4_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_12_lpi_1_dfm_1[7:4]),
      4'b1111, FpMul_8U_23U_is_inf_12_lpi_1_dfm_2);
  assign FpMul_8U_23U_is_inf_12_lpi_1_dfm_2 = ~(FpMul_8U_23U_FpMul_8U_23U_and_74_itm_2
      | FpMul_8U_23U_lor_29_lpi_1_dfm_7);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_22_nl = (~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_11)
      & mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_23_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_11
      & mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_12_lpi_1_dfm_1 = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_12_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_12_sva_1, {(~ mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs_2)
      , (FpMantWidthDec_8U_47U_23U_0U_0U_and_22_nl) , (FpMantWidthDec_8U_47U_23U_0U_0U_and_23_nl)});
  assign nl_mul_loop_mul_13_FpMul_8U_23U_else_2_else_if_if_acc_nl = ({reg_FpMul_8U_23U_p_expo_13_itm
      , reg_FpMul_8U_23U_p_expo_13_2_itm}) + 8'b1;
  assign mul_loop_mul_13_FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_mul_loop_mul_13_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign FpMul_8U_23U_p_expo_13_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((mul_loop_mul_13_FpMul_8U_23U_else_2_else_if_if_acc_nl),
      ({reg_FpMul_8U_23U_p_expo_13_itm , reg_FpMul_8U_23U_p_expo_13_2_itm}), FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_12_itm_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_51_nl
      = ~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_12;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_13_lpi_1_dfm = MUX_v_23_2_2(FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_13_sva,
      23'b11111111111111111111111, (FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_51_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_12 = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_13_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_13_sva_1 = FpMul_8U_23U_p_expo_13_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_13_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_13_sva_1[7:0];
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_13_sva = mul_loop_mul_13_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_13_sva_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_13_sva = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_13_sva[22:0];
  assign FpMul_8U_23U_o_expo_3_0_13_lpi_1_dfm_mx1 = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_13_lpi_1_dfm_1[3:0]),
      or_tmp_1869);
  assign FpMul_8U_23U_lor_45_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_7_4_13_lpi_1_dfm!=4'b0000)
      | (FpMul_8U_23U_o_expo_3_0_13_lpi_1_dfm_mx1!=4'b0000))) | FpMul_8U_23U_lor_30_lpi_1_dfm_7;
  assign FpMul_8U_23U_o_expo_7_4_13_lpi_1_dfm = MUX_v_4_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_13_lpi_1_dfm_1[7:4]),
      4'b1111, FpMul_8U_23U_is_inf_13_lpi_1_dfm_2);
  assign FpMul_8U_23U_is_inf_13_lpi_1_dfm_2 = ~(FpMul_8U_23U_FpMul_8U_23U_and_75_itm_2
      | FpMul_8U_23U_lor_30_lpi_1_dfm_7);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_24_nl = (~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_12)
      & mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_25_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_12
      & mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_13_lpi_1_dfm_1 = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_13_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_13_sva_1, {(~ mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs_2)
      , (FpMantWidthDec_8U_47U_23U_0U_0U_and_24_nl) , (FpMantWidthDec_8U_47U_23U_0U_0U_and_25_nl)});
  assign nl_mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_nl = ({reg_FpMul_8U_23U_p_expo_14_itm
      , reg_FpMul_8U_23U_p_expo_14_2_itm}) + 8'b1;
  assign mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign FpMul_8U_23U_p_expo_14_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_nl),
      ({reg_FpMul_8U_23U_p_expo_14_itm , reg_FpMul_8U_23U_p_expo_14_2_itm}), FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_13_itm_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_50_nl
      = ~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_13;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_14_lpi_1_dfm = MUX_v_23_2_2(FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_14_sva,
      23'b11111111111111111111111, (FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_50_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_13 = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_14_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_14_sva_1 = FpMul_8U_23U_p_expo_14_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_14_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_14_sva_1[7:0];
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_14_sva = mul_loop_mul_14_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_14_sva_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_14_sva = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_14_sva[22:0];
  assign FpMul_8U_23U_o_expo_3_0_14_lpi_1_dfm_mx1 = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_14_lpi_1_dfm_1[3:0]),
      or_tmp_1957);
  assign FpMul_8U_23U_lor_46_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_7_4_14_lpi_1_dfm!=4'b0000)
      | (FpMul_8U_23U_o_expo_3_0_14_lpi_1_dfm_mx1!=4'b0000))) | FpMul_8U_23U_lor_31_lpi_1_dfm_7;
  assign FpMul_8U_23U_o_expo_7_4_14_lpi_1_dfm = MUX_v_4_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_14_lpi_1_dfm_1[7:4]),
      4'b1111, FpMul_8U_23U_is_inf_14_lpi_1_dfm_2);
  assign FpMul_8U_23U_is_inf_14_lpi_1_dfm_2 = ~(FpMul_8U_23U_FpMul_8U_23U_and_76_itm_2
      | FpMul_8U_23U_lor_31_lpi_1_dfm_7);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_26_nl = (~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_13)
      & mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_27_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_13
      & mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_14_lpi_1_dfm_1 = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_14_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_14_sva_1, {(~ mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs_2)
      , (FpMantWidthDec_8U_47U_23U_0U_0U_and_26_nl) , (FpMantWidthDec_8U_47U_23U_0U_0U_and_27_nl)});
  assign nl_mul_loop_mul_15_FpMul_8U_23U_else_2_else_if_if_acc_nl = ({reg_FpMul_8U_23U_p_expo_15_itm
      , reg_FpMul_8U_23U_p_expo_15_2_itm}) + 8'b1;
  assign mul_loop_mul_15_FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_mul_loop_mul_15_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign FpMul_8U_23U_p_expo_15_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((mul_loop_mul_15_FpMul_8U_23U_else_2_else_if_if_acc_nl),
      ({reg_FpMul_8U_23U_p_expo_15_itm , reg_FpMul_8U_23U_p_expo_15_2_itm}), FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_14_itm_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_49_nl
      = ~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_14;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_15_lpi_1_dfm = MUX_v_23_2_2(FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_15_sva,
      23'b11111111111111111111111, (FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_49_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_14 = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_15_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_15_sva_1 = FpMul_8U_23U_p_expo_15_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_15_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_15_sva_1[7:0];
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_15_sva = mul_loop_mul_15_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_15_sva_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_15_sva = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_15_sva[22:0];
  assign FpMul_8U_23U_o_expo_3_0_15_lpi_1_dfm_mx1 = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_15_lpi_1_dfm_1[3:0]),
      or_tmp_2036);
  assign FpMul_8U_23U_lor_47_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_7_4_15_lpi_1_dfm!=4'b0000)
      | (FpMul_8U_23U_o_expo_3_0_15_lpi_1_dfm_mx1!=4'b0000))) | FpMul_8U_23U_lor_32_lpi_1_dfm_7;
  assign FpMul_8U_23U_o_expo_7_4_15_lpi_1_dfm = MUX_v_4_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_15_lpi_1_dfm_1[7:4]),
      4'b1111, FpMul_8U_23U_is_inf_15_lpi_1_dfm_2);
  assign FpMul_8U_23U_is_inf_15_lpi_1_dfm_2 = ~(FpMul_8U_23U_FpMul_8U_23U_and_77_itm_2
      | FpMul_8U_23U_lor_32_lpi_1_dfm_7);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_28_nl = (~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_14)
      & mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_29_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_14
      & mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_15_lpi_1_dfm_1 = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_15_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_15_sva_1, {(~ mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs_2)
      , (FpMantWidthDec_8U_47U_23U_0U_0U_and_28_nl) , (FpMantWidthDec_8U_47U_23U_0U_0U_and_29_nl)});
  assign nl_mul_loop_mul_16_FpMul_8U_23U_else_2_else_if_if_acc_nl = ({reg_FpMul_8U_23U_p_expo_itm
      , reg_FpMul_8U_23U_p_expo_2_itm_1}) + 8'b1;
  assign mul_loop_mul_16_FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_mul_loop_mul_16_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign FpMul_8U_23U_p_expo_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((mul_loop_mul_16_FpMul_8U_23U_else_2_else_if_if_acc_nl),
      ({reg_FpMul_8U_23U_p_expo_itm , reg_FpMul_8U_23U_p_expo_2_itm_1}), FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_15_itm_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_48_nl
      = ~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_15;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_lpi_1_dfm = MUX_v_23_2_2(FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_sva,
      23'b11111111111111111111111, (FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_FpMantWidthDec_8U_47U_23U_0U_0U_if_1_not_48_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_15 = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1 = FpMul_8U_23U_p_expo_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1[7:0];
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_sva = mul_loop_mul_16_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_sva_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_sva = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_sva[22:0];
  assign FpMul_8U_23U_o_expo_3_0_lpi_1_dfm_mx1 = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_lpi_1_dfm_1[3:0]),
      or_tmp_2118);
  assign FpMul_8U_23U_lor_2_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_7_4_lpi_1_dfm!=4'b0000)
      | (FpMul_8U_23U_o_expo_3_0_lpi_1_dfm_mx1!=4'b0000))) | FpMul_8U_23U_lor_1_lpi_1_dfm_7;
  assign FpMul_8U_23U_o_expo_7_4_lpi_1_dfm = MUX_v_4_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_lpi_1_dfm_1[7:4]),
      4'b1111, FpMul_8U_23U_is_inf_lpi_1_dfm_2);
  assign FpMul_8U_23U_is_inf_lpi_1_dfm_2 = ~(FpMul_8U_23U_FpMul_8U_23U_and_78_itm_2
      | FpMul_8U_23U_lor_1_lpi_1_dfm_7);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_30_nl = (~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_15)
      & mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_31_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_15
      & mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_lpi_1_dfm_1 = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1, {(~ mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs_2)
      , (FpMantWidthDec_8U_47U_23U_0U_0U_and_30_nl) , (FpMantWidthDec_8U_47U_23U_0U_0U_and_31_nl)});
  assign and_116_ssc = (~ mul_loop_mul_if_land_1_lpi_1_dfm_10) & nor_m1c;
  assign or_17_ssc = (mul_loop_mul_if_land_1_lpi_1_dfm_10 & nor_m1c) | (mul_loop_mul_else_land_1_lpi_1_dfm_10
      & and_1_m1c) | io_read_cfg_mul_bypass_rsc_svs_8;
  assign and_1_m1c = else_unequal_tmp & (~ io_read_cfg_mul_bypass_rsc_svs_8);
  assign nor_m1c = ~(else_unequal_tmp | io_read_cfg_mul_bypass_rsc_svs_8);
  assign and_51_ssc = (~ mul_loop_mul_if_land_2_lpi_1_dfm_10) & nor_m1c;
  assign or_1_ssc = (mul_loop_mul_if_land_2_lpi_1_dfm_10 & nor_m1c) | (mul_loop_mul_else_land_2_lpi_1_dfm_10
      & and_1_m1c) | io_read_cfg_mul_bypass_rsc_svs_8;
  assign and_55_ssc = (~ mul_loop_mul_if_land_3_lpi_1_dfm_10) & nor_m1c;
  assign or_2_ssc = (mul_loop_mul_if_land_3_lpi_1_dfm_10 & nor_m1c) | (mul_loop_mul_else_land_3_lpi_1_dfm_10
      & and_1_m1c) | io_read_cfg_mul_bypass_rsc_svs_8;
  assign and_59_ssc = (~ mul_loop_mul_if_land_4_lpi_1_dfm_10) & nor_m1c;
  assign or_3_ssc = (mul_loop_mul_if_land_4_lpi_1_dfm_10 & nor_m1c) | (mul_loop_mul_else_land_4_lpi_1_dfm_10
      & and_1_m1c) | io_read_cfg_mul_bypass_rsc_svs_8;
  assign and_63_ssc = (~ mul_loop_mul_if_land_5_lpi_1_dfm_10) & nor_m1c;
  assign or_4_ssc = (mul_loop_mul_if_land_5_lpi_1_dfm_10 & nor_m1c) | (mul_loop_mul_else_land_5_lpi_1_dfm_10
      & and_1_m1c) | io_read_cfg_mul_bypass_rsc_svs_8;
  assign and_67_ssc = (~ mul_loop_mul_if_land_6_lpi_1_dfm_10) & nor_m1c;
  assign or_5_ssc = (mul_loop_mul_if_land_6_lpi_1_dfm_10 & nor_m1c) | (mul_loop_mul_else_land_6_lpi_1_dfm_10
      & and_1_m1c) | io_read_cfg_mul_bypass_rsc_svs_8;
  assign and_71_ssc = (~ mul_loop_mul_if_land_7_lpi_1_dfm_10) & nor_m1c;
  assign or_6_ssc = (mul_loop_mul_if_land_7_lpi_1_dfm_10 & nor_m1c) | (mul_loop_mul_else_land_7_lpi_1_dfm_10
      & and_1_m1c) | io_read_cfg_mul_bypass_rsc_svs_8;
  assign and_75_ssc = (~ mul_loop_mul_if_land_8_lpi_1_dfm_10) & nor_m1c;
  assign or_7_ssc = (mul_loop_mul_if_land_8_lpi_1_dfm_10 & nor_m1c) | (mul_loop_mul_else_land_8_lpi_1_dfm_10
      & and_1_m1c) | io_read_cfg_mul_bypass_rsc_svs_8;
  assign and_79_ssc = (~ mul_loop_mul_if_land_9_lpi_1_dfm_10) & nor_m1c;
  assign or_8_ssc = (mul_loop_mul_if_land_9_lpi_1_dfm_10 & nor_m1c) | (mul_loop_mul_else_land_9_lpi_1_dfm_10
      & and_1_m1c) | io_read_cfg_mul_bypass_rsc_svs_8;
  assign and_83_ssc = (~ mul_loop_mul_if_land_10_lpi_1_dfm_10) & nor_m1c;
  assign or_9_ssc = (mul_loop_mul_if_land_10_lpi_1_dfm_10 & nor_m1c) | (mul_loop_mul_else_land_10_lpi_1_dfm_10
      & and_1_m1c) | io_read_cfg_mul_bypass_rsc_svs_8;
  assign and_87_ssc = (~ mul_loop_mul_if_land_11_lpi_1_dfm_10) & nor_m1c;
  assign or_10_ssc = (mul_loop_mul_if_land_11_lpi_1_dfm_10 & nor_m1c) | (mul_loop_mul_else_land_11_lpi_1_dfm_10
      & and_1_m1c) | io_read_cfg_mul_bypass_rsc_svs_8;
  assign and_91_ssc = (~ mul_loop_mul_if_land_12_lpi_1_dfm_10) & nor_m1c;
  assign or_11_ssc = (mul_loop_mul_if_land_12_lpi_1_dfm_10 & nor_m1c) | (mul_loop_mul_else_land_12_lpi_1_dfm_10
      & and_1_m1c) | io_read_cfg_mul_bypass_rsc_svs_8;
  assign and_95_ssc = (~ mul_loop_mul_if_land_13_lpi_1_dfm_10) & nor_m1c;
  assign or_12_ssc = (mul_loop_mul_if_land_13_lpi_1_dfm_10 & nor_m1c) | (mul_loop_mul_else_land_13_lpi_1_dfm_10
      & and_1_m1c) | io_read_cfg_mul_bypass_rsc_svs_8;
  assign and_99_ssc = (~ mul_loop_mul_if_land_14_lpi_1_dfm_10) & nor_m1c;
  assign or_13_ssc = (mul_loop_mul_if_land_14_lpi_1_dfm_10 & nor_m1c) | (mul_loop_mul_else_land_14_lpi_1_dfm_10
      & and_1_m1c) | io_read_cfg_mul_bypass_rsc_svs_8;
  assign and_103_ssc = (~ mul_loop_mul_if_land_15_lpi_1_dfm_10) & nor_m1c;
  assign or_14_ssc = (mul_loop_mul_if_land_15_lpi_1_dfm_10 & nor_m1c) | (mul_loop_mul_else_land_15_lpi_1_dfm_10
      & and_1_m1c) | io_read_cfg_mul_bypass_rsc_svs_8;
  assign and_107_ssc = (~ mul_loop_mul_if_land_lpi_1_dfm_10) & nor_m1c;
  assign or_15_ssc = (mul_loop_mul_if_land_lpi_1_dfm_10 & nor_m1c) | (mul_loop_mul_else_land_lpi_1_dfm_10
      & and_1_m1c) | io_read_cfg_mul_bypass_rsc_svs_8;
  assign main_stage_en_1 = chn_mul_in_rsci_bawt & (chn_mul_op_rsci_bawt | (~(cfg_mul_src_1_sva_st_1
      & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) & main_stage_v_1))) & (cfg_mul_src_rsc_triosy_obj_bawt
      | (~ main_stage_v_1)) & (cfg_mul_prelu_rsc_triosy_obj_bawt | (~ main_stage_v_1))
      & (cfg_mul_bypass_rsc_triosy_obj_bawt | (~ main_stage_v_1)) & (cfg_mul_op_rsc_triosy_obj_bawt
      | (~ main_stage_v_1)) & or_309_cse;
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_sva_1 = conv_u2u_3_4({2'b11
      , (mul_nan_to_zero_op_expo_1_lpi_1_dfm[4])}) + 4'b1;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_sva_1 = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_sva_1[3:0];
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_1_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_16)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_1_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_1_sva[5:0];
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_ssc =
      ~(IsDenorm_5U_23U_land_1_lpi_1_dfm | IsInf_5U_23U_land_1_lpi_1_dfm);
  assign IsInf_5U_23U_land_1_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_1_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_1_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_cse);
  assign IsNaN_5U_23U_nor_tmp = ~((mul_nan_to_zero_op_mant_1_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_1_lpi_1_dfm = ~(IsNaN_5U_23U_nor_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_cse);
  assign IsNaN_5U_23U_aelse_not_32_nl = ~ IsNaN_5U_23U_land_1_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_1_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_1_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_32_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_1_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_1_lpi_1_dfm, IsNaN_5U_23U_land_1_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_cse = ~((mul_nan_to_zero_op_expo_1_lpi_1_dfm==5'b11111));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_sva_1 = conv_u2u_3_4({2'b11
      , (mul_nan_to_zero_op_expo_2_lpi_1_dfm[4])}) + 4'b1;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_sva_1 = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_sva_1[3:0];
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_2_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_17)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_2_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_2_sva[5:0];
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_2_ssc
      = ~(IsDenorm_5U_23U_land_2_lpi_1_dfm | IsInf_5U_23U_land_2_lpi_1_dfm);
  assign IsInf_5U_23U_land_2_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_2_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_2_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_1_cse);
  assign IsNaN_5U_23U_nor_1_tmp = ~((mul_nan_to_zero_op_mant_2_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_2_lpi_1_dfm = ~(IsNaN_5U_23U_nor_1_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_1_cse);
  assign IsNaN_5U_23U_aelse_not_33_nl = ~ IsNaN_5U_23U_land_2_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_2_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_2_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_33_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_2_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_2_lpi_1_dfm, IsNaN_5U_23U_land_2_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_1_cse = ~((mul_nan_to_zero_op_expo_2_lpi_1_dfm==5'b11111));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_sva_1 = conv_u2u_3_4({2'b11
      , (mul_nan_to_zero_op_expo_3_lpi_1_dfm[4])}) + 4'b1;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_sva_1 = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_sva_1[3:0];
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_3_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_18)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_3_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_3_sva[5:0];
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_4_ssc
      = ~(IsDenorm_5U_23U_land_3_lpi_1_dfm | IsInf_5U_23U_land_3_lpi_1_dfm);
  assign IsInf_5U_23U_land_3_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_3_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_3_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_2_cse);
  assign IsNaN_5U_23U_nor_2_tmp = ~((mul_nan_to_zero_op_mant_3_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_3_lpi_1_dfm = ~(IsNaN_5U_23U_nor_2_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_2_cse);
  assign IsNaN_5U_23U_aelse_not_34_nl = ~ IsNaN_5U_23U_land_3_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_3_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_3_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_34_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_3_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_3_lpi_1_dfm, IsNaN_5U_23U_land_3_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_2_cse = ~((mul_nan_to_zero_op_expo_3_lpi_1_dfm==5'b11111));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_sva_1 = conv_u2u_3_4({2'b11
      , (mul_nan_to_zero_op_expo_4_lpi_1_dfm[4])}) + 4'b1;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_sva_1 = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_sva_1[3:0];
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_4_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_19)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_4_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_4_sva[5:0];
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_6_ssc
      = ~(IsDenorm_5U_23U_land_4_lpi_1_dfm | IsInf_5U_23U_land_4_lpi_1_dfm);
  assign IsInf_5U_23U_land_4_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_4_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_4_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_3_cse);
  assign IsNaN_5U_23U_nor_3_tmp = ~((mul_nan_to_zero_op_mant_4_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_4_lpi_1_dfm = ~(IsNaN_5U_23U_nor_3_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_3_cse);
  assign IsNaN_5U_23U_aelse_not_35_nl = ~ IsNaN_5U_23U_land_4_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_4_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_4_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_35_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_4_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_4_lpi_1_dfm, IsNaN_5U_23U_land_4_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_3_cse = ~((mul_nan_to_zero_op_expo_4_lpi_1_dfm==5'b11111));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_sva_1 = conv_u2u_3_4({2'b11
      , (mul_nan_to_zero_op_expo_5_lpi_1_dfm[4])}) + 4'b1;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_sva_1 = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_sva_1[3:0];
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_5_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_20)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_5_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_5_sva[5:0];
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_8_ssc
      = ~(IsDenorm_5U_23U_land_5_lpi_1_dfm | IsInf_5U_23U_land_5_lpi_1_dfm);
  assign IsInf_5U_23U_land_5_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_5_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_5_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_4_cse);
  assign IsNaN_5U_23U_nor_4_tmp = ~((mul_nan_to_zero_op_mant_5_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_5_lpi_1_dfm = ~(IsNaN_5U_23U_nor_4_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_4_cse);
  assign IsNaN_5U_23U_aelse_not_36_nl = ~ IsNaN_5U_23U_land_5_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_5_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_5_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_36_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_5_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_5_lpi_1_dfm, IsNaN_5U_23U_land_5_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_4_cse = ~((mul_nan_to_zero_op_expo_5_lpi_1_dfm==5'b11111));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_sva_1 = conv_u2u_3_4({2'b11
      , (mul_nan_to_zero_op_expo_6_lpi_1_dfm[4])}) + 4'b1;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_sva_1 = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_sva_1[3:0];
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_6_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_21)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_6_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_6_sva[5:0];
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_10_ssc
      = ~(IsDenorm_5U_23U_land_6_lpi_1_dfm | IsInf_5U_23U_land_6_lpi_1_dfm);
  assign IsInf_5U_23U_land_6_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_6_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_6_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_5_cse);
  assign IsNaN_5U_23U_nor_5_tmp = ~((mul_nan_to_zero_op_mant_6_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_6_lpi_1_dfm = ~(IsNaN_5U_23U_nor_5_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_5_cse);
  assign IsNaN_5U_23U_aelse_not_37_nl = ~ IsNaN_5U_23U_land_6_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_6_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_6_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_37_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_6_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_6_lpi_1_dfm, IsNaN_5U_23U_land_6_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_5_cse = ~((mul_nan_to_zero_op_expo_6_lpi_1_dfm==5'b11111));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_sva_1 = conv_u2u_3_4({2'b11
      , (mul_nan_to_zero_op_expo_7_lpi_1_dfm[4])}) + 4'b1;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_sva_1 = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_sva_1[3:0];
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_7_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_22)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_7_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_7_sva[5:0];
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_12_ssc
      = ~(IsDenorm_5U_23U_land_7_lpi_1_dfm | IsInf_5U_23U_land_7_lpi_1_dfm);
  assign IsInf_5U_23U_land_7_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_7_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_7_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_6_cse);
  assign IsNaN_5U_23U_nor_6_tmp = ~((mul_nan_to_zero_op_mant_7_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_7_lpi_1_dfm = ~(IsNaN_5U_23U_nor_6_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_6_cse);
  assign IsNaN_5U_23U_aelse_not_38_nl = ~ IsNaN_5U_23U_land_7_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_7_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_7_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_38_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_7_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_7_lpi_1_dfm, IsNaN_5U_23U_land_7_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_6_cse = ~((mul_nan_to_zero_op_expo_7_lpi_1_dfm==5'b11111));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_sva_1 = conv_u2u_3_4({2'b11
      , (mul_nan_to_zero_op_expo_8_lpi_1_dfm[4])}) + 4'b1;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_sva_1 = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_sva_1[3:0];
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_8_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_23)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_8_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_8_sva[5:0];
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_14_ssc
      = ~(IsDenorm_5U_23U_land_8_lpi_1_dfm | IsInf_5U_23U_land_8_lpi_1_dfm);
  assign IsInf_5U_23U_land_8_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_8_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_8_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_7_cse);
  assign IsNaN_5U_23U_nor_7_tmp = ~((mul_nan_to_zero_op_mant_8_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_8_lpi_1_dfm = ~(IsNaN_5U_23U_nor_7_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_7_cse);
  assign IsNaN_5U_23U_aelse_not_39_nl = ~ IsNaN_5U_23U_land_8_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_8_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_8_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_39_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_8_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_8_lpi_1_dfm, IsNaN_5U_23U_land_8_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_7_cse = ~((mul_nan_to_zero_op_expo_8_lpi_1_dfm==5'b11111));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_sva_1 = conv_u2u_3_4({2'b11
      , (mul_nan_to_zero_op_expo_9_lpi_1_dfm[4])}) + 4'b1;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_sva_1 = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_sva_1[3:0];
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_9_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_24)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_9_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_9_sva[5:0];
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_16_ssc
      = ~(IsDenorm_5U_23U_land_9_lpi_1_dfm | IsInf_5U_23U_land_9_lpi_1_dfm);
  assign IsInf_5U_23U_land_9_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_9_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_9_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_8_cse);
  assign IsNaN_5U_23U_nor_8_tmp = ~((mul_nan_to_zero_op_mant_9_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_9_lpi_1_dfm = ~(IsNaN_5U_23U_nor_8_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_8_cse);
  assign IsNaN_5U_23U_aelse_not_40_nl = ~ IsNaN_5U_23U_land_9_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_9_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_9_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_40_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_9_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_9_lpi_1_dfm, IsNaN_5U_23U_land_9_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_8_cse = ~((mul_nan_to_zero_op_expo_9_lpi_1_dfm==5'b11111));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_sva_1 = conv_u2u_3_4({2'b11
      , (mul_nan_to_zero_op_expo_10_lpi_1_dfm[4])}) + 4'b1;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_sva_1 = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_sva_1[3:0];
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_10_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_25)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_10_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_10_sva[5:0];
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_18_ssc
      = ~(IsDenorm_5U_23U_land_10_lpi_1_dfm | IsInf_5U_23U_land_10_lpi_1_dfm);
  assign IsInf_5U_23U_land_10_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_10_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_10_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_9_cse);
  assign IsNaN_5U_23U_nor_9_tmp = ~((mul_nan_to_zero_op_mant_10_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_10_lpi_1_dfm = ~(IsNaN_5U_23U_nor_9_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_9_cse);
  assign IsNaN_5U_23U_aelse_not_41_nl = ~ IsNaN_5U_23U_land_10_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_10_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_10_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_41_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_10_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_10_lpi_1_dfm, IsNaN_5U_23U_land_10_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_9_cse = ~((mul_nan_to_zero_op_expo_10_lpi_1_dfm==5'b11111));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_sva_1 = conv_u2u_3_4({2'b11
      , (mul_nan_to_zero_op_expo_11_lpi_1_dfm[4])}) + 4'b1;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_sva_1 = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_sva_1[3:0];
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_11_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_26)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_11_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_11_sva[5:0];
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_20_ssc
      = ~(IsDenorm_5U_23U_land_11_lpi_1_dfm | IsInf_5U_23U_land_11_lpi_1_dfm);
  assign IsInf_5U_23U_land_11_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_11_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_11_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_10_cse);
  assign IsNaN_5U_23U_nor_10_tmp = ~((mul_nan_to_zero_op_mant_11_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_11_lpi_1_dfm = ~(IsNaN_5U_23U_nor_10_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_10_cse);
  assign IsNaN_5U_23U_aelse_not_42_nl = ~ IsNaN_5U_23U_land_11_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_11_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_11_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_42_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_11_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_11_lpi_1_dfm, IsNaN_5U_23U_land_11_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_10_cse = ~((mul_nan_to_zero_op_expo_11_lpi_1_dfm==5'b11111));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_sva_1 = conv_u2u_3_4({2'b11
      , (mul_nan_to_zero_op_expo_12_lpi_1_dfm[4])}) + 4'b1;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_sva_1 = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_sva_1[3:0];
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_12_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_27)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_12_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_12_sva[5:0];
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_22_ssc
      = ~(IsDenorm_5U_23U_land_12_lpi_1_dfm | IsInf_5U_23U_land_12_lpi_1_dfm);
  assign IsInf_5U_23U_land_12_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_12_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_12_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_11_cse);
  assign IsNaN_5U_23U_nor_11_tmp = ~((mul_nan_to_zero_op_mant_12_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_12_lpi_1_dfm = ~(IsNaN_5U_23U_nor_11_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_11_cse);
  assign IsNaN_5U_23U_aelse_not_43_nl = ~ IsNaN_5U_23U_land_12_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_12_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_12_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_43_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_12_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_12_lpi_1_dfm, IsNaN_5U_23U_land_12_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_11_cse = ~((mul_nan_to_zero_op_expo_12_lpi_1_dfm==5'b11111));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_sva_1 = conv_u2u_3_4({2'b11
      , (mul_nan_to_zero_op_expo_13_lpi_1_dfm[4])}) + 4'b1;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_sva_1 = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_sva_1[3:0];
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_13_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_28)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_13_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_13_sva[5:0];
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_24_ssc
      = ~(IsDenorm_5U_23U_land_13_lpi_1_dfm | IsInf_5U_23U_land_13_lpi_1_dfm);
  assign IsInf_5U_23U_land_13_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_13_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_13_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_12_cse);
  assign IsNaN_5U_23U_nor_12_tmp = ~((mul_nan_to_zero_op_mant_13_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_13_lpi_1_dfm = ~(IsNaN_5U_23U_nor_12_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_12_cse);
  assign IsNaN_5U_23U_aelse_not_44_nl = ~ IsNaN_5U_23U_land_13_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_13_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_13_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_44_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_13_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_13_lpi_1_dfm, IsNaN_5U_23U_land_13_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_12_cse = ~((mul_nan_to_zero_op_expo_13_lpi_1_dfm==5'b11111));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_sva_1 = conv_u2u_3_4({2'b11
      , (mul_nan_to_zero_op_expo_14_lpi_1_dfm[4])}) + 4'b1;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_sva_1 = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_sva_1[3:0];
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_14_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_29)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_14_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_14_sva[5:0];
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_26_ssc
      = ~(IsDenorm_5U_23U_land_14_lpi_1_dfm | IsInf_5U_23U_land_14_lpi_1_dfm);
  assign IsInf_5U_23U_land_14_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_14_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_14_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_13_cse);
  assign IsNaN_5U_23U_nor_13_tmp = ~((mul_nan_to_zero_op_mant_14_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_14_lpi_1_dfm = ~(IsNaN_5U_23U_nor_13_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_13_cse);
  assign IsNaN_5U_23U_aelse_not_45_nl = ~ IsNaN_5U_23U_land_14_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_14_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_14_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_45_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_14_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_14_lpi_1_dfm, IsNaN_5U_23U_land_14_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_13_cse = ~((mul_nan_to_zero_op_expo_14_lpi_1_dfm==5'b11111));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_sva_1 = conv_u2u_3_4({2'b11
      , (mul_nan_to_zero_op_expo_15_lpi_1_dfm[4])}) + 4'b1;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_sva_1 = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_sva_1[3:0];
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_15_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_30)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_15_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_15_sva[5:0];
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_28_ssc
      = ~(IsDenorm_5U_23U_land_15_lpi_1_dfm | IsInf_5U_23U_land_15_lpi_1_dfm);
  assign IsInf_5U_23U_land_15_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_15_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_15_lpi_1_dfm!=10'b0000000000)
      | IsNaN_5U_23U_IsNaN_5U_23U_nand_14_cse);
  assign IsNaN_5U_23U_nor_14_tmp = ~((mul_nan_to_zero_op_mant_15_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_15_lpi_1_dfm = ~(IsNaN_5U_23U_nor_14_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_14_cse);
  assign IsNaN_5U_23U_aelse_not_46_nl = ~ IsNaN_5U_23U_land_15_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_15_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_15_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_46_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_15_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_15_lpi_1_dfm, IsNaN_5U_23U_land_15_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_14_cse = ~((mul_nan_to_zero_op_expo_15_lpi_1_dfm==5'b11111));
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_sva_1 = conv_u2u_3_4({2'b11
      , (mul_nan_to_zero_op_expo_lpi_1_dfm[4])}) + 4'b1;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_sva_1 = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_sva_1[3:0];
  assign nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_sva = ({1'b1 , (~ libraries_leading_sign_23_0_5aae14ba1d9c4916020dde6af2ddf1395444_31)})
      + 6'b110001;
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_sva = nl_FpExpoWidthInc_5U_8U_23U_1U_1U_if_1_if_acc_psp_sva[5:0];
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_nor_30_ssc
      = ~(IsDenorm_5U_23U_land_lpi_1_dfm | IsInf_5U_23U_land_lpi_1_dfm);
  assign IsInf_5U_23U_land_lpi_1_dfm = ~((FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_lpi_1_dfm!=10'b0000000000) |
      IsNaN_5U_23U_IsNaN_5U_23U_nand_15_cse);
  assign IsNaN_5U_23U_nor_15_tmp = ~((mul_nan_to_zero_op_mant_lpi_1_dfm!=10'b0000000000));
  assign IsNaN_5U_23U_land_lpi_1_dfm = ~(IsNaN_5U_23U_nor_15_tmp | IsNaN_5U_23U_IsNaN_5U_23U_nand_15_cse);
  assign IsNaN_5U_23U_aelse_not_47_nl = ~ IsNaN_5U_23U_land_lpi_1_dfm;
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_lpi_1_dfm, (IsNaN_5U_23U_aelse_not_47_nl));
  assign FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      mul_nan_to_zero_op_mant_lpi_1_dfm, IsNaN_5U_23U_land_lpi_1_dfm);
  assign IsNaN_5U_23U_IsNaN_5U_23U_nand_15_cse = ~((mul_nan_to_zero_op_expo_lpi_1_dfm==5'b11111));
  assign nl_mul_loop_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_1_sva_1_mx0w0[7:1])})
      + 8'b1;
  assign mul_loop_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_mul_loop_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign mul_loop_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 = readslicef_8_1_7((mul_loop_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign or_4383_cse = (~ mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_18_lpi_1_dfm_st_3;
  assign mux_1664_nl = MUX_s_1_2_2((mul_loop_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
      (FpMul_8U_23U_p_mant_p1_1_sva[47]), or_4383_cse);
  assign FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_1_sva_mx1[45:0]),
      (FpMul_8U_23U_p_mant_p1_1_sva_mx1[46:1]), mux_1664_nl);
  assign nl_mul_loop_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_2_sva_1_mx0w0[7:1])})
      + 8'b1;
  assign mul_loop_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_mul_loop_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign mul_loop_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 = readslicef_8_1_7((mul_loop_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign or_4384_cse = (~ mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_19_lpi_1_dfm_st_3;
  assign mux_1665_nl = MUX_s_1_2_2((mul_loop_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
      (FpMul_8U_23U_p_mant_p1_2_sva[47]), or_4384_cse);
  assign FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_2_sva_mx1[45:0]),
      (FpMul_8U_23U_p_mant_p1_2_sva_mx1[46:1]), mux_1665_nl);
  assign nl_mul_loop_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_3_sva_1_mx0w0[7:1])})
      + 8'b1;
  assign mul_loop_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_mul_loop_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign mul_loop_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 = readslicef_8_1_7((mul_loop_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign or_4385_cse = (~ mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_20_lpi_1_dfm_st_3;
  assign mux_1666_nl = MUX_s_1_2_2((mul_loop_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
      (FpMul_8U_23U_p_mant_p1_3_sva[47]), or_4385_cse);
  assign FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_3_sva_mx1[45:0]),
      (FpMul_8U_23U_p_mant_p1_3_sva_mx1[46:1]), mux_1666_nl);
  assign nl_mul_loop_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_4_sva_1_mx0w0[7:1])})
      + 8'b1;
  assign mul_loop_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_mul_loop_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign mul_loop_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 = readslicef_8_1_7((mul_loop_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign mux_1667_nl = MUX_s_1_2_2((mul_loop_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
      (FpMul_8U_23U_p_mant_p1_4_sva[47]), or_1253_cse);
  assign FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_4_sva_mx1[45:0]),
      (FpMul_8U_23U_p_mant_p1_4_sva_mx1[46:1]), mux_1667_nl);
  assign nl_mul_loop_mul_5_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_5_sva_1_mx0w0[7:1])})
      + 8'b1;
  assign mul_loop_mul_5_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_mul_loop_mul_5_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign mul_loop_mul_5_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 = readslicef_8_1_7((mul_loop_mul_5_FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign or_4387_cse = (~ mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_22_lpi_1_dfm_st_3;
  assign mux_1668_nl = MUX_s_1_2_2((mul_loop_mul_5_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
      (FpMul_8U_23U_p_mant_p1_5_sva[47]), or_4387_cse);
  assign FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_5_sva_mx1[45:0]),
      (FpMul_8U_23U_p_mant_p1_5_sva_mx1[46:1]), mux_1668_nl);
  assign nl_mul_loop_mul_6_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_6_sva_1_mx0w0[7:1])})
      + 8'b1;
  assign mul_loop_mul_6_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_mul_loop_mul_6_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign mul_loop_mul_6_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 = readslicef_8_1_7((mul_loop_mul_6_FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign mux_1669_nl = MUX_s_1_2_2((mul_loop_mul_6_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
      (FpMul_8U_23U_p_mant_p1_6_sva[47]), or_2342_cse);
  assign FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_6_sva_mx1[45:0]),
      (FpMul_8U_23U_p_mant_p1_6_sva_mx1[46:1]), mux_1669_nl);
  assign nl_mul_loop_mul_7_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_7_sva_1_mx0w0[7:1])})
      + 8'b1;
  assign mul_loop_mul_7_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_mul_loop_mul_7_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign mul_loop_mul_7_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 = readslicef_8_1_7((mul_loop_mul_7_FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign or_4389_cse = (~ mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_24_lpi_1_dfm_st_3;
  assign mux_1670_nl = MUX_s_1_2_2((mul_loop_mul_7_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
      (FpMul_8U_23U_p_mant_p1_7_sva[47]), or_4389_cse);
  assign FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_7_sva_mx1[45:0]),
      (FpMul_8U_23U_p_mant_p1_7_sva_mx1[46:1]), mux_1670_nl);
  assign nl_mul_loop_mul_8_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_8_sva_1_mx0w0[7:1])})
      + 8'b1;
  assign mul_loop_mul_8_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_mul_loop_mul_8_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign mul_loop_mul_8_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 = readslicef_8_1_7((mul_loop_mul_8_FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign or_4390_cse = (~ mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_25_lpi_1_dfm_st_3;
  assign mux_1671_nl = MUX_s_1_2_2((mul_loop_mul_8_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
      (FpMul_8U_23U_p_mant_p1_8_sva[47]), or_4390_cse);
  assign FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_8_sva_mx1[45:0]),
      (FpMul_8U_23U_p_mant_p1_8_sva_mx1[46:1]), mux_1671_nl);
  assign nl_mul_loop_mul_9_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_9_sva_1_mx0w0[7:1])})
      + 8'b1;
  assign mul_loop_mul_9_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_mul_loop_mul_9_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign mul_loop_mul_9_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 = readslicef_8_1_7((mul_loop_mul_9_FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign or_4391_cse = (~ mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_26_lpi_1_dfm_st_3;
  assign mux_1672_nl = MUX_s_1_2_2((mul_loop_mul_9_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
      (FpMul_8U_23U_p_mant_p1_9_sva[47]), or_4391_cse);
  assign FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_9_sva_mx1[45:0]),
      (FpMul_8U_23U_p_mant_p1_9_sva_mx1[46:1]), mux_1672_nl);
  assign nl_mul_loop_mul_10_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_10_sva_1_mx0w0[7:1])})
      + 8'b1;
  assign mul_loop_mul_10_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_mul_loop_mul_10_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign mul_loop_mul_10_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 = readslicef_8_1_7((mul_loop_mul_10_FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign mux_1673_nl = MUX_s_1_2_2((mul_loop_mul_10_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
      (FpMul_8U_23U_p_mant_p1_10_sva[47]), or_2386_cse);
  assign FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_10_sva_mx1[45:0]),
      (FpMul_8U_23U_p_mant_p1_10_sva_mx1[46:1]), mux_1673_nl);
  assign nl_mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_11_sva_1_mx0w0[7:1])})
      + 8'b1;
  assign mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 = readslicef_8_1_7((mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign nor_606_nl = ~((~ or_1819_cse) | (FpMul_8U_23U_p_mant_p1_11_sva[47]));
  assign nand_170_nl = ~(or_1819_cse & (FpMul_8U_23U_p_mant_p1_11_sva[47]));
  assign mux_1674_nl = MUX_s_1_2_2((nand_170_nl), (nor_606_nl), mul_loop_mul_11_FpMul_8U_23U_p_mant_p1_mul_tmp[47]);
  assign FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_11_sva_mx1[46:1]),
      (FpMul_8U_23U_p_mant_p1_11_sva_mx1[45:0]), mux_1674_nl);
  assign nl_mul_loop_mul_12_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_12_sva_1_mx0w0[7:1])})
      + 8'b1;
  assign mul_loop_mul_12_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_mul_loop_mul_12_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign mul_loop_mul_12_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 = readslicef_8_1_7((mul_loop_mul_12_FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign mux_1675_nl = MUX_s_1_2_2((mul_loop_mul_12_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
      (FpMul_8U_23U_p_mant_p1_12_sva[47]), or_1898_cse);
  assign FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_12_sva_mx1[45:0]),
      (FpMul_8U_23U_p_mant_p1_12_sva_mx1[46:1]), mux_1675_nl);
  assign nl_mul_loop_mul_13_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_13_sva_1_mx0w0[7:1])})
      + 8'b1;
  assign mul_loop_mul_13_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_mul_loop_mul_13_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign mul_loop_mul_13_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 = readslicef_8_1_7((mul_loop_mul_13_FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign mux_1676_nl = MUX_s_1_2_2((mul_loop_mul_13_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
      (FpMul_8U_23U_p_mant_p1_13_sva[47]), or_1981_cse);
  assign FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_13_sva_mx1[45:0]),
      (FpMul_8U_23U_p_mant_p1_13_sva_mx1[46:1]), mux_1676_nl);
  assign nl_mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_14_sva_1_mx0w0[7:1])})
      + 8'b1;
  assign mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 = readslicef_8_1_7((mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign or_4398_cse = (~ mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_31_lpi_1_dfm_st_3;
  assign mux_1677_nl = MUX_s_1_2_2((mul_loop_mul_14_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
      (FpMul_8U_23U_p_mant_p1_14_sva[47]), or_4398_cse);
  assign FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_14_sva_mx1[45:0]),
      (FpMul_8U_23U_p_mant_p1_14_sva_mx1[46:1]), mux_1677_nl);
  assign nl_mul_loop_mul_15_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_15_sva_1_mx0w0[7:1])})
      + 8'b1;
  assign mul_loop_mul_15_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_mul_loop_mul_15_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign mul_loop_mul_15_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 = readslicef_8_1_7((mul_loop_mul_15_FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign or_4399_cse = (~ mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_32_lpi_1_dfm_st_3;
  assign mux_1678_nl = MUX_s_1_2_2((mul_loop_mul_15_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
      (FpMul_8U_23U_p_mant_p1_15_sva[47]), or_4399_cse);
  assign FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_15_sva_mx1[45:0]),
      (FpMul_8U_23U_p_mant_p1_15_sva_mx1[46:1]), mux_1678_nl);
  assign nl_mul_loop_mul_16_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_sva_1_mx0w0[7:1])})
      + 8'b1;
  assign mul_loop_mul_16_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_mul_loop_mul_16_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign mul_loop_mul_16_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 = readslicef_8_1_7((mul_loop_mul_16_FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign or_4400_cse = (~ mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
  assign mux_1679_nl = MUX_s_1_2_2((mul_loop_mul_16_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
      (FpMul_8U_23U_p_mant_p1_sva[47]), or_4400_cse);
  assign FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_sva_mx1[45:0]),
      (FpMul_8U_23U_p_mant_p1_sva_mx1[46:1]), mux_1679_nl);
  assign else_MulOp_data_0_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_mul_op_1_sva_1[15]),
      (chn_mul_op_rsci_d_mxwt[15]), cfg_mul_src_1_sva_1);
  assign else_MulOp_data_1_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_mul_op_1_sva_1[15]),
      (chn_mul_op_rsci_d_mxwt[31]), cfg_mul_src_1_sva_1);
  assign else_MulOp_data_2_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_mul_op_1_sva_1[15]),
      (chn_mul_op_rsci_d_mxwt[47]), cfg_mul_src_1_sva_1);
  assign else_MulOp_data_3_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_mul_op_1_sva_1[15]),
      (chn_mul_op_rsci_d_mxwt[63]), cfg_mul_src_1_sva_1);
  assign else_MulOp_data_4_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_mul_op_1_sva_1[15]),
      (chn_mul_op_rsci_d_mxwt[79]), cfg_mul_src_1_sva_1);
  assign else_MulOp_data_5_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_mul_op_1_sva_1[15]),
      (chn_mul_op_rsci_d_mxwt[95]), cfg_mul_src_1_sva_1);
  assign else_MulOp_data_6_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_mul_op_1_sva_1[15]),
      (chn_mul_op_rsci_d_mxwt[111]), cfg_mul_src_1_sva_1);
  assign else_MulOp_data_7_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_mul_op_1_sva_1[15]),
      (chn_mul_op_rsci_d_mxwt[127]), cfg_mul_src_1_sva_1);
  assign else_MulOp_data_8_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_mul_op_1_sva_1[15]),
      (chn_mul_op_rsci_d_mxwt[143]), cfg_mul_src_1_sva_1);
  assign else_MulOp_data_9_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_mul_op_1_sva_1[15]),
      (chn_mul_op_rsci_d_mxwt[159]), cfg_mul_src_1_sva_1);
  assign else_MulOp_data_10_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_mul_op_1_sva_1[15]),
      (chn_mul_op_rsci_d_mxwt[175]), cfg_mul_src_1_sva_1);
  assign else_MulOp_data_11_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_mul_op_1_sva_1[15]),
      (chn_mul_op_rsci_d_mxwt[191]), cfg_mul_src_1_sva_1);
  assign else_MulOp_data_12_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_mul_op_1_sva_1[15]),
      (chn_mul_op_rsci_d_mxwt[207]), cfg_mul_src_1_sva_1);
  assign else_MulOp_data_13_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_mul_op_1_sva_1[15]),
      (chn_mul_op_rsci_d_mxwt[223]), cfg_mul_src_1_sva_1);
  assign else_MulOp_data_14_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_mul_op_1_sva_1[15]),
      (chn_mul_op_rsci_d_mxwt[239]), cfg_mul_src_1_sva_1);
  assign else_MulOp_data_15_15_lpi_1_dfm_mx0 = MUX_s_1_2_2((cfg_mul_op_1_sva_1[15]),
      (chn_mul_op_rsci_d_mxwt[255]), cfg_mul_src_1_sva_1);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_exs_261_0 = (mul_nan_to_zero_op_mant_1_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_1_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_exs_267_0 = (mul_nan_to_zero_op_mant_2_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_2_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_exs_273_0 = (mul_nan_to_zero_op_mant_3_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_3_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_exs_279_0 = (mul_nan_to_zero_op_mant_4_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_4_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_exs_285_0 = (mul_nan_to_zero_op_mant_5_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_5_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_exs_291_0 = (mul_nan_to_zero_op_mant_6_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_6_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_exs_297_0 = (mul_nan_to_zero_op_mant_7_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_7_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_exs_303_0 = (mul_nan_to_zero_op_mant_8_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_8_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_exs_309_0 = (mul_nan_to_zero_op_mant_9_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_9_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_exs_315_0 = (mul_nan_to_zero_op_mant_10_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_10_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_exs_321_0 = (mul_nan_to_zero_op_mant_11_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_11_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_exs_327_0 = (mul_nan_to_zero_op_mant_12_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_12_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_exs_333_0 = (mul_nan_to_zero_op_mant_13_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_13_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_exs_339_0 = (mul_nan_to_zero_op_mant_14_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_14_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_exs_345_0 = (mul_nan_to_zero_op_mant_15_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_15_sva);
  assign FpExpoWidthInc_5U_8U_23U_1U_1U_exs_351_0 = (mul_nan_to_zero_op_mant_lpi_1_dfm!=10'b0000000000)
      | (~ IsZero_5U_23U_IsZero_5U_23U_nor_cse_sva);
  assign asn_1163 = (~ mul_loop_mul_else_land_1_lpi_1_dfm_10) & and_1_m1c;
  assign asn_1165 = (~ IsNaN_8U_23U_land_1_lpi_1_dfm_11) & and_116_ssc;
  assign asn_1173 = (~ mul_loop_mul_else_land_2_lpi_1_dfm_10) & and_1_m1c;
  assign asn_1175 = (~ IsNaN_8U_23U_land_2_lpi_1_dfm_11) & and_51_ssc;
  assign asn_1183 = (~ mul_loop_mul_else_land_3_lpi_1_dfm_10) & and_1_m1c;
  assign asn_1185 = (~ IsNaN_8U_23U_land_3_lpi_1_dfm_11) & and_55_ssc;
  assign asn_1193 = (~ mul_loop_mul_else_land_4_lpi_1_dfm_10) & and_1_m1c;
  assign asn_1195 = (~ IsNaN_8U_23U_land_4_lpi_1_dfm_11) & and_59_ssc;
  assign asn_1203 = (~ mul_loop_mul_else_land_5_lpi_1_dfm_10) & and_1_m1c;
  assign asn_1205 = (~ IsNaN_8U_23U_land_5_lpi_1_dfm_11) & and_63_ssc;
  assign asn_1213 = (~ mul_loop_mul_else_land_6_lpi_1_dfm_10) & and_1_m1c;
  assign asn_1215 = (~ IsNaN_8U_23U_land_6_lpi_1_dfm_11) & and_67_ssc;
  assign asn_1223 = (~ mul_loop_mul_else_land_7_lpi_1_dfm_10) & and_1_m1c;
  assign asn_1225 = (~ IsNaN_8U_23U_land_7_lpi_1_dfm_11) & and_71_ssc;
  assign asn_1233 = (~ mul_loop_mul_else_land_8_lpi_1_dfm_10) & and_1_m1c;
  assign asn_1235 = (~ IsNaN_8U_23U_land_8_lpi_1_dfm_11) & and_75_ssc;
  assign asn_1243 = (~ mul_loop_mul_else_land_9_lpi_1_dfm_10) & and_1_m1c;
  assign asn_1245 = (~ IsNaN_8U_23U_land_9_lpi_1_dfm_11) & and_79_ssc;
  assign asn_1253 = (~ mul_loop_mul_else_land_10_lpi_1_dfm_10) & and_1_m1c;
  assign asn_1255 = (~ IsNaN_8U_23U_land_10_lpi_1_dfm_11) & and_83_ssc;
  assign asn_1263 = (~ mul_loop_mul_else_land_11_lpi_1_dfm_10) & and_1_m1c;
  assign asn_1265 = (~ IsNaN_8U_23U_land_11_lpi_1_dfm_11) & and_87_ssc;
  assign asn_1273 = (~ mul_loop_mul_else_land_12_lpi_1_dfm_10) & and_1_m1c;
  assign asn_1275 = (~ IsNaN_8U_23U_land_12_lpi_1_dfm_11) & and_91_ssc;
  assign asn_1283 = (~ mul_loop_mul_else_land_13_lpi_1_dfm_10) & and_1_m1c;
  assign asn_1285 = (~ IsNaN_8U_23U_land_13_lpi_1_dfm_11) & and_95_ssc;
  assign asn_1293 = (~ mul_loop_mul_else_land_14_lpi_1_dfm_10) & and_1_m1c;
  assign asn_1295 = (~ IsNaN_8U_23U_land_14_lpi_1_dfm_11) & and_99_ssc;
  assign asn_1303 = (~ mul_loop_mul_else_land_15_lpi_1_dfm_10) & and_1_m1c;
  assign asn_1305 = (~ IsNaN_8U_23U_land_15_lpi_1_dfm_11) & and_103_ssc;
  assign asn_1313 = (~ mul_loop_mul_else_land_lpi_1_dfm_10) & and_1_m1c;
  assign asn_1315 = (~ IsNaN_8U_23U_land_lpi_1_dfm_11) & and_107_ssc;
  assign else_mux_47_tmp = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]), (chn_mul_op_rsci_d_mxwt[254:250]),
      cfg_mul_src_1_sva_1);
  assign else_mux_44_tmp = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]), (chn_mul_op_rsci_d_mxwt[238:234]),
      cfg_mul_src_1_sva_1);
  assign else_mux_41_tmp = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]), (chn_mul_op_rsci_d_mxwt[222:218]),
      cfg_mul_src_1_sva_1);
  assign else_mux_38_tmp = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]), (chn_mul_op_rsci_d_mxwt[206:202]),
      cfg_mul_src_1_sva_1);
  assign else_mux_35_tmp = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]), (chn_mul_op_rsci_d_mxwt[190:186]),
      cfg_mul_src_1_sva_1);
  assign else_mux_32_tmp = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]), (chn_mul_op_rsci_d_mxwt[174:170]),
      cfg_mul_src_1_sva_1);
  assign else_mux_29_tmp = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]), (chn_mul_op_rsci_d_mxwt[158:154]),
      cfg_mul_src_1_sva_1);
  assign else_mux_26_tmp = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]), (chn_mul_op_rsci_d_mxwt[142:138]),
      cfg_mul_src_1_sva_1);
  assign else_mux_23_tmp = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]), (chn_mul_op_rsci_d_mxwt[126:122]),
      cfg_mul_src_1_sva_1);
  assign else_mux_20_tmp = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]), (chn_mul_op_rsci_d_mxwt[110:106]),
      cfg_mul_src_1_sva_1);
  assign else_mux_17_tmp = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]), (chn_mul_op_rsci_d_mxwt[94:90]),
      cfg_mul_src_1_sva_1);
  assign else_mux_14_tmp = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]), (chn_mul_op_rsci_d_mxwt[78:74]),
      cfg_mul_src_1_sva_1);
  assign else_mux_11_tmp = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]), (chn_mul_op_rsci_d_mxwt[62:58]),
      cfg_mul_src_1_sva_1);
  assign else_mux_8_tmp = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]), (chn_mul_op_rsci_d_mxwt[46:42]),
      cfg_mul_src_1_sva_1);
  assign else_mux_5_tmp = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]), (chn_mul_op_rsci_d_mxwt[30:26]),
      cfg_mul_src_1_sva_1);
  assign else_mux_2_tmp = MUX_v_5_2_2((cfg_mul_op_1_sva_1[14:10]), (chn_mul_op_rsci_d_mxwt[14:10]),
      cfg_mul_src_1_sva_1);
  assign and_dcpl_2 = (~(cfg_mul_bypass_rsci_d | (cfg_precision[0]))) & (cfg_precision[1])
      & chn_mul_in_rsci_bawt;
  assign and_dcpl_3 = cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt;
  assign and_dcpl_4 = cfg_mul_op_rsc_triosy_obj_bawt & cfg_mul_bypass_rsc_triosy_obj_bawt;
  assign and_dcpl_5 = and_dcpl_4 & and_dcpl_3;
  assign or_dcpl_4 = ~((~(and_dcpl_5 & or_4649_cse)) & main_stage_v_1);
  assign and_dcpl_7 = or_dcpl_4 & or_309_cse;
  assign or_tmp_4 = mul_loop_mul_if_land_1_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign or_tmp_5 = or_tmp_4 | (~ main_stage_v_1);
  assign or_4664_nl = mul_loop_mul_if_land_1_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | (~ main_stage_v_1) | and_dcpl_5;
  assign mux_7_nl = MUX_s_1_2_2(or_tmp_5, (or_4664_nl), or_2575_cse);
  assign mux_tmp_1 = MUX_s_1_2_2(or_tmp_5, (mux_7_nl), or_309_cse);
  assign nand_tmp_1 = ~(main_stage_v_1 & (~ and_dcpl_5));
  assign or_tmp_8 = cfg_mul_bypass_rsci_d | (~ nand_tmp_1);
  assign nand_tmp_2 = io_read_cfg_mul_bypass_rsc_svs_st_1 | (~ main_stage_v_1) |
      and_dcpl_5;
  assign not_tmp_8 = io_read_cfg_mul_bypass_rsc_svs_st_1 & main_stage_v_1 & (~ and_dcpl_5);
  assign mux_tmp_2 = MUX_s_1_2_2(not_tmp_8, nand_tmp_2, cfg_mul_bypass_rsci_d);
  assign mux_11_nl = MUX_s_1_2_2(main_stage_v_1, (~ nand_tmp_1), io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign or_tmp_9 = cfg_mul_bypass_rsci_d | (mux_11_nl);
  assign or_tmp_10 = io_read_cfg_mul_bypass_rsc_svs_st_1 | (~ main_stage_v_1);
  assign mux_tmp_5 = MUX_s_1_2_2(not_tmp_8, or_tmp_10, cfg_mul_bypass_rsci_d);
  assign mux_10_nl = MUX_s_1_2_2(mux_tmp_2, or_tmp_8, mul_loop_mul_if_land_1_lpi_1_dfm_st_5);
  assign mux_13_nl = MUX_s_1_2_2(mux_tmp_5, or_tmp_9, mul_loop_mul_if_land_1_lpi_1_dfm_st_5);
  assign mux_14_nl = MUX_s_1_2_2((mux_13_nl), (mux_10_nl), or_2575_cse);
  assign mux_tmp_8 = MUX_s_1_2_2(or_tmp_5, (mux_14_nl), or_309_cse);
  assign or_tmp_14 = mul_loop_mul_if_land_2_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign or_tmp_15 = or_tmp_14 | (~ main_stage_v_1);
  assign or_4662_nl = mul_loop_mul_if_land_2_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | (~ main_stage_v_1) | and_dcpl_5;
  assign mux_20_nl = MUX_s_1_2_2(or_tmp_15, (or_4662_nl), or_2575_cse);
  assign mux_tmp_14 = MUX_s_1_2_2(or_tmp_15, (mux_20_nl), or_309_cse);
  assign mux_22_nl = MUX_s_1_2_2(mux_tmp_2, or_tmp_8, mul_loop_mul_if_land_2_lpi_1_dfm_st_5);
  assign mux_23_nl = MUX_s_1_2_2(mux_tmp_5, or_tmp_9, mul_loop_mul_if_land_2_lpi_1_dfm_st_5);
  assign mux_24_nl = MUX_s_1_2_2((mux_23_nl), (mux_22_nl), or_2575_cse);
  assign mux_tmp_18 = MUX_s_1_2_2(or_tmp_15, (mux_24_nl), or_309_cse);
  assign or_tmp_21 = mul_loop_mul_if_land_3_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign or_tmp_22 = or_tmp_21 | (~ main_stage_v_1);
  assign or_4661_nl = mul_loop_mul_if_land_3_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | (~ main_stage_v_1) | and_dcpl_5;
  assign mux_30_nl = MUX_s_1_2_2(or_tmp_22, (or_4661_nl), or_2575_cse);
  assign mux_tmp_24 = MUX_s_1_2_2(or_tmp_22, (mux_30_nl), or_309_cse);
  assign mux_32_nl = MUX_s_1_2_2(mux_tmp_2, or_tmp_8, mul_loop_mul_if_land_3_lpi_1_dfm_st_5);
  assign mux_33_nl = MUX_s_1_2_2(mux_tmp_5, or_tmp_9, mul_loop_mul_if_land_3_lpi_1_dfm_st_5);
  assign mux_34_nl = MUX_s_1_2_2((mux_33_nl), (mux_32_nl), or_2575_cse);
  assign mux_tmp_28 = MUX_s_1_2_2(or_tmp_22, (mux_34_nl), or_309_cse);
  assign mux_tmp_33 = MUX_s_1_2_2(or_tmp_10, nand_tmp_2, or_2575_cse);
  assign or_tmp_29 = mul_loop_mul_if_land_4_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign or_tmp_30 = or_tmp_29 | (~ main_stage_v_1);
  assign or_117_nl = mul_loop_mul_if_land_4_lpi_1_dfm_st_5 | mux_tmp_33;
  assign mux_tmp_34 = MUX_s_1_2_2(or_tmp_30, (or_117_nl), or_309_cse);
  assign mux_tmp_35 = MUX_s_1_2_2(or_tmp_9, or_tmp_8, or_2575_cse);
  assign mux_tmp_36 = MUX_s_1_2_2(mux_tmp_5, mux_tmp_2, or_2575_cse);
  assign mux_44_nl = MUX_s_1_2_2(mux_tmp_36, mux_tmp_35, mul_loop_mul_if_land_4_lpi_1_dfm_st_5);
  assign mux_tmp_38 = MUX_s_1_2_2(or_tmp_30, (mux_44_nl), or_309_cse);
  assign or_tmp_37 = mul_loop_mul_if_land_5_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign or_tmp_38 = or_tmp_37 | (~ main_stage_v_1);
  assign or_4660_nl = mul_loop_mul_if_land_5_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | (~ main_stage_v_1) | and_dcpl_5;
  assign mux_50_nl = MUX_s_1_2_2(or_tmp_38, (or_4660_nl), or_2575_cse);
  assign mux_tmp_44 = MUX_s_1_2_2(or_tmp_38, (mux_50_nl), or_309_cse);
  assign mux_52_nl = MUX_s_1_2_2(mux_tmp_2, or_tmp_8, mul_loop_mul_if_land_5_lpi_1_dfm_st_5);
  assign mux_53_nl = MUX_s_1_2_2(mux_tmp_5, or_tmp_9, mul_loop_mul_if_land_5_lpi_1_dfm_st_5);
  assign mux_54_nl = MUX_s_1_2_2((mux_53_nl), (mux_52_nl), or_2575_cse);
  assign mux_tmp_48 = MUX_s_1_2_2(or_tmp_38, (mux_54_nl), or_309_cse);
  assign or_tmp_44 = mul_loop_mul_if_land_6_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign or_tmp_45 = or_tmp_44 | (~ main_stage_v_1);
  assign or_132_nl = mul_loop_mul_if_land_6_lpi_1_dfm_st_5 | mux_tmp_33;
  assign mux_tmp_53 = MUX_s_1_2_2(or_tmp_45, (or_132_nl), or_309_cse);
  assign mux_61_nl = MUX_s_1_2_2(mux_tmp_36, mux_tmp_35, mul_loop_mul_if_land_6_lpi_1_dfm_st_5);
  assign mux_tmp_55 = MUX_s_1_2_2(or_tmp_45, (mux_61_nl), or_309_cse);
  assign or_tmp_50 = mul_loop_mul_if_land_7_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign or_tmp_51 = or_tmp_50 | (~ main_stage_v_1);
  assign or_138_nl = mul_loop_mul_if_land_7_lpi_1_dfm_st_5 | mux_tmp_33;
  assign mux_tmp_60 = MUX_s_1_2_2(or_tmp_51, (or_138_nl), or_309_cse);
  assign mux_68_nl = MUX_s_1_2_2(mux_tmp_36, mux_tmp_35, mul_loop_mul_if_land_7_lpi_1_dfm_st_5);
  assign mux_tmp_62 = MUX_s_1_2_2(or_tmp_51, (mux_68_nl), or_309_cse);
  assign or_tmp_56 = mul_loop_mul_if_land_8_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign or_tmp_57 = or_tmp_56 | (~ main_stage_v_1);
  assign or_4659_nl = mul_loop_mul_if_land_8_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | (~ main_stage_v_1) | and_dcpl_5;
  assign mux_74_nl = MUX_s_1_2_2(or_tmp_57, (or_4659_nl), or_2575_cse);
  assign mux_tmp_68 = MUX_s_1_2_2(or_tmp_57, (mux_74_nl), or_309_cse);
  assign mux_76_nl = MUX_s_1_2_2(mux_tmp_2, or_tmp_8, mul_loop_mul_if_land_8_lpi_1_dfm_st_5);
  assign mux_77_nl = MUX_s_1_2_2(mux_tmp_5, or_tmp_9, mul_loop_mul_if_land_8_lpi_1_dfm_st_5);
  assign mux_78_nl = MUX_s_1_2_2((mux_77_nl), (mux_76_nl), or_2575_cse);
  assign mux_tmp_72 = MUX_s_1_2_2(or_tmp_57, (mux_78_nl), or_309_cse);
  assign or_tmp_63 = mul_loop_mul_if_land_9_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign or_tmp_64 = or_tmp_63 | (~ main_stage_v_1);
  assign or_4658_nl = mul_loop_mul_if_land_9_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | (~ main_stage_v_1) | and_dcpl_5;
  assign mux_84_nl = MUX_s_1_2_2(or_tmp_64, (or_4658_nl), or_2575_cse);
  assign mux_tmp_78 = MUX_s_1_2_2(or_tmp_64, (mux_84_nl), or_309_cse);
  assign mux_86_nl = MUX_s_1_2_2(mux_tmp_2, or_tmp_8, mul_loop_mul_if_land_9_lpi_1_dfm_st_5);
  assign mux_87_nl = MUX_s_1_2_2(mux_tmp_5, or_tmp_9, mul_loop_mul_if_land_9_lpi_1_dfm_st_5);
  assign mux_88_nl = MUX_s_1_2_2((mux_87_nl), (mux_86_nl), or_2575_cse);
  assign mux_tmp_82 = MUX_s_1_2_2(or_tmp_64, (mux_88_nl), or_309_cse);
  assign or_tmp_70 = mul_loop_mul_if_land_10_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign or_tmp_71 = or_tmp_70 | (~ main_stage_v_1);
  assign or_158_nl = mul_loop_mul_if_land_10_lpi_1_dfm_st_5 | mux_tmp_33;
  assign mux_tmp_87 = MUX_s_1_2_2(or_tmp_71, (or_158_nl), or_309_cse);
  assign mux_95_nl = MUX_s_1_2_2(mux_tmp_36, mux_tmp_35, mul_loop_mul_if_land_10_lpi_1_dfm_st_5);
  assign mux_tmp_89 = MUX_s_1_2_2(or_tmp_71, (mux_95_nl), or_309_cse);
  assign or_tmp_76 = mul_loop_mul_if_land_11_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign or_tmp_77 = or_tmp_76 | (~ main_stage_v_1);
  assign or_164_nl = mul_loop_mul_if_land_11_lpi_1_dfm_st_5 | mux_tmp_33;
  assign mux_tmp_94 = MUX_s_1_2_2(or_tmp_77, (or_164_nl), or_309_cse);
  assign mux_102_nl = MUX_s_1_2_2(mux_tmp_36, mux_tmp_35, mul_loop_mul_if_land_11_lpi_1_dfm_st_5);
  assign mux_tmp_96 = MUX_s_1_2_2(or_tmp_77, (mux_102_nl), or_309_cse);
  assign or_tmp_82 = mul_loop_mul_if_land_12_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign or_tmp_83 = or_tmp_82 | (~ main_stage_v_1);
  assign or_170_nl = mul_loop_mul_if_land_12_lpi_1_dfm_st_5 | mux_tmp_33;
  assign mux_tmp_101 = MUX_s_1_2_2(or_tmp_83, (or_170_nl), or_309_cse);
  assign mux_109_nl = MUX_s_1_2_2(mux_tmp_36, mux_tmp_35, mul_loop_mul_if_land_12_lpi_1_dfm_st_5);
  assign mux_tmp_103 = MUX_s_1_2_2(or_tmp_83, (mux_109_nl), or_309_cse);
  assign or_tmp_88 = mul_loop_mul_if_land_13_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign or_tmp_89 = or_tmp_88 | (~ main_stage_v_1);
  assign or_4657_nl = mul_loop_mul_if_land_13_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | (~ main_stage_v_1) | and_dcpl_5;
  assign mux_115_nl = MUX_s_1_2_2(or_tmp_89, (or_4657_nl), or_2575_cse);
  assign mux_tmp_109 = MUX_s_1_2_2(or_tmp_89, (mux_115_nl), or_309_cse);
  assign mux_117_nl = MUX_s_1_2_2(mux_tmp_2, or_tmp_8, mul_loop_mul_if_land_13_lpi_1_dfm_st_5);
  assign mux_118_nl = MUX_s_1_2_2(mux_tmp_5, or_tmp_9, mul_loop_mul_if_land_13_lpi_1_dfm_st_5);
  assign mux_119_nl = MUX_s_1_2_2((mux_118_nl), (mux_117_nl), or_2575_cse);
  assign mux_tmp_113 = MUX_s_1_2_2(or_tmp_89, (mux_119_nl), or_309_cse);
  assign or_tmp_95 = mul_loop_mul_if_land_14_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign or_tmp_96 = or_tmp_95 | (~ main_stage_v_1);
  assign or_183_nl = mul_loop_mul_if_land_14_lpi_1_dfm_st_5 | mux_tmp_33;
  assign mux_tmp_118 = MUX_s_1_2_2(or_tmp_96, (or_183_nl), or_309_cse);
  assign mux_126_nl = MUX_s_1_2_2(mux_tmp_36, mux_tmp_35, mul_loop_mul_if_land_14_lpi_1_dfm_st_5);
  assign mux_tmp_120 = MUX_s_1_2_2(or_tmp_96, (mux_126_nl), or_309_cse);
  assign or_tmp_101 = mul_loop_mul_if_land_15_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign or_tmp_102 = or_tmp_101 | (~ main_stage_v_1);
  assign or_4656_nl = mul_loop_mul_if_land_15_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | (~ main_stage_v_1) | and_dcpl_5;
  assign mux_132_nl = MUX_s_1_2_2(or_tmp_102, (or_4656_nl), or_2575_cse);
  assign mux_tmp_126 = MUX_s_1_2_2(or_tmp_102, (mux_132_nl), or_309_cse);
  assign mux_134_nl = MUX_s_1_2_2(mux_tmp_2, or_tmp_8, mul_loop_mul_if_land_15_lpi_1_dfm_st_5);
  assign mux_135_nl = MUX_s_1_2_2(mux_tmp_5, or_tmp_9, mul_loop_mul_if_land_15_lpi_1_dfm_st_5);
  assign mux_136_nl = MUX_s_1_2_2((mux_135_nl), (mux_134_nl), or_2575_cse);
  assign mux_tmp_130 = MUX_s_1_2_2(or_tmp_102, (mux_136_nl), or_309_cse);
  assign or_tmp_108 = mul_loop_mul_if_land_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign or_tmp_109 = or_tmp_108 | (~ main_stage_v_1);
  assign or_4655_nl = mul_loop_mul_if_land_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | (~ main_stage_v_1) | and_dcpl_5;
  assign mux_142_nl = MUX_s_1_2_2(or_tmp_109, (or_4655_nl), or_2575_cse);
  assign mux_tmp_136 = MUX_s_1_2_2(or_tmp_109, (mux_142_nl), or_309_cse);
  assign mux_144_nl = MUX_s_1_2_2(mux_tmp_2, or_tmp_8, mul_loop_mul_if_land_lpi_1_dfm_st_5);
  assign mux_145_nl = MUX_s_1_2_2(mux_tmp_5, or_tmp_9, mul_loop_mul_if_land_lpi_1_dfm_st_5);
  assign mux_146_nl = MUX_s_1_2_2((mux_145_nl), (mux_144_nl), or_2575_cse);
  assign mux_tmp_140 = MUX_s_1_2_2(or_tmp_109, (mux_146_nl), or_309_cse);
  assign or_tmp_115 = (~ main_stage_v_1) | io_read_cfg_mul_bypass_rsc_svs_st_1 |
      (or_2575_cse & cfg_mul_op_rsc_triosy_obj_bawt & cfg_mul_bypass_rsc_triosy_obj_bawt
      & cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt & or_309_cse);
  assign and_2250_nl = or_4649_cse & main_stage_v_1 & cfg_mul_src_rsc_triosy_obj_bawt
      & cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_bypass_rsc_triosy_obj_bawt &
      cfg_mul_op_rsc_triosy_obj_bawt;
  assign mux_tmp_148 = MUX_s_1_2_2(main_stage_v_2, (and_2250_nl), or_309_cse);
  assign not_tmp_30 = ~(main_stage_v_1 & cfg_mul_src_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_op_rsc_triosy_obj_bawt);
  assign or_tmp_122 = mul_loop_mul_if_land_1_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5;
  assign or_tmp_123 = or_tmp_122 | (~ main_stage_v_2);
  assign or_210_nl = nor_749_cse | mul_loop_mul_if_land_1_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | not_tmp_30;
  assign mux_156_itm = MUX_s_1_2_2(or_tmp_123, (or_210_nl), or_309_cse);
  assign or_tmp_128 = mul_loop_mul_if_land_2_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5;
  assign or_tmp_129 = or_tmp_128 | (~ main_stage_v_2);
  assign or_216_nl = nor_749_cse | mul_loop_mul_if_land_2_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | not_tmp_30;
  assign mux_157_itm = MUX_s_1_2_2(or_tmp_129, (or_216_nl), or_309_cse);
  assign or_tmp_134 = mul_loop_mul_if_land_3_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5;
  assign or_tmp_135 = or_tmp_134 | (~ main_stage_v_2);
  assign or_222_nl = nor_749_cse | mul_loop_mul_if_land_3_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | not_tmp_30;
  assign mux_158_itm = MUX_s_1_2_2(or_tmp_135, (or_222_nl), or_309_cse);
  assign or_tmp_139 = nor_749_cse | io_read_cfg_mul_bypass_rsc_svs_st_1 | not_tmp_30;
  assign or_tmp_141 = mul_loop_mul_if_land_4_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5;
  assign or_tmp_142 = or_tmp_141 | (~ main_stage_v_2);
  assign or_229_nl = mul_loop_mul_if_land_4_lpi_1_dfm_st_5 | or_tmp_139;
  assign mux_159_itm = MUX_s_1_2_2(or_tmp_142, (or_229_nl), or_309_cse);
  assign or_tmp_147 = mul_loop_mul_if_land_5_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5;
  assign or_tmp_148 = or_tmp_147 | (~ main_stage_v_2);
  assign or_235_nl = nor_749_cse | mul_loop_mul_if_land_5_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | not_tmp_30;
  assign mux_160_itm = MUX_s_1_2_2(or_tmp_148, (or_235_nl), or_309_cse);
  assign or_tmp_151 = mul_loop_mul_if_land_6_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5;
  assign or_tmp_152 = or_tmp_151 | (~ main_stage_v_2);
  assign or_239_nl = mul_loop_mul_if_land_6_lpi_1_dfm_st_5 | or_tmp_139;
  assign mux_161_itm = MUX_s_1_2_2(or_tmp_152, (or_239_nl), or_309_cse);
  assign or_tmp_155 = mul_loop_mul_if_land_7_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5;
  assign or_tmp_156 = or_tmp_155 | (~ main_stage_v_2);
  assign or_243_nl = mul_loop_mul_if_land_7_lpi_1_dfm_st_5 | or_tmp_139;
  assign mux_162_itm = MUX_s_1_2_2(or_tmp_156, (or_243_nl), or_309_cse);
  assign or_tmp_161 = mul_loop_mul_if_land_8_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5;
  assign or_tmp_162 = or_tmp_161 | (~ main_stage_v_2);
  assign or_249_nl = nor_749_cse | mul_loop_mul_if_land_8_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | not_tmp_30;
  assign mux_163_itm = MUX_s_1_2_2(or_tmp_162, (or_249_nl), or_309_cse);
  assign or_tmp_167 = mul_loop_mul_if_land_9_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5;
  assign or_tmp_168 = or_tmp_167 | (~ main_stage_v_2);
  assign or_255_nl = nor_749_cse | mul_loop_mul_if_land_9_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | not_tmp_30;
  assign mux_164_itm = MUX_s_1_2_2(or_tmp_168, (or_255_nl), or_309_cse);
  assign or_tmp_171 = mul_loop_mul_if_land_10_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5;
  assign or_tmp_172 = or_tmp_171 | (~ main_stage_v_2);
  assign or_259_nl = mul_loop_mul_if_land_10_lpi_1_dfm_st_5 | or_tmp_139;
  assign mux_165_itm = MUX_s_1_2_2(or_tmp_172, (or_259_nl), or_309_cse);
  assign or_tmp_175 = mul_loop_mul_if_land_11_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5;
  assign or_tmp_176 = or_tmp_175 | (~ main_stage_v_2);
  assign or_263_nl = mul_loop_mul_if_land_11_lpi_1_dfm_st_5 | or_tmp_139;
  assign mux_166_itm = MUX_s_1_2_2(or_tmp_176, (or_263_nl), or_309_cse);
  assign or_tmp_179 = mul_loop_mul_if_land_12_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5;
  assign or_tmp_180 = or_tmp_179 | (~ main_stage_v_2);
  assign or_267_nl = mul_loop_mul_if_land_12_lpi_1_dfm_st_5 | or_tmp_139;
  assign mux_167_itm = MUX_s_1_2_2(or_tmp_180, (or_267_nl), or_309_cse);
  assign or_tmp_185 = mul_loop_mul_if_land_13_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5;
  assign or_tmp_186 = or_tmp_185 | (~ main_stage_v_2);
  assign or_273_nl = nor_749_cse | mul_loop_mul_if_land_13_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | not_tmp_30;
  assign mux_168_itm = MUX_s_1_2_2(or_tmp_186, (or_273_nl), or_309_cse);
  assign or_tmp_189 = mul_loop_mul_if_land_14_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5;
  assign or_tmp_190 = or_tmp_189 | (~ main_stage_v_2);
  assign or_277_nl = mul_loop_mul_if_land_14_lpi_1_dfm_st_5 | or_tmp_139;
  assign mux_169_itm = MUX_s_1_2_2(or_tmp_190, (or_277_nl), or_309_cse);
  assign or_tmp_195 = mul_loop_mul_if_land_15_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5;
  assign or_tmp_196 = or_tmp_195 | (~ main_stage_v_2);
  assign or_283_nl = nor_749_cse | mul_loop_mul_if_land_15_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | not_tmp_30;
  assign mux_170_itm = MUX_s_1_2_2(or_tmp_196, (or_283_nl), or_309_cse);
  assign or_tmp_201 = mul_loop_mul_if_land_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5;
  assign or_tmp_202 = or_tmp_201 | (~ main_stage_v_2);
  assign or_289_nl = nor_749_cse | mul_loop_mul_if_land_lpi_1_dfm_st_5 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | not_tmp_30;
  assign mux_171_itm = MUX_s_1_2_2(or_tmp_202, (or_289_nl), or_309_cse);
  assign or_tmp_204 = io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign nor_50_cse = ~(reg_FpMul_8U_23U_lor_3_lpi_1_dfm_4_cse | (~ mul_loop_mul_1_FpMul_8U_23U_else_2_if_acc_itm_8_1));
  assign or_tmp_213 = IsNaN_8U_23U_land_1_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_6
      | (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_7) | mul_loop_mul_if_land_1_lpi_1_dfm_8
      | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_1_lpi_1_dfm_st_6;
  assign or_tmp_228 = mul_loop_mul_if_land_1_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_187_itm = MUX_s_1_2_2(or_tmp_228, or_tmp_123, or_309_cse);
  assign nor_55_cse = ~(reg_FpMul_8U_23U_lor_4_lpi_1_dfm_4_cse | (~ mul_loop_mul_2_FpMul_8U_23U_else_2_if_acc_itm_8_1));
  assign or_tmp_236 = IsNaN_8U_23U_land_2_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_6
      | (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_7) | mul_loop_mul_if_land_2_lpi_1_dfm_8
      | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_2_lpi_1_dfm_st_6;
  assign or_tmp_248 = FpMul_8U_23U_lor_19_lpi_1_dfm_st_3 | mul_loop_mul_if_land_2_lpi_1_dfm_st_7
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | (~ main_stage_v_3);
  assign or_tmp_256 = mul_loop_mul_if_land_2_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_202_itm = MUX_s_1_2_2(or_tmp_256, or_tmp_129, or_309_cse);
  assign nor_59_cse = ~(reg_FpMul_8U_23U_lor_5_lpi_1_dfm_4_cse | (~ mul_loop_mul_3_FpMul_8U_23U_else_2_if_acc_itm_8_1));
  assign or_tmp_264 = IsNaN_8U_23U_land_3_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_6
      | (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_7) | mul_loop_mul_if_land_3_lpi_1_dfm_8
      | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_3_lpi_1_dfm_st_6;
  assign or_tmp_279 = mul_loop_mul_if_land_3_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_216_itm = MUX_s_1_2_2(or_tmp_279, or_tmp_135, or_309_cse);
  assign nor_64_cse = ~(reg_FpMul_8U_23U_lor_6_lpi_1_dfm_4_cse | (~ mul_loop_mul_4_FpMul_8U_23U_else_2_if_acc_itm_8_1));
  assign or_tmp_287 = IsNaN_8U_23U_land_4_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_6
      | (~ IsNaN_8U_23U_1_land_4_lpi_1_dfm_7) | mul_loop_mul_if_land_4_lpi_1_dfm_8
      | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_4_lpi_1_dfm_st_6;
  assign or_378_cse = (~ mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_21_lpi_1_dfm_st;
  assign or_tmp_302 = mul_loop_mul_if_land_4_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_230_itm = MUX_s_1_2_2(or_tmp_302, or_tmp_142, or_309_cse);
  assign nor_69_cse = ~(reg_FpMul_8U_23U_lor_7_lpi_1_dfm_4_cse | (~ mul_loop_mul_5_FpMul_8U_23U_else_2_if_acc_itm_8_1));
  assign or_tmp_310 = IsNaN_8U_23U_land_5_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_6
      | (~ IsNaN_8U_23U_1_land_5_lpi_1_dfm_7) | mul_loop_mul_if_land_5_lpi_1_dfm_8
      | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_5_lpi_1_dfm_st_6;
  assign or_tmp_321 = FpMul_8U_23U_lor_22_lpi_1_dfm_st_3 | mul_loop_mul_if_land_5_lpi_1_dfm_st_7
      | io_read_cfg_mul_bypass_rsc_svs_st_6;
  assign or_tmp_322 = or_tmp_321 | (~ main_stage_v_3);
  assign or_tmp_331 = mul_loop_mul_if_land_5_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_245_itm = MUX_s_1_2_2(or_tmp_331, or_tmp_148, or_309_cse);
  assign nor_73_cse = ~(reg_FpMul_8U_23U_lor_8_lpi_1_dfm_4_cse | (~ mul_loop_mul_6_FpMul_8U_23U_else_2_if_acc_itm_8_1));
  assign or_tmp_339 = IsNaN_8U_23U_land_6_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_6
      | (~ IsNaN_8U_23U_1_land_6_lpi_1_dfm_7) | mul_loop_mul_if_land_6_lpi_1_dfm_8
      | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_6_lpi_1_dfm_st_6;
  assign or_430_cse = (~ mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_23_lpi_1_dfm_st;
  assign or_tmp_354 = mul_loop_mul_if_land_6_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_259_itm = MUX_s_1_2_2(or_tmp_354, or_tmp_152, or_309_cse);
  assign nor_78_cse = ~(reg_FpMul_8U_23U_lor_9_lpi_1_dfm_4_cse | (~ mul_loop_mul_7_FpMul_8U_23U_else_2_if_acc_itm_8_1));
  assign or_tmp_362 = IsNaN_8U_23U_land_7_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_6
      | (~ IsNaN_8U_23U_1_land_7_lpi_1_dfm_7) | mul_loop_mul_if_land_7_lpi_1_dfm_8
      | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_7_lpi_1_dfm_st_6;
  assign or_453_cse = (~ mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_24_lpi_1_dfm_st;
  assign or_tmp_377 = mul_loop_mul_if_land_7_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_273_itm = MUX_s_1_2_2(or_tmp_377, or_tmp_156, or_309_cse);
  assign nor_83_cse = ~(reg_FpMul_8U_23U_lor_10_lpi_1_dfm_4_cse | (~ mul_loop_mul_8_FpMul_8U_23U_else_2_if_acc_itm_8_1));
  assign or_tmp_385 = IsNaN_8U_23U_land_8_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_6
      | (~ IsNaN_8U_23U_1_land_8_lpi_1_dfm_7) | mul_loop_mul_if_land_8_lpi_1_dfm_8
      | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_8_lpi_1_dfm_st_6;
  assign or_tmp_397 = FpMul_8U_23U_lor_25_lpi_1_dfm_st_3 | mul_loop_mul_if_land_8_lpi_1_dfm_st_7
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | (~ main_stage_v_3);
  assign or_tmp_405 = mul_loop_mul_if_land_8_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_288_itm = MUX_s_1_2_2(or_tmp_405, or_tmp_162, or_309_cse);
  assign nor_87_cse = ~(reg_FpMul_8U_23U_lor_11_lpi_1_dfm_4_cse | (~ mul_loop_mul_9_FpMul_8U_23U_else_2_if_acc_itm_8_1));
  assign or_tmp_413 = IsNaN_8U_23U_land_9_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_6
      | (~ IsNaN_8U_23U_1_land_9_lpi_1_dfm_7) | mul_loop_mul_if_land_9_lpi_1_dfm_8
      | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_9_lpi_1_dfm_st_6;
  assign or_tmp_424 = FpMul_8U_23U_lor_26_lpi_1_dfm_st_3 | mul_loop_mul_if_land_9_lpi_1_dfm_st_7
      | io_read_cfg_mul_bypass_rsc_svs_st_6;
  assign or_tmp_425 = or_tmp_424 | (~ main_stage_v_3);
  assign or_tmp_434 = mul_loop_mul_if_land_9_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_303_itm = MUX_s_1_2_2(or_tmp_434, or_tmp_168, or_309_cse);
  assign nor_91_cse = ~(reg_FpMul_8U_23U_lor_12_lpi_1_dfm_4_cse | (~ mul_loop_mul_10_FpMul_8U_23U_else_2_if_acc_itm_8_1));
  assign or_tmp_442 = IsNaN_8U_23U_land_10_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_6
      | (~ IsNaN_8U_23U_1_land_10_lpi_1_dfm_7) | mul_loop_mul_if_land_10_lpi_1_dfm_8
      | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_10_lpi_1_dfm_st_6;
  assign or_533_cse = (~ mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_27_lpi_1_dfm_st;
  assign or_tmp_453 = FpMul_8U_23U_lor_27_lpi_1_dfm_st_3 | mul_loop_mul_if_land_10_lpi_1_dfm_st_7
      | io_read_cfg_mul_bypass_rsc_svs_st_6;
  assign or_tmp_454 = or_tmp_453 | (~ main_stage_v_3);
  assign or_tmp_460 = reg_FpMul_8U_23U_lor_12_lpi_1_dfm_4_cse | mul_loop_mul_10_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | mul_loop_mul_if_land_10_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign or_tmp_463 = mul_loop_mul_if_land_10_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_318_itm = MUX_s_1_2_2(or_tmp_463, or_tmp_172, or_309_cse);
  assign nor_95_cse = ~(reg_FpMul_8U_23U_lor_13_lpi_1_dfm_4_cse | (~ mul_loop_mul_11_FpMul_8U_23U_else_2_if_acc_itm_8_1));
  assign or_tmp_471 = IsNaN_8U_23U_land_11_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_6
      | (~ IsNaN_8U_23U_1_land_11_lpi_1_dfm_7) | mul_loop_mul_if_land_11_lpi_1_dfm_8
      | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_11_lpi_1_dfm_st_6;
  assign or_562_cse = (~ mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_28_lpi_1_dfm_st;
  assign or_tmp_486 = mul_loop_mul_if_land_11_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_332_itm = MUX_s_1_2_2(or_tmp_486, or_tmp_176, or_309_cse);
  assign nor_100_cse = ~(reg_FpMul_8U_23U_lor_14_lpi_1_dfm_4_cse | (~ mul_loop_mul_12_FpMul_8U_23U_else_2_if_acc_itm_8_1));
  assign or_tmp_494 = IsNaN_8U_23U_land_12_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_6
      | (~ IsNaN_8U_23U_1_land_12_lpi_1_dfm_7) | mul_loop_mul_if_land_12_lpi_1_dfm_8
      | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_12_lpi_1_dfm_st_6;
  assign or_585_cse = (~ mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_29_lpi_1_dfm_st;
  assign or_tmp_509 = mul_loop_mul_if_land_12_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_346_itm = MUX_s_1_2_2(or_tmp_509, or_tmp_180, or_309_cse);
  assign nor_105_cse = ~(reg_FpMul_8U_23U_lor_15_lpi_1_dfm_4_cse | (~ mul_loop_mul_13_FpMul_8U_23U_else_2_if_acc_itm_8_1));
  assign or_tmp_517 = IsNaN_8U_23U_land_13_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_6
      | (~ IsNaN_8U_23U_1_land_13_lpi_1_dfm_7) | mul_loop_mul_if_land_13_lpi_1_dfm_8
      | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_13_lpi_1_dfm_st_6;
  assign or_tmp_532 = mul_loop_mul_if_land_13_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_360_itm = MUX_s_1_2_2(or_tmp_532, or_tmp_186, or_309_cse);
  assign nor_110_cse = ~(reg_FpMul_8U_23U_lor_16_lpi_1_dfm_4_cse | (~ mul_loop_mul_14_FpMul_8U_23U_else_2_if_acc_itm_8_1));
  assign or_tmp_540 = IsNaN_8U_23U_land_14_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_6
      | (~ IsNaN_8U_23U_1_land_14_lpi_1_dfm_7) | mul_loop_mul_if_land_14_lpi_1_dfm_8
      | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_14_lpi_1_dfm_st_6;
  assign or_631_cse = (~ mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st)
      | FpMul_8U_23U_lor_31_lpi_1_dfm_st;
  assign or_tmp_555 = mul_loop_mul_if_land_14_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_374_itm = MUX_s_1_2_2(or_tmp_555, or_tmp_190, or_309_cse);
  assign nor_115_cse = ~(reg_FpMul_8U_23U_lor_17_lpi_1_dfm_4_cse | (~ mul_loop_mul_15_FpMul_8U_23U_else_2_if_acc_itm_8_1));
  assign or_tmp_563 = IsNaN_8U_23U_land_15_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_6
      | (~ IsNaN_8U_23U_1_land_15_lpi_1_dfm_7) | mul_loop_mul_if_land_15_lpi_1_dfm_8
      | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_15_lpi_1_dfm_st_6;
  assign or_tmp_578 = mul_loop_mul_if_land_15_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_388_itm = MUX_s_1_2_2(or_tmp_578, or_tmp_196, or_309_cse);
  assign nor_120_cse = ~(reg_FpMul_8U_23U_lor_lpi_1_dfm_4_cse | (~ mul_loop_mul_16_FpMul_8U_23U_else_2_if_acc_itm_8_1));
  assign or_tmp_586 = IsNaN_8U_23U_land_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_6
      | (~ IsNaN_8U_23U_1_land_lpi_1_dfm_7) | mul_loop_mul_if_land_lpi_1_dfm_8 |
      (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_lpi_1_dfm_st_6;
  assign or_tmp_597 = FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | mul_loop_mul_if_land_lpi_1_dfm_st_7
      | io_read_cfg_mul_bypass_rsc_svs_st_6;
  assign or_tmp_598 = or_tmp_597 | (~ main_stage_v_3);
  assign or_tmp_606 = mul_loop_mul_if_land_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_403_itm = MUX_s_1_2_2(or_tmp_606, or_tmp_202, or_309_cse);
  assign or_tmp_608 = io_read_cfg_mul_bypass_rsc_svs_st_6 | (~ main_stage_v_3);
  assign mux_tmp_399 = mul_loop_mul_if_land_1_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | (~ main_stage_v_3);
  assign mux_tmp_402 = mul_loop_mul_else_land_1_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_tmp_403 = io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_tmp_406 = mul_loop_mul_if_land_2_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | (~ main_stage_v_3);
  assign mux_tmp_409 = mul_loop_mul_else_land_2_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_tmp_412 = mul_loop_mul_if_land_3_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | (~ main_stage_v_3);
  assign mux_tmp_415 = mul_loop_mul_else_land_3_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | (~ main_stage_v_3);
  assign mux_tmp_418 = mul_loop_mul_if_land_4_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | (~ main_stage_v_3);
  assign mux_tmp_421 = mul_loop_mul_else_land_4_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | (~ main_stage_v_3);
  assign mux_tmp_424 = mul_loop_mul_if_land_5_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | (~ main_stage_v_3);
  assign mux_tmp_427 = mul_loop_mul_else_land_5_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | (~ main_stage_v_3);
  assign mux_tmp_430 = mul_loop_mul_if_land_6_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | (~ main_stage_v_3);
  assign mux_tmp_433 = mul_loop_mul_else_land_6_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | (~ main_stage_v_3);
  assign mux_tmp_436 = mul_loop_mul_if_land_7_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | (~ main_stage_v_3);
  assign mux_tmp_439 = mul_loop_mul_else_land_7_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | (~ main_stage_v_3);
  assign mux_tmp_442 = mul_loop_mul_if_land_8_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | (~ main_stage_v_3);
  assign mux_tmp_445 = mul_loop_mul_else_land_8_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | (~ main_stage_v_3);
  assign mux_tmp_448 = mul_loop_mul_if_land_9_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | (~ main_stage_v_3);
  assign mux_tmp_451 = mul_loop_mul_else_land_9_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | (~ main_stage_v_3);
  assign mux_tmp_454 = mul_loop_mul_if_land_10_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | (~ main_stage_v_3);
  assign mux_tmp_457 = mul_loop_mul_else_land_10_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | (~ main_stage_v_3);
  assign mux_tmp_460 = mul_loop_mul_if_land_11_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | (~ main_stage_v_3);
  assign mux_tmp_463 = mul_loop_mul_else_land_11_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_tmp_466 = mul_loop_mul_if_land_12_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | (~ main_stage_v_3);
  assign mux_tmp_469 = mul_loop_mul_else_land_12_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_tmp_472 = mul_loop_mul_if_land_13_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | (~ main_stage_v_3);
  assign mux_tmp_475 = mul_loop_mul_else_land_13_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_tmp_478 = mul_loop_mul_if_land_14_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | (~ main_stage_v_3);
  assign mux_tmp_481 = mul_loop_mul_else_land_14_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_tmp_484 = mul_loop_mul_if_land_15_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | (~ main_stage_v_3);
  assign mux_tmp_487 = mul_loop_mul_else_land_15_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_tmp_490 = mul_loop_mul_if_land_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | (~ main_stage_v_3);
  assign mux_tmp_493 = mul_loop_mul_else_land_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | (~ main_stage_v_3);
  assign or_tmp_893 = FpMul_8U_23U_FpMul_8U_23U_and_itm | FpMul_8U_23U_lor_18_lpi_1_dfm_6;
  assign or_tmp_898 = FpMul_8U_23U_lor_18_lpi_1_dfm_7 | FpMul_8U_23U_FpMul_8U_23U_and_itm_2;
  assign or_tmp_932 = mul_loop_mul_if_land_1_lpi_1_dfm_st_7 | mul_loop_mul_if_land_1_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1044_nl = mul_loop_mul_if_land_1_lpi_1_dfm_st_8 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | (~ main_stage_v_4);
  assign mux_522_itm = MUX_s_1_2_2((or_1044_nl), or_tmp_228, or_309_cse);
  assign or_tmp_958 = IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 | IsNaN_8U_23U_land_1_lpi_1_dfm_10
      | mul_loop_mul_if_land_1_lpi_1_dfm_st_7 | mul_loop_mul_if_land_1_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1049_nl = IsNaN_8U_23U_1_land_1_lpi_1_dfm_9 | IsNaN_8U_23U_land_1_lpi_1_dfm_11
      | mul_loop_mul_if_land_1_lpi_1_dfm_st_8 | mul_loop_mul_if_land_1_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_523_itm = MUX_s_1_2_2((or_1049_nl), or_tmp_958, or_309_cse);
  assign or_tmp_975 = FpMul_8U_23U_FpMul_8U_23U_and_64_itm | FpMul_8U_23U_lor_19_lpi_1_dfm_6;
  assign or_tmp_980 = FpMul_8U_23U_lor_19_lpi_1_dfm_7 | FpMul_8U_23U_FpMul_8U_23U_and_64_itm_2;
  assign or_tmp_1012 = mul_loop_mul_if_land_2_lpi_1_dfm_st_7 | mul_loop_mul_if_land_2_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1124_nl = mul_loop_mul_if_land_2_lpi_1_dfm_st_8 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | (~ main_stage_v_4);
  assign mux_546_itm = MUX_s_1_2_2((or_1124_nl), or_tmp_256, or_309_cse);
  assign or_tmp_1038 = IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 | IsNaN_8U_23U_land_2_lpi_1_dfm_10
      | mul_loop_mul_if_land_2_lpi_1_dfm_st_7 | mul_loop_mul_if_land_2_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1129_nl = IsNaN_8U_23U_1_land_2_lpi_1_dfm_9 | IsNaN_8U_23U_land_2_lpi_1_dfm_11
      | mul_loop_mul_if_land_2_lpi_1_dfm_st_8 | mul_loop_mul_if_land_2_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_547_itm = MUX_s_1_2_2((or_1129_nl), or_tmp_1038, or_309_cse);
  assign or_tmp_1055 = FpMul_8U_23U_FpMul_8U_23U_and_65_itm | FpMul_8U_23U_lor_20_lpi_1_dfm_6;
  assign or_tmp_1060 = FpMul_8U_23U_lor_20_lpi_1_dfm_7 | FpMul_8U_23U_FpMul_8U_23U_and_65_itm_2;
  assign or_tmp_1088 = FpMul_8U_23U_lor_20_lpi_1_dfm_st_3 | mul_loop_mul_if_land_3_lpi_1_dfm_st_7
      | io_read_cfg_mul_bypass_rsc_svs_st_6;
  assign or_tmp_1094 = mul_loop_mul_if_land_3_lpi_1_dfm_st_7 | mul_loop_mul_if_land_3_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1206_nl = mul_loop_mul_if_land_3_lpi_1_dfm_st_8 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | (~ main_stage_v_4);
  assign mux_570_itm = MUX_s_1_2_2((or_1206_nl), or_tmp_279, or_309_cse);
  assign or_tmp_1120 = IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 | IsNaN_8U_23U_land_3_lpi_1_dfm_10
      | mul_loop_mul_if_land_3_lpi_1_dfm_st_7 | mul_loop_mul_if_land_3_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1211_nl = IsNaN_8U_23U_1_land_3_lpi_1_dfm_9 | IsNaN_8U_23U_land_3_lpi_1_dfm_11
      | mul_loop_mul_if_land_3_lpi_1_dfm_st_8 | mul_loop_mul_if_land_3_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_571_itm = MUX_s_1_2_2((or_1211_nl), or_tmp_1120, or_309_cse);
  assign or_tmp_1137 = FpMul_8U_23U_FpMul_8U_23U_and_66_itm | FpMul_8U_23U_lor_21_lpi_1_dfm_6;
  assign or_tmp_1142 = FpMul_8U_23U_lor_21_lpi_1_dfm_7 | FpMul_8U_23U_FpMul_8U_23U_and_66_itm_2;
  assign or_tmp_1177 = mul_loop_mul_if_land_4_lpi_1_dfm_st_7 | mul_loop_mul_if_land_4_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1289_nl = mul_loop_mul_if_land_4_lpi_1_dfm_st_8 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | (~ main_stage_v_4);
  assign mux_596_itm = MUX_s_1_2_2((or_1289_nl), or_tmp_302, or_309_cse);
  assign or_tmp_1203 = IsNaN_8U_23U_land_4_lpi_1_dfm_10 | IsNaN_8U_23U_1_land_4_lpi_1_dfm_8
      | mul_loop_mul_if_land_4_lpi_1_dfm_st_7 | mul_loop_mul_if_land_4_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1294_nl = IsNaN_8U_23U_1_land_4_lpi_1_dfm_9 | IsNaN_8U_23U_land_4_lpi_1_dfm_11
      | mul_loop_mul_if_land_4_lpi_1_dfm_st_8 | mul_loop_mul_if_land_4_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_597_itm = MUX_s_1_2_2((or_1294_nl), or_tmp_1203, or_309_cse);
  assign or_tmp_1220 = FpMul_8U_23U_FpMul_8U_23U_and_67_itm | FpMul_8U_23U_lor_22_lpi_1_dfm_6;
  assign or_tmp_1225 = FpMul_8U_23U_lor_22_lpi_1_dfm_7 | FpMul_8U_23U_FpMul_8U_23U_and_67_itm_2;
  assign or_tmp_1257 = mul_loop_mul_if_land_5_lpi_1_dfm_st_7 | mul_loop_mul_if_land_5_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1369_nl = mul_loop_mul_if_land_5_lpi_1_dfm_st_8 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | (~ main_stage_v_4);
  assign mux_620_itm = MUX_s_1_2_2((or_1369_nl), or_tmp_331, or_309_cse);
  assign or_tmp_1283 = IsNaN_8U_23U_1_land_5_lpi_1_dfm_8 | IsNaN_8U_23U_land_5_lpi_1_dfm_10
      | mul_loop_mul_if_land_5_lpi_1_dfm_st_7 | mul_loop_mul_if_land_5_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1374_nl = IsNaN_8U_23U_land_5_lpi_1_dfm_11 | IsNaN_8U_23U_1_land_5_lpi_1_dfm_9
      | mul_loop_mul_if_land_5_lpi_1_dfm_st_8 | mul_loop_mul_if_land_5_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_621_itm = MUX_s_1_2_2((or_1374_nl), or_tmp_1283, or_309_cse);
  assign or_tmp_1300 = FpMul_8U_23U_FpMul_8U_23U_and_68_itm | FpMul_8U_23U_lor_23_lpi_1_dfm_6;
  assign or_tmp_1305 = FpMul_8U_23U_lor_23_lpi_1_dfm_7 | FpMul_8U_23U_FpMul_8U_23U_and_68_itm_2;
  assign or_tmp_1333 = FpMul_8U_23U_lor_23_lpi_1_dfm_st_3 | mul_loop_mul_if_land_6_lpi_1_dfm_st_7
      | io_read_cfg_mul_bypass_rsc_svs_st_6;
  assign or_tmp_1339 = mul_loop_mul_if_land_6_lpi_1_dfm_st_7 | mul_loop_mul_if_land_6_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1451_nl = mul_loop_mul_if_land_6_lpi_1_dfm_st_8 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | (~ main_stage_v_4);
  assign mux_644_itm = MUX_s_1_2_2((or_1451_nl), or_tmp_354, or_309_cse);
  assign or_tmp_1365 = IsNaN_8U_23U_1_land_6_lpi_1_dfm_8 | IsNaN_8U_23U_land_6_lpi_1_dfm_10
      | mul_loop_mul_if_land_6_lpi_1_dfm_st_7 | mul_loop_mul_if_land_6_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1456_nl = IsNaN_8U_23U_1_land_6_lpi_1_dfm_9 | IsNaN_8U_23U_land_6_lpi_1_dfm_11
      | mul_loop_mul_if_land_6_lpi_1_dfm_st_8 | mul_loop_mul_if_land_6_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_645_itm = MUX_s_1_2_2((or_1456_nl), or_tmp_1365, or_309_cse);
  assign or_tmp_1382 = FpMul_8U_23U_FpMul_8U_23U_and_69_itm | FpMul_8U_23U_lor_24_lpi_1_dfm_6;
  assign or_tmp_1387 = FpMul_8U_23U_lor_24_lpi_1_dfm_7 | FpMul_8U_23U_FpMul_8U_23U_and_69_itm_2;
  assign or_tmp_1415 = FpMul_8U_23U_lor_24_lpi_1_dfm_st_3 | mul_loop_mul_if_land_7_lpi_1_dfm_st_7
      | io_read_cfg_mul_bypass_rsc_svs_st_6;
  assign or_tmp_1421 = mul_loop_mul_if_land_7_lpi_1_dfm_st_7 | mul_loop_mul_if_land_7_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1533_nl = mul_loop_mul_if_land_7_lpi_1_dfm_st_8 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | (~ main_stage_v_4);
  assign mux_668_itm = MUX_s_1_2_2((or_1533_nl), or_tmp_377, or_309_cse);
  assign or_tmp_1447 = IsNaN_8U_23U_1_land_7_lpi_1_dfm_8 | IsNaN_8U_23U_land_7_lpi_1_dfm_10
      | mul_loop_mul_if_land_7_lpi_1_dfm_st_7 | mul_loop_mul_if_land_7_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1538_nl = IsNaN_8U_23U_1_land_7_lpi_1_dfm_9 | IsNaN_8U_23U_land_7_lpi_1_dfm_11
      | mul_loop_mul_if_land_7_lpi_1_dfm_st_8 | mul_loop_mul_if_land_7_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_669_itm = MUX_s_1_2_2((or_1538_nl), or_tmp_1447, or_309_cse);
  assign or_tmp_1464 = FpMul_8U_23U_FpMul_8U_23U_and_70_itm | FpMul_8U_23U_lor_25_lpi_1_dfm_6;
  assign or_tmp_1469 = FpMul_8U_23U_lor_25_lpi_1_dfm_7 | FpMul_8U_23U_FpMul_8U_23U_and_70_itm_2;
  assign or_tmp_1501 = mul_loop_mul_if_land_8_lpi_1_dfm_st_7 | mul_loop_mul_if_land_8_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1613_nl = mul_loop_mul_if_land_8_lpi_1_dfm_st_8 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | (~ main_stage_v_4);
  assign mux_692_itm = MUX_s_1_2_2((or_1613_nl), or_tmp_405, or_309_cse);
  assign or_tmp_1527 = IsNaN_8U_23U_1_land_8_lpi_1_dfm_8 | IsNaN_8U_23U_land_8_lpi_1_dfm_10
      | mul_loop_mul_if_land_8_lpi_1_dfm_st_7 | mul_loop_mul_if_land_8_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1618_nl = IsNaN_8U_23U_1_land_8_lpi_1_dfm_9 | IsNaN_8U_23U_land_8_lpi_1_dfm_11
      | mul_loop_mul_if_land_8_lpi_1_dfm_st_8 | mul_loop_mul_if_land_8_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_693_itm = MUX_s_1_2_2((or_1618_nl), or_tmp_1527, or_309_cse);
  assign or_tmp_1544 = FpMul_8U_23U_FpMul_8U_23U_and_71_itm | FpMul_8U_23U_lor_26_lpi_1_dfm_6;
  assign or_tmp_1549 = FpMul_8U_23U_lor_26_lpi_1_dfm_7 | FpMul_8U_23U_FpMul_8U_23U_and_71_itm_2;
  assign or_tmp_1581 = mul_loop_mul_if_land_9_lpi_1_dfm_st_7 | mul_loop_mul_if_land_9_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1693_nl = mul_loop_mul_if_land_9_lpi_1_dfm_st_8 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | (~ main_stage_v_4);
  assign mux_716_itm = MUX_s_1_2_2((or_1693_nl), or_tmp_434, or_309_cse);
  assign or_tmp_1607 = IsNaN_8U_23U_1_land_9_lpi_1_dfm_8 | IsNaN_8U_23U_land_9_lpi_1_dfm_10
      | mul_loop_mul_if_land_9_lpi_1_dfm_st_7 | mul_loop_mul_if_land_9_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1698_nl = IsNaN_8U_23U_1_land_9_lpi_1_dfm_9 | IsNaN_8U_23U_land_9_lpi_1_dfm_11
      | mul_loop_mul_if_land_9_lpi_1_dfm_st_8 | mul_loop_mul_if_land_9_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_717_itm = MUX_s_1_2_2((or_1698_nl), or_tmp_1607, or_309_cse);
  assign or_tmp_1624 = FpMul_8U_23U_FpMul_8U_23U_and_72_itm | FpMul_8U_23U_lor_27_lpi_1_dfm_6;
  assign or_tmp_1629 = FpMul_8U_23U_lor_27_lpi_1_dfm_7 | FpMul_8U_23U_FpMul_8U_23U_and_72_itm_2;
  assign or_tmp_1661 = mul_loop_mul_if_land_10_lpi_1_dfm_st_7 | mul_loop_mul_if_land_10_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1773_nl = mul_loop_mul_if_land_10_lpi_1_dfm_st_8 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | (~ main_stage_v_4);
  assign mux_740_itm = MUX_s_1_2_2((or_1773_nl), or_tmp_463, or_309_cse);
  assign or_tmp_1687 = IsNaN_8U_23U_land_10_lpi_1_dfm_10 | IsNaN_8U_23U_1_land_10_lpi_1_dfm_8
      | mul_loop_mul_if_land_10_lpi_1_dfm_st_7 | mul_loop_mul_if_land_10_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1778_nl = IsNaN_8U_23U_1_land_10_lpi_1_dfm_9 | IsNaN_8U_23U_land_10_lpi_1_dfm_11
      | mul_loop_mul_if_land_10_lpi_1_dfm_st_8 | mul_loop_mul_if_land_10_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_741_itm = MUX_s_1_2_2((or_1778_nl), or_tmp_1687, or_309_cse);
  assign or_tmp_1703 = FpMul_8U_23U_FpMul_8U_23U_and_73_itm | FpMul_8U_23U_lor_28_lpi_1_dfm_6;
  assign or_tmp_1709 = FpMul_8U_23U_lor_28_lpi_1_dfm_7 | FpMul_8U_23U_FpMul_8U_23U_and_73_itm_2;
  assign or_tmp_1736 = nor_872_cse | mul_loop_mul_if_land_11_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign or_1828_nl = mul_loop_mul_if_land_11_lpi_1_dfm_st_8 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | (~ main_stage_v_4);
  assign mux_tmp_748 = MUX_s_1_2_2((or_1828_nl), or_tmp_486, or_309_cse);
  assign or_tmp_1744 = mul_loop_mul_if_land_11_lpi_1_dfm_st_7 | mul_loop_mul_if_land_11_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_tmp_1765 = IsNaN_8U_23U_1_land_11_lpi_1_dfm_8 | IsNaN_8U_23U_land_11_lpi_1_dfm_10
      | mul_loop_mul_if_land_11_lpi_1_dfm_st_7 | mul_loop_mul_if_land_11_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1856_nl = IsNaN_8U_23U_1_land_11_lpi_1_dfm_9 | IsNaN_8U_23U_land_11_lpi_1_dfm_11
      | mul_loop_mul_if_land_11_lpi_1_dfm_st_8 | mul_loop_mul_if_land_11_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_767_itm = MUX_s_1_2_2((or_1856_nl), or_tmp_1765, or_309_cse);
  assign or_tmp_1782 = FpMul_8U_23U_FpMul_8U_23U_and_74_itm | FpMul_8U_23U_lor_29_lpi_1_dfm_6;
  assign or_tmp_1786 = FpMul_8U_23U_lor_29_lpi_1_dfm_7 | FpMul_8U_23U_FpMul_8U_23U_and_74_itm_2;
  assign or_tmp_1822 = mul_loop_mul_if_land_12_lpi_1_dfm_st_7 | mul_loop_mul_if_land_12_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1934_nl = mul_loop_mul_if_land_12_lpi_1_dfm_st_8 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | (~ main_stage_v_4);
  assign mux_793_itm = MUX_s_1_2_2((or_1934_nl), or_tmp_509, or_309_cse);
  assign or_tmp_1848 = IsNaN_8U_23U_1_land_12_lpi_1_dfm_8 | IsNaN_8U_23U_land_12_lpi_1_dfm_10
      | mul_loop_mul_if_land_12_lpi_1_dfm_st_7 | mul_loop_mul_if_land_12_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_1939_nl = IsNaN_8U_23U_1_land_12_lpi_1_dfm_9 | IsNaN_8U_23U_land_12_lpi_1_dfm_11
      | mul_loop_mul_if_land_12_lpi_1_dfm_st_8 | mul_loop_mul_if_land_12_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_794_itm = MUX_s_1_2_2((or_1939_nl), or_tmp_1848, or_309_cse);
  assign or_tmp_1865 = FpMul_8U_23U_FpMul_8U_23U_and_75_itm | FpMul_8U_23U_lor_30_lpi_1_dfm_6;
  assign or_tmp_1869 = FpMul_8U_23U_lor_30_lpi_1_dfm_7 | FpMul_8U_23U_FpMul_8U_23U_and_75_itm_2;
  assign or_tmp_1905 = mul_loop_mul_if_land_13_lpi_1_dfm_st_7 | mul_loop_mul_if_land_13_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_2017_nl = mul_loop_mul_if_land_13_lpi_1_dfm_st_8 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | (~ main_stage_v_4);
  assign mux_820_itm = MUX_s_1_2_2((or_2017_nl), or_tmp_532, or_309_cse);
  assign or_tmp_1931 = IsNaN_8U_23U_1_land_13_lpi_1_dfm_8 | IsNaN_8U_23U_land_13_lpi_1_dfm_10
      | mul_loop_mul_if_land_13_lpi_1_dfm_st_7 | mul_loop_mul_if_land_13_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_2022_nl = IsNaN_8U_23U_1_land_13_lpi_1_dfm_9 | IsNaN_8U_23U_land_13_lpi_1_dfm_11
      | mul_loop_mul_if_land_13_lpi_1_dfm_st_8 | mul_loop_mul_if_land_13_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_821_itm = MUX_s_1_2_2((or_2022_nl), or_tmp_1931, or_309_cse);
  assign or_tmp_1947 = FpMul_8U_23U_FpMul_8U_23U_and_76_itm | FpMul_8U_23U_lor_31_lpi_1_dfm_6;
  assign or_tmp_1957 = FpMul_8U_23U_FpMul_8U_23U_and_76_itm_2 | FpMul_8U_23U_lor_31_lpi_1_dfm_7;
  assign or_tmp_1985 = FpMul_8U_23U_lor_31_lpi_1_dfm_st_3 | mul_loop_mul_if_land_14_lpi_1_dfm_st_7
      | io_read_cfg_mul_bypass_rsc_svs_st_6;
  assign or_tmp_1991 = mul_loop_mul_if_land_14_lpi_1_dfm_st_7 | mul_loop_mul_if_land_14_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_2101_nl = mul_loop_mul_if_land_14_lpi_1_dfm_st_8 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | (~ main_stage_v_4);
  assign mux_845_itm = MUX_s_1_2_2((or_2101_nl), or_tmp_555, or_309_cse);
  assign or_tmp_2015 = IsNaN_8U_23U_1_land_14_lpi_1_dfm_8 | IsNaN_8U_23U_land_14_lpi_1_dfm_10
      | mul_loop_mul_if_land_14_lpi_1_dfm_st_7 | mul_loop_mul_if_land_14_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_2106_nl = IsNaN_8U_23U_1_land_14_lpi_1_dfm_9 | IsNaN_8U_23U_land_14_lpi_1_dfm_11
      | mul_loop_mul_if_land_14_lpi_1_dfm_st_8 | mul_loop_mul_if_land_14_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_846_itm = MUX_s_1_2_2((or_2106_nl), or_tmp_2015, or_309_cse);
  assign or_tmp_2032 = FpMul_8U_23U_FpMul_8U_23U_and_77_itm | FpMul_8U_23U_lor_32_lpi_1_dfm_6;
  assign or_tmp_2036 = FpMul_8U_23U_lor_32_lpi_1_dfm_7 | FpMul_8U_23U_FpMul_8U_23U_and_77_itm_2;
  assign or_tmp_2065 = FpMul_8U_23U_lor_32_lpi_1_dfm_st_3 | mul_loop_mul_if_land_15_lpi_1_dfm_st_7
      | io_read_cfg_mul_bypass_rsc_svs_st_6;
  assign or_tmp_2071 = mul_loop_mul_if_land_15_lpi_1_dfm_st_7 | mul_loop_mul_if_land_15_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_2183_nl = mul_loop_mul_if_land_15_lpi_1_dfm_st_8 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | (~ main_stage_v_4);
  assign mux_870_itm = MUX_s_1_2_2((or_2183_nl), or_tmp_578, or_309_cse);
  assign or_tmp_2097 = IsNaN_8U_23U_1_land_15_lpi_1_dfm_8 | IsNaN_8U_23U_land_15_lpi_1_dfm_10
      | mul_loop_mul_if_land_15_lpi_1_dfm_st_7 | mul_loop_mul_if_land_15_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_2188_nl = IsNaN_8U_23U_1_land_15_lpi_1_dfm_9 | IsNaN_8U_23U_land_15_lpi_1_dfm_11
      | mul_loop_mul_if_land_15_lpi_1_dfm_st_8 | mul_loop_mul_if_land_15_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_871_itm = MUX_s_1_2_2((or_2188_nl), or_tmp_2097, or_309_cse);
  assign or_tmp_2114 = FpMul_8U_23U_FpMul_8U_23U_and_78_itm | FpMul_8U_23U_lor_1_lpi_1_dfm_6;
  assign or_tmp_2118 = FpMul_8U_23U_lor_1_lpi_1_dfm_7 | FpMul_8U_23U_FpMul_8U_23U_and_78_itm_2;
  assign or_tmp_2151 = mul_loop_mul_if_land_lpi_1_dfm_st_7 | mul_loop_mul_if_land_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_2263_nl = mul_loop_mul_if_land_lpi_1_dfm_st_8 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | (~ main_stage_v_4);
  assign mux_895_itm = MUX_s_1_2_2((or_2263_nl), or_tmp_606, or_309_cse);
  assign or_tmp_2177 = IsNaN_8U_23U_1_land_lpi_1_dfm_8 | IsNaN_8U_23U_land_lpi_1_dfm_10
      | mul_loop_mul_if_land_lpi_1_dfm_st_7 | mul_loop_mul_if_land_lpi_1_dfm_9 |
      io_read_cfg_mul_bypass_rsc_svs_7 | io_read_cfg_mul_bypass_rsc_svs_st_6 | (~
      main_stage_v_3);
  assign or_2268_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_9 | IsNaN_8U_23U_land_lpi_1_dfm_11
      | mul_loop_mul_if_land_lpi_1_dfm_st_8 | mul_loop_mul_if_land_lpi_1_dfm_10 |
      io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~
      main_stage_v_4);
  assign mux_896_itm = MUX_s_1_2_2((or_2268_nl), or_tmp_2177, or_309_cse);
  assign or_tmp_2227 = nor_872_cse | mul_loop_mul_if_land_4_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign or_tmp_2254 = FpMul_8U_23U_FpMul_8U_23U_and_68_itm | (~ or_tmp_354);
  assign and_tmp_72 = FpMul_8U_23U_FpMul_8U_23U_and_68_itm & or_tmp_354;
  assign or_tmp_2298 = FpMul_8U_23U_FpMul_8U_23U_and_72_itm | (~ or_tmp_463);
  assign and_tmp_76 = FpMul_8U_23U_FpMul_8U_23U_and_72_itm & or_tmp_463;
  assign or_tmp_2310 = nor_872_cse | mul_loop_mul_if_land_12_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign or_tmp_2319 = nor_872_cse | mul_loop_mul_if_land_13_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign or_tmp_2358 = IsNaN_8U_23U_land_1_lpi_1_dfm_st_6 | IsNaN_8U_23U_land_1_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_6 | (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_7)
      | mul_loop_mul_if_land_1_lpi_1_dfm_8 | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_1_lpi_1_dfm_st_6;
  assign or_tmp_2366 = IsNaN_8U_23U_land_2_lpi_1_dfm_st_6 | IsNaN_8U_23U_land_2_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_6 | (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_7)
      | mul_loop_mul_if_land_2_lpi_1_dfm_8 | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_2_lpi_1_dfm_st_6;
  assign or_tmp_2376 = io_read_cfg_mul_bypass_rsc_svs_6 | (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_7)
      | mul_loop_mul_if_land_3_lpi_1_dfm_8 | (~ main_stage_v_2);
  assign or_tmp_2384 = io_read_cfg_mul_bypass_rsc_svs_6 | (~ IsNaN_8U_23U_1_land_4_lpi_1_dfm_7)
      | mul_loop_mul_if_land_4_lpi_1_dfm_8 | (~ main_stage_v_2);
  assign or_tmp_2392 = io_read_cfg_mul_bypass_rsc_svs_6 | (~ IsNaN_8U_23U_1_land_5_lpi_1_dfm_7)
      | mul_loop_mul_if_land_5_lpi_1_dfm_8 | (~ main_stage_v_2);
  assign or_tmp_2400 = io_read_cfg_mul_bypass_rsc_svs_6 | (~ IsNaN_8U_23U_1_land_6_lpi_1_dfm_7)
      | mul_loop_mul_if_land_6_lpi_1_dfm_8 | (~ main_stage_v_2);
  assign or_tmp_2408 = io_read_cfg_mul_bypass_rsc_svs_6 | (~ IsNaN_8U_23U_1_land_7_lpi_1_dfm_7)
      | mul_loop_mul_if_land_7_lpi_1_dfm_8 | (~ main_stage_v_2);
  assign or_tmp_2414 = IsNaN_8U_23U_land_8_lpi_1_dfm_st_6 | IsNaN_8U_23U_land_8_lpi_1_dfm_9
      | io_read_cfg_mul_bypass_rsc_svs_6 | (~ IsNaN_8U_23U_1_land_8_lpi_1_dfm_7)
      | mul_loop_mul_if_land_8_lpi_1_dfm_8 | (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_8_lpi_1_dfm_st_6;
  assign or_tmp_2424 = io_read_cfg_mul_bypass_rsc_svs_6 | (~ IsNaN_8U_23U_1_land_9_lpi_1_dfm_7)
      | mul_loop_mul_if_land_9_lpi_1_dfm_8 | (~ main_stage_v_2);
  assign or_tmp_2432 = io_read_cfg_mul_bypass_rsc_svs_6 | (~ IsNaN_8U_23U_1_land_10_lpi_1_dfm_7)
      | mul_loop_mul_if_land_10_lpi_1_dfm_8 | (~ main_stage_v_2);
  assign or_tmp_2440 = io_read_cfg_mul_bypass_rsc_svs_6 | (~ IsNaN_8U_23U_1_land_11_lpi_1_dfm_7)
      | mul_loop_mul_if_land_11_lpi_1_dfm_8 | (~ main_stage_v_2);
  assign or_tmp_2448 = io_read_cfg_mul_bypass_rsc_svs_6 | (~ IsNaN_8U_23U_1_land_12_lpi_1_dfm_7)
      | mul_loop_mul_if_land_12_lpi_1_dfm_8 | (~ main_stage_v_2);
  assign or_tmp_2456 = io_read_cfg_mul_bypass_rsc_svs_6 | (~ IsNaN_8U_23U_1_land_13_lpi_1_dfm_7)
      | mul_loop_mul_if_land_13_lpi_1_dfm_8 | (~ main_stage_v_2);
  assign or_tmp_2464 = io_read_cfg_mul_bypass_rsc_svs_6 | (~ IsNaN_8U_23U_1_land_14_lpi_1_dfm_7)
      | mul_loop_mul_if_land_14_lpi_1_dfm_8 | (~ main_stage_v_2);
  assign or_tmp_2472 = io_read_cfg_mul_bypass_rsc_svs_6 | (~ IsNaN_8U_23U_1_land_15_lpi_1_dfm_7)
      | mul_loop_mul_if_land_15_lpi_1_dfm_8 | (~ main_stage_v_2);
  assign or_tmp_2480 = io_read_cfg_mul_bypass_rsc_svs_6 | (~ IsNaN_8U_23U_1_land_lpi_1_dfm_7)
      | mul_loop_mul_if_land_lpi_1_dfm_8 | (~ main_stage_v_2);
  assign or_tmp_2490 = FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_tmp | (~ or_309_cse);
  assign or_tmp_2492 = FpMul_8U_23U_lor_3_lpi_1_dfm_st | (~ or_309_cse);
  assign and_tmp_86 = FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_tmp & or_309_cse;
  assign or_2591_nl = reg_FpMul_8U_23U_lor_3_lpi_1_dfm_4_cse | (~ reg_chn_mul_out_rsci_ld_core_psct_cse)
      | chn_mul_out_rsci_bawt;
  assign mux_1138_nl = MUX_s_1_2_2(or_309_cse, (or_2591_nl), or_2577_cse);
  assign or_tmp_2503 = (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 |
      mul_loop_mul_if_land_1_lpi_1_dfm_st_6 | (mux_1138_nl);
  assign or_tmp_2521 = FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_2_tmp | (~ or_309_cse);
  assign or_tmp_2523 = FpMul_8U_23U_lor_4_lpi_1_dfm_st | (~ or_309_cse);
  assign and_tmp_90 = FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_2_tmp & or_309_cse;
  assign or_2622_nl = reg_FpMul_8U_23U_lor_4_lpi_1_dfm_4_cse | (~ reg_chn_mul_out_rsci_ld_core_psct_cse)
      | chn_mul_out_rsci_bawt;
  assign mux_1160_nl = MUX_s_1_2_2(or_309_cse, (or_2622_nl), or_2608_cse);
  assign or_tmp_2534 = (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 |
      mul_loop_mul_if_land_2_lpi_1_dfm_st_6 | (mux_1160_nl);
  assign or_tmp_2538 = FpMul_8U_23U_lor_19_lpi_1_dfm_st | (~ or_tmp_129);
  assign or_tmp_2544 = FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_4_tmp | (~ or_309_cse);
  assign or_tmp_2546 = FpMul_8U_23U_lor_5_lpi_1_dfm_st | (~ or_309_cse);
  assign and_tmp_95 = FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_4_tmp & or_309_cse;
  assign or_2645_nl = reg_FpMul_8U_23U_lor_5_lpi_1_dfm_4_cse | (~ reg_chn_mul_out_rsci_ld_core_psct_cse)
      | chn_mul_out_rsci_bawt;
  assign mux_1183_nl = MUX_s_1_2_2(or_309_cse, (or_2645_nl), or_2631_cse);
  assign or_tmp_2557 = (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 |
      mul_loop_mul_if_land_3_lpi_1_dfm_st_6 | (mux_1183_nl);
  assign or_tmp_2588 = FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_8_tmp | (~ or_309_cse);
  assign or_tmp_2590 = FpMul_8U_23U_lor_7_lpi_1_dfm_st | (~ or_309_cse);
  assign and_tmp_99 = FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_8_tmp & or_309_cse;
  assign or_2689_nl = reg_FpMul_8U_23U_lor_7_lpi_1_dfm_4_cse | (~ reg_chn_mul_out_rsci_ld_core_psct_cse)
      | chn_mul_out_rsci_bawt;
  assign mux_1210_nl = MUX_s_1_2_2(or_309_cse, (or_2689_nl), or_2675_cse);
  assign or_tmp_2601 = (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 |
      mul_loop_mul_if_land_5_lpi_1_dfm_st_6 | (mux_1210_nl);
  assign or_tmp_2604 = FpMul_8U_23U_lor_22_lpi_1_dfm_st | (~ or_tmp_148);
  assign or_tmp_2635 = FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_14_tmp | (~ or_309_cse);
  assign or_tmp_2637 = FpMul_8U_23U_lor_10_lpi_1_dfm_st | (~ or_309_cse);
  assign and_tmp_104 = FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_14_tmp & or_309_cse;
  assign or_2736_nl = reg_FpMul_8U_23U_lor_10_lpi_1_dfm_4_cse | (~ reg_chn_mul_out_rsci_ld_core_psct_cse)
      | chn_mul_out_rsci_bawt;
  assign mux_1244_nl = MUX_s_1_2_2(or_309_cse, (or_2736_nl), or_2722_cse);
  assign or_tmp_2648 = (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 |
      mul_loop_mul_if_land_8_lpi_1_dfm_st_6 | (mux_1244_nl);
  assign or_tmp_2652 = FpMul_8U_23U_lor_25_lpi_1_dfm_st | (~ or_tmp_162);
  assign or_tmp_2658 = FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_16_tmp | (~ or_309_cse);
  assign or_tmp_2660 = FpMul_8U_23U_lor_11_lpi_1_dfm_st | (~ or_309_cse);
  assign and_tmp_109 = FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_16_tmp & or_309_cse;
  assign or_2759_nl = reg_FpMul_8U_23U_lor_11_lpi_1_dfm_4_cse | (~ reg_chn_mul_out_rsci_ld_core_psct_cse)
      | chn_mul_out_rsci_bawt;
  assign mux_1267_nl = MUX_s_1_2_2(or_309_cse, (or_2759_nl), or_2745_cse);
  assign or_tmp_2671 = (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 |
      mul_loop_mul_if_land_9_lpi_1_dfm_st_6 | (mux_1267_nl);
  assign or_tmp_2674 = FpMul_8U_23U_lor_26_lpi_1_dfm_st | (~ or_tmp_168);
  assign or_tmp_2711 = FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_24_tmp | (~ or_309_cse);
  assign or_tmp_2713 = FpMul_8U_23U_lor_15_lpi_1_dfm_st | (~ or_309_cse);
  assign and_tmp_114 = FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_24_tmp & or_309_cse;
  assign or_2812_nl = reg_FpMul_8U_23U_lor_15_lpi_1_dfm_4_cse | (~ reg_chn_mul_out_rsci_ld_core_psct_cse)
      | chn_mul_out_rsci_bawt;
  assign mux_1306_nl = MUX_s_1_2_2(or_309_cse, (or_2812_nl), or_2798_cse);
  assign or_tmp_2724 = (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 |
      mul_loop_mul_if_land_13_lpi_1_dfm_st_6 | (mux_1306_nl);
  assign or_tmp_2728 = FpMul_8U_23U_lor_30_lpi_1_dfm_st | (~ or_tmp_186);
  assign or_tmp_2747 = FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_28_tmp | (~ or_309_cse);
  assign or_tmp_2749 = FpMul_8U_23U_lor_17_lpi_1_dfm_st | (~ or_309_cse);
  assign and_tmp_119 = FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_28_tmp & or_309_cse;
  assign or_2848_nl = reg_FpMul_8U_23U_lor_17_lpi_1_dfm_4_cse | (~ reg_chn_mul_out_rsci_ld_core_psct_cse)
      | chn_mul_out_rsci_bawt;
  assign mux_1334_nl = MUX_s_1_2_2(or_309_cse, (or_2848_nl), or_2834_cse);
  assign or_tmp_2760 = (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 |
      mul_loop_mul_if_land_15_lpi_1_dfm_st_6 | (mux_1334_nl);
  assign or_tmp_2778 = FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_30_tmp | (~ or_309_cse);
  assign or_tmp_2780 = FpMul_8U_23U_lor_lpi_1_dfm_st | (~ or_309_cse);
  assign and_tmp_123 = FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_30_tmp & or_309_cse;
  assign or_2879_nl = reg_FpMul_8U_23U_lor_lpi_1_dfm_4_cse | (~ reg_chn_mul_out_rsci_ld_core_psct_cse)
      | chn_mul_out_rsci_bawt;
  assign mux_1356_nl = MUX_s_1_2_2(or_309_cse, (or_2879_nl), or_2865_cse);
  assign or_tmp_2791 = (~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5 |
      mul_loop_mul_if_land_lpi_1_dfm_st_6 | (mux_1356_nl);
  assign or_tmp_2795 = FpMul_8U_23U_lor_1_lpi_1_dfm_st | (~ or_tmp_202);
  assign or_2950_nl = (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt
      | main_stage_v_1;
  assign mux_1428_nl = MUX_s_1_2_2(main_stage_v_1, (~ or_dcpl_4), or_309_cse);
  assign mux_tmp_1422 = MUX_s_1_2_2((mux_1428_nl), (or_2950_nl), chn_mul_in_rsci_bawt);
  assign not_tmp_845 = ~(main_stage_v_2 | (~ or_2577_cse));
  assign or_2958_nl = nor_821_cse | FpMul_8U_23U_lor_18_lpi_1_dfm_st | (~ mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st);
  assign mux_1431_nl = MUX_s_1_2_2(not_tmp_845, or_2577_cse, or_tmp_122);
  assign or_2961_nl = mul_loop_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1 | (~ mul_loop_mul_1_FpMul_8U_23U_else_2_if_acc_itm_8_1)
      | reg_FpMul_8U_23U_lor_3_lpi_1_dfm_4_cse;
  assign mux_tmp_1427 = MUX_s_1_2_2((mux_1431_nl), (or_2958_nl), or_2961_nl);
  assign mux_tmp_1430 = mux_tmp_1427 & FpMul_8U_23U_lor_3_lpi_1_dfm_st;
  assign or_tmp_2894 = mul_loop_mul_if_land_15_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_6;
  assign or_tmp_2905 = mul_loop_mul_if_land_14_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_6;
  assign or_tmp_2916 = mul_loop_mul_if_land_13_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_6;
  assign or_tmp_2927 = mul_loop_mul_if_land_12_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_6;
  assign or_tmp_2938 = mul_loop_mul_if_land_11_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_6;
  assign or_tmp_2949 = mul_loop_mul_if_land_10_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_6;
  assign or_tmp_2960 = mul_loop_mul_if_land_9_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_6;
  assign or_tmp_2971 = mul_loop_mul_if_land_8_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_6;
  assign or_tmp_2982 = mul_loop_mul_if_land_7_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_6;
  assign or_tmp_2993 = mul_loop_mul_if_land_6_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_6;
  assign or_tmp_3004 = mul_loop_mul_if_land_5_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_6;
  assign or_tmp_3015 = mul_loop_mul_if_land_4_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_6;
  assign or_tmp_3026 = mul_loop_mul_if_land_3_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_6;
  assign or_tmp_3037 = mul_loop_mul_if_land_2_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_6;
  assign or_tmp_3048 = mul_loop_mul_if_land_1_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_6;
  assign mux_tmp_1504 = mul_loop_mul_else_land_15_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | io_read_cfg_mul_bypass_rsc_svs_6 | (~ main_stage_v_2);
  assign mux_tmp_1507 = mul_loop_mul_else_land_14_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | io_read_cfg_mul_bypass_rsc_svs_6 | (~ main_stage_v_2);
  assign mux_tmp_1510 = mul_loop_mul_else_land_13_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | io_read_cfg_mul_bypass_rsc_svs_6 | (~ main_stage_v_2);
  assign mux_tmp_1513 = mul_loop_mul_else_land_12_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | io_read_cfg_mul_bypass_rsc_svs_6 | (~ main_stage_v_2);
  assign mux_tmp_1516 = mul_loop_mul_else_land_11_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | io_read_cfg_mul_bypass_rsc_svs_6 | (~ main_stage_v_2);
  assign mux_tmp_1535 = mul_loop_mul_else_land_2_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | io_read_cfg_mul_bypass_rsc_svs_6 | (~ main_stage_v_2);
  assign mux_tmp_1538 = mul_loop_mul_else_land_1_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | io_read_cfg_mul_bypass_rsc_svs_6 | (~ main_stage_v_2);
  assign and_dcpl_47 = chn_mul_out_rsci_bawt & reg_chn_mul_out_rsci_ld_core_psct_cse;
  assign and_dcpl_50 = (~ chn_mul_out_rsci_bawt) & reg_chn_mul_out_rsci_ld_core_psct_cse;
  assign and_dcpl_52 = (~ io_read_cfg_mul_bypass_rsc_svs_st_1) & (~ chn_mul_op_rsci_bawt)
      & cfg_mul_src_1_sva_st_1;
  assign or_dcpl_27 = (~(cfg_mul_op_rsc_triosy_obj_bawt & cfg_mul_bypass_rsc_triosy_obj_bawt))
      | (~(cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt));
  assign and_dcpl_53 = (or_dcpl_27 | and_dcpl_52) & main_stage_v_1;
  assign and_dcpl_56 = or_309_cse & main_stage_v_4;
  assign and_dcpl_58 = (~ main_stage_v_4) & chn_mul_out_rsci_bawt & reg_chn_mul_out_rsci_ld_core_psct_cse;
  assign and_dcpl_59 = (~ cfg_mul_bypass_rsci_d) & chn_mul_in_rsci_bawt;
  assign or_dcpl_31 = cfg_mul_bypass_rsci_d | (~ chn_mul_in_rsci_bawt);
  assign and_dcpl_67 = (~ io_read_cfg_mul_bypass_rsc_svs_st_1) & chn_mul_op_rsci_bawt
      & cfg_mul_src_1_sva_st_1;
  assign nor_tmp_568 = main_stage_v_1 & cfg_mul_src_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_op_rsc_triosy_obj_bawt;
  assign and_dcpl_72 = and_dcpl_3 & main_stage_v_1;
  assign and_dcpl_75 = or_4649_cse & and_dcpl_4 & and_dcpl_72 & or_309_cse;
  assign and_dcpl_85 = (cfg_precision==2'b10);
  assign and_dcpl_87 = and_dcpl_7 & or_90_cse;
  assign or_dcpl_46 = and_dcpl_53 | and_dcpl_50;
  assign and_dcpl_91 = cfg_mul_bypass_rsci_d & chn_mul_in_rsci_bawt;
  assign and_dcpl_95 = or_309_cse & main_stage_v_2;
  assign and_dcpl_100 = or_309_cse & (~ io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign and_dcpl_102 = (or_tmp_4 | or_90_cse) & or_309_cse;
  assign and_dcpl_104 = or_309_cse & or_90_cse;
  assign and_dcpl_108 = (or_tmp_14 | or_90_cse) & or_309_cse;
  assign and_dcpl_112 = (or_tmp_21 | or_90_cse) & or_309_cse;
  assign and_dcpl_116 = (or_tmp_29 | or_90_cse) & or_309_cse;
  assign and_dcpl_120 = (or_tmp_37 | or_90_cse) & or_309_cse;
  assign and_dcpl_124 = (or_tmp_44 | or_90_cse) & or_309_cse;
  assign and_dcpl_128 = (or_tmp_50 | or_90_cse) & or_309_cse;
  assign and_dcpl_132 = (or_tmp_56 | or_90_cse) & or_309_cse;
  assign and_dcpl_136 = (or_tmp_63 | or_90_cse) & or_309_cse;
  assign and_dcpl_140 = (or_tmp_70 | or_90_cse) & or_309_cse;
  assign and_dcpl_144 = (or_tmp_76 | or_90_cse) & or_309_cse;
  assign and_dcpl_148 = (or_tmp_82 | or_90_cse) & or_309_cse;
  assign and_dcpl_152 = (or_tmp_88 | or_90_cse) & or_309_cse;
  assign and_dcpl_156 = (or_tmp_95 | or_90_cse) & or_309_cse;
  assign and_dcpl_160 = (or_tmp_101 | or_90_cse) & or_309_cse;
  assign and_dcpl_164 = (or_tmp_108 | or_90_cse) & or_309_cse;
  assign and_dcpl_172 = or_309_cse & (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_8);
  assign and_dcpl_177 = or_309_cse & (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_8);
  assign and_dcpl_182 = or_309_cse & (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_8);
  assign and_dcpl_187 = or_309_cse & (~ IsNaN_8U_23U_1_land_4_lpi_1_dfm_8);
  assign and_dcpl_192 = or_309_cse & (~ IsNaN_8U_23U_1_land_5_lpi_1_dfm_8);
  assign and_dcpl_197 = or_309_cse & (~ IsNaN_8U_23U_1_land_6_lpi_1_dfm_8);
  assign and_dcpl_202 = or_309_cse & (~ IsNaN_8U_23U_1_land_7_lpi_1_dfm_8);
  assign and_dcpl_207 = or_309_cse & (~ IsNaN_8U_23U_1_land_8_lpi_1_dfm_8);
  assign and_dcpl_212 = or_309_cse & (~ IsNaN_8U_23U_1_land_9_lpi_1_dfm_8);
  assign and_dcpl_217 = or_309_cse & (~ IsNaN_8U_23U_1_land_10_lpi_1_dfm_8);
  assign and_dcpl_222 = or_309_cse & (~ IsNaN_8U_23U_1_land_11_lpi_1_dfm_8);
  assign and_dcpl_227 = or_309_cse & (~ IsNaN_8U_23U_1_land_12_lpi_1_dfm_8);
  assign and_dcpl_232 = or_309_cse & (~ IsNaN_8U_23U_1_land_13_lpi_1_dfm_8);
  assign and_dcpl_237 = or_309_cse & (~ IsNaN_8U_23U_1_land_14_lpi_1_dfm_8);
  assign and_dcpl_242 = or_309_cse & (~ IsNaN_8U_23U_1_land_15_lpi_1_dfm_8);
  assign and_dcpl_247 = or_309_cse & (~ IsNaN_8U_23U_1_land_lpi_1_dfm_8);
  assign or_dcpl_87 = and_dcpl_50 | or_90_cse;
  assign or_dcpl_92 = or_tmp_608 | mul_loop_mul_if_land_1_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_18_lpi_1_dfm_st_3
      | (~ mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | or_dcpl_87;
  assign or_dcpl_95 = or_tmp_608 | and_dcpl_50;
  assign or_dcpl_96 = or_dcpl_95 | mul_loop_mul_if_land_1_lpi_1_dfm_st_7 | (cfg_precision!=2'b10);
  assign or_dcpl_100 = or_tmp_608 | mul_loop_mul_if_land_2_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_19_lpi_1_dfm_st_3
      | (~ mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | or_dcpl_87;
  assign or_dcpl_103 = or_dcpl_95 | mul_loop_mul_if_land_2_lpi_1_dfm_st_7 | (cfg_precision!=2'b10);
  assign or_dcpl_107 = or_tmp_608 | mul_loop_mul_if_land_3_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_20_lpi_1_dfm_st_3
      | (~ mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | or_dcpl_87;
  assign or_dcpl_110 = or_dcpl_95 | mul_loop_mul_if_land_3_lpi_1_dfm_st_7 | (cfg_precision!=2'b10);
  assign or_dcpl_115 = or_tmp_608 | mul_loop_mul_if_land_4_lpi_1_dfm_st_7 | and_dcpl_50
      | FpMul_8U_23U_lor_21_lpi_1_dfm_st_3 | (~ mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | or_90_cse;
  assign or_dcpl_118 = or_dcpl_95 | mul_loop_mul_if_land_4_lpi_1_dfm_st_7 | (cfg_precision!=2'b10);
  assign or_dcpl_122 = or_tmp_608 | mul_loop_mul_if_land_5_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_22_lpi_1_dfm_st_3
      | (~ mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | or_dcpl_87;
  assign or_dcpl_125 = or_dcpl_95 | mul_loop_mul_if_land_5_lpi_1_dfm_st_7 | (cfg_precision!=2'b10);
  assign or_dcpl_129 = or_tmp_608 | mul_loop_mul_if_land_6_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_23_lpi_1_dfm_st_3
      | (~ mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | or_dcpl_87;
  assign or_dcpl_132 = or_dcpl_95 | mul_loop_mul_if_land_6_lpi_1_dfm_st_7 | (cfg_precision!=2'b10);
  assign or_dcpl_136 = or_tmp_608 | mul_loop_mul_if_land_7_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_24_lpi_1_dfm_st_3
      | (~ mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | or_dcpl_87;
  assign or_dcpl_139 = or_dcpl_95 | mul_loop_mul_if_land_7_lpi_1_dfm_st_7 | (cfg_precision!=2'b10);
  assign or_dcpl_143 = or_tmp_608 | mul_loop_mul_if_land_8_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_25_lpi_1_dfm_st_3
      | (~ mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | or_dcpl_87;
  assign or_dcpl_146 = or_dcpl_95 | mul_loop_mul_if_land_8_lpi_1_dfm_st_7 | (cfg_precision!=2'b10);
  assign or_dcpl_150 = or_tmp_608 | mul_loop_mul_if_land_9_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_26_lpi_1_dfm_st_3
      | (~ mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | or_dcpl_87;
  assign or_dcpl_153 = or_dcpl_95 | mul_loop_mul_if_land_9_lpi_1_dfm_st_7 | (cfg_precision!=2'b10);
  assign or_dcpl_157 = or_tmp_608 | mul_loop_mul_if_land_10_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_27_lpi_1_dfm_st_3
      | (~ mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | or_dcpl_87;
  assign or_dcpl_160 = or_dcpl_95 | mul_loop_mul_if_land_10_lpi_1_dfm_st_7 | (cfg_precision!=2'b10);
  assign or_dcpl_165 = or_tmp_608 | mul_loop_mul_if_land_11_lpi_1_dfm_st_7 | and_dcpl_50
      | FpMul_8U_23U_lor_28_lpi_1_dfm_st_3 | (~ mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | or_90_cse;
  assign or_dcpl_168 = or_dcpl_95 | mul_loop_mul_if_land_11_lpi_1_dfm_st_7 | (cfg_precision!=2'b10);
  assign or_dcpl_173 = or_tmp_608 | mul_loop_mul_if_land_12_lpi_1_dfm_st_7 | and_dcpl_50
      | FpMul_8U_23U_lor_29_lpi_1_dfm_st_3 | (~ mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | or_90_cse;
  assign or_dcpl_176 = or_dcpl_95 | mul_loop_mul_if_land_12_lpi_1_dfm_st_7 | (cfg_precision!=2'b10);
  assign or_dcpl_181 = or_tmp_608 | mul_loop_mul_if_land_13_lpi_1_dfm_st_7 | and_dcpl_50
      | FpMul_8U_23U_lor_30_lpi_1_dfm_st_3 | (~ mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | or_90_cse;
  assign or_dcpl_184 = or_dcpl_95 | mul_loop_mul_if_land_13_lpi_1_dfm_st_7 | (cfg_precision!=2'b10);
  assign or_dcpl_188 = or_tmp_608 | mul_loop_mul_if_land_14_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_31_lpi_1_dfm_st_3
      | (~ mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | or_dcpl_87;
  assign or_dcpl_191 = or_dcpl_95 | mul_loop_mul_if_land_14_lpi_1_dfm_st_7 | (cfg_precision!=2'b10);
  assign or_dcpl_195 = or_tmp_608 | mul_loop_mul_if_land_15_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_32_lpi_1_dfm_st_3
      | (~ mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | or_dcpl_87;
  assign or_dcpl_198 = or_dcpl_95 | mul_loop_mul_if_land_15_lpi_1_dfm_st_7 | (cfg_precision!=2'b10);
  assign or_dcpl_202 = or_tmp_608 | mul_loop_mul_if_land_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3
      | (~ mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | or_dcpl_87;
  assign or_dcpl_205 = or_dcpl_95 | mul_loop_mul_if_land_lpi_1_dfm_st_7 | (cfg_precision!=2'b10);
  assign and_dcpl_254 = (else_mux_2_tmp[3:2]==2'b11);
  assign and_dcpl_255 = (cfg_precision[1]) & (else_mux_2_tmp[4]);
  assign and_dcpl_258 = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_loop_mul_if_land_1_lpi_1_dfm_st_5);
  assign and_dcpl_259 = and_dcpl_258 & (~ (cfg_precision[0]));
  assign or_dcpl_206 = (~ cfg_nan_to_zero) | IsNaN_5U_10U_nor_tmp;
  assign and_dcpl_262 = or_309_cse & or_dcpl_206 & and_dcpl_259 & and_dcpl_255 &
      and_dcpl_254 & (else_mux_2_tmp[1:0]==2'b11) & (~ IsNaN_5U_23U_nor_tmp);
  assign and_dcpl_263 = and_dcpl_258 & and_dcpl_85;
  assign or_dcpl_212 = (cfg_nan_to_zero & (~ IsNaN_5U_10U_nor_tmp)) | (else_mux_2_tmp!=5'b11111)
      | IsNaN_5U_23U_nor_tmp;
  assign and_dcpl_266 = or_dcpl_212 & or_309_cse & and_dcpl_263;
  assign or_dcpl_216 = or_tmp_204 | and_dcpl_50;
  assign or_dcpl_217 = or_dcpl_216 | mul_loop_mul_if_land_1_lpi_1_dfm_st_6 | (cfg_precision!=2'b10);
  assign and_dcpl_269 = (else_mux_5_tmp[3:2]==2'b11);
  assign and_dcpl_270 = (cfg_precision[1]) & (else_mux_5_tmp[4]);
  assign and_dcpl_273 = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_loop_mul_if_land_2_lpi_1_dfm_st_5);
  assign and_dcpl_274 = and_dcpl_273 & (~ (cfg_precision[0]));
  assign or_dcpl_218 = IsNaN_5U_10U_nor_1_tmp | (~ cfg_nan_to_zero);
  assign and_dcpl_277 = or_309_cse & or_dcpl_218 & and_dcpl_274 & and_dcpl_270 &
      and_dcpl_269 & (else_mux_5_tmp[1:0]==2'b11) & (~ IsNaN_5U_23U_nor_1_tmp);
  assign and_dcpl_278 = and_dcpl_273 & and_dcpl_85;
  assign or_dcpl_224 = ((~ IsNaN_5U_10U_nor_1_tmp) & cfg_nan_to_zero) | (else_mux_5_tmp!=5'b11111)
      | IsNaN_5U_23U_nor_1_tmp;
  assign and_dcpl_281 = or_dcpl_224 & or_309_cse & and_dcpl_278;
  assign or_dcpl_227 = or_dcpl_216 | mul_loop_mul_if_land_2_lpi_1_dfm_st_6 | (cfg_precision!=2'b10);
  assign and_dcpl_284 = (else_mux_8_tmp[3:2]==2'b11);
  assign and_dcpl_285 = (cfg_precision[1]) & (else_mux_8_tmp[4]);
  assign and_dcpl_288 = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_loop_mul_if_land_3_lpi_1_dfm_st_5);
  assign and_dcpl_289 = and_dcpl_288 & (~ (cfg_precision[0]));
  assign or_dcpl_228 = IsNaN_5U_10U_nor_2_tmp | (~ cfg_nan_to_zero);
  assign and_dcpl_292 = or_309_cse & or_dcpl_228 & and_dcpl_289 & and_dcpl_285 &
      and_dcpl_284 & (else_mux_8_tmp[1:0]==2'b11) & (~ IsNaN_5U_23U_nor_2_tmp);
  assign and_dcpl_293 = and_dcpl_288 & and_dcpl_85;
  assign or_dcpl_234 = ((~ IsNaN_5U_10U_nor_2_tmp) & cfg_nan_to_zero) | (else_mux_8_tmp!=5'b11111)
      | IsNaN_5U_23U_nor_2_tmp;
  assign and_dcpl_296 = or_dcpl_234 & or_309_cse & and_dcpl_293;
  assign or_dcpl_237 = or_dcpl_216 | mul_loop_mul_if_land_3_lpi_1_dfm_st_6 | (cfg_precision!=2'b10);
  assign and_dcpl_299 = (else_mux_11_tmp[3:2]==2'b11);
  assign and_dcpl_300 = (cfg_precision[1]) & (else_mux_11_tmp[4]);
  assign and_dcpl_303 = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_loop_mul_if_land_4_lpi_1_dfm_st_5);
  assign and_dcpl_304 = and_dcpl_303 & (~ (cfg_precision[0]));
  assign or_dcpl_238 = IsNaN_5U_10U_nor_3_tmp | (~ cfg_nan_to_zero);
  assign and_dcpl_307 = or_309_cse & or_dcpl_238 & and_dcpl_304 & and_dcpl_300 &
      and_dcpl_299 & (else_mux_11_tmp[1:0]==2'b11) & (~ IsNaN_5U_23U_nor_3_tmp);
  assign and_dcpl_308 = and_dcpl_303 & and_dcpl_85;
  assign or_dcpl_244 = ((~ IsNaN_5U_10U_nor_3_tmp) & cfg_nan_to_zero) | (else_mux_11_tmp!=5'b11111)
      | IsNaN_5U_23U_nor_3_tmp;
  assign and_dcpl_311 = or_dcpl_244 & or_309_cse & and_dcpl_308;
  assign or_dcpl_247 = or_dcpl_216 | mul_loop_mul_if_land_4_lpi_1_dfm_st_6 | (cfg_precision!=2'b10);
  assign and_dcpl_314 = (else_mux_14_tmp[3:2]==2'b11);
  assign and_dcpl_315 = (cfg_precision[1]) & (else_mux_14_tmp[4]);
  assign and_dcpl_318 = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_loop_mul_if_land_5_lpi_1_dfm_st_5);
  assign and_dcpl_319 = and_dcpl_318 & (~ (cfg_precision[0]));
  assign or_dcpl_248 = IsNaN_5U_10U_nor_4_tmp | (~ cfg_nan_to_zero);
  assign and_dcpl_322 = or_309_cse & or_dcpl_248 & and_dcpl_319 & and_dcpl_315 &
      and_dcpl_314 & (else_mux_14_tmp[1:0]==2'b11) & (~ IsNaN_5U_23U_nor_4_tmp);
  assign and_dcpl_323 = and_dcpl_318 & and_dcpl_85;
  assign or_dcpl_254 = ((~ IsNaN_5U_10U_nor_4_tmp) & cfg_nan_to_zero) | (else_mux_14_tmp!=5'b11111)
      | IsNaN_5U_23U_nor_4_tmp;
  assign and_dcpl_326 = or_dcpl_254 & or_309_cse & and_dcpl_323;
  assign or_dcpl_257 = or_dcpl_216 | mul_loop_mul_if_land_5_lpi_1_dfm_st_6 | (cfg_precision!=2'b10);
  assign and_dcpl_329 = (else_mux_17_tmp[3:2]==2'b11);
  assign and_dcpl_330 = (cfg_precision[1]) & (else_mux_17_tmp[4]);
  assign and_dcpl_333 = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_loop_mul_if_land_6_lpi_1_dfm_st_5);
  assign and_dcpl_334 = and_dcpl_333 & (~ (cfg_precision[0]));
  assign or_dcpl_258 = IsNaN_5U_10U_nor_5_tmp | (~ cfg_nan_to_zero);
  assign and_dcpl_337 = or_309_cse & or_dcpl_258 & and_dcpl_334 & and_dcpl_330 &
      and_dcpl_329 & (else_mux_17_tmp[1:0]==2'b11) & (~ IsNaN_5U_23U_nor_5_tmp);
  assign and_dcpl_338 = and_dcpl_333 & and_dcpl_85;
  assign or_dcpl_264 = ((~ IsNaN_5U_10U_nor_5_tmp) & cfg_nan_to_zero) | (else_mux_17_tmp!=5'b11111)
      | IsNaN_5U_23U_nor_5_tmp;
  assign and_dcpl_341 = or_dcpl_264 & or_309_cse & and_dcpl_338;
  assign or_dcpl_267 = or_dcpl_216 | mul_loop_mul_if_land_6_lpi_1_dfm_st_6 | (cfg_precision!=2'b10);
  assign and_dcpl_344 = (else_mux_20_tmp[1:0]==2'b11);
  assign and_dcpl_345 = (else_mux_20_tmp[4:3]==2'b11);
  assign or_dcpl_268 = IsNaN_5U_10U_nor_6_tmp | (~ cfg_nan_to_zero);
  assign and_dcpl_349 = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_loop_mul_if_land_7_lpi_1_dfm_st_5);
  assign and_dcpl_352 = and_dcpl_349 & or_309_cse & or_dcpl_268 & (else_mux_20_tmp[2])
      & and_dcpl_345 & and_dcpl_344 & (~ IsNaN_5U_23U_nor_6_tmp) & (cfg_precision==2'b10);
  assign and_dcpl_353 = and_dcpl_349 & and_dcpl_85;
  assign or_dcpl_274 = (else_mux_20_tmp!=5'b11111) | IsNaN_5U_23U_nor_6_tmp | ((~
      IsNaN_5U_10U_nor_6_tmp) & cfg_nan_to_zero);
  assign and_dcpl_356 = or_dcpl_274 & or_309_cse & and_dcpl_353;
  assign or_dcpl_277 = or_dcpl_216 | mul_loop_mul_if_land_7_lpi_1_dfm_st_6 | (cfg_precision!=2'b10);
  assign and_dcpl_359 = (else_mux_23_tmp[1:0]==2'b11);
  assign and_dcpl_360 = (else_mux_23_tmp[3:2]==2'b11);
  assign or_dcpl_278 = IsNaN_5U_10U_nor_7_tmp | (~ cfg_nan_to_zero);
  assign and_dcpl_364 = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_loop_mul_if_land_8_lpi_1_dfm_st_5);
  assign and_dcpl_367 = and_dcpl_364 & or_309_cse & or_dcpl_278 & (else_mux_23_tmp[4])
      & and_dcpl_360 & and_dcpl_359 & (~ IsNaN_5U_23U_nor_7_tmp) & (cfg_precision==2'b10);
  assign and_dcpl_368 = and_dcpl_364 & and_dcpl_85;
  assign or_dcpl_284 = (else_mux_23_tmp!=5'b11111) | IsNaN_5U_23U_nor_7_tmp | ((~
      IsNaN_5U_10U_nor_7_tmp) & cfg_nan_to_zero);
  assign and_dcpl_371 = or_dcpl_284 & or_309_cse & and_dcpl_368;
  assign or_dcpl_287 = or_dcpl_216 | mul_loop_mul_if_land_8_lpi_1_dfm_st_6 | (cfg_precision!=2'b10);
  assign and_dcpl_374 = (else_mux_26_tmp[1:0]==2'b11);
  assign and_dcpl_375 = (else_mux_26_tmp[3:2]==2'b11);
  assign or_dcpl_288 = IsNaN_5U_10U_nor_8_tmp | (~ cfg_nan_to_zero);
  assign and_dcpl_379 = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_loop_mul_if_land_9_lpi_1_dfm_st_5);
  assign and_dcpl_382 = and_dcpl_379 & or_309_cse & or_dcpl_288 & (else_mux_26_tmp[4])
      & and_dcpl_375 & and_dcpl_374 & (~ IsNaN_5U_23U_nor_8_tmp) & (cfg_precision==2'b10);
  assign and_dcpl_383 = and_dcpl_379 & and_dcpl_85;
  assign or_dcpl_294 = (else_mux_26_tmp!=5'b11111) | IsNaN_5U_23U_nor_8_tmp | ((~
      IsNaN_5U_10U_nor_8_tmp) & cfg_nan_to_zero);
  assign and_dcpl_386 = or_dcpl_294 & or_309_cse & and_dcpl_383;
  assign or_dcpl_297 = or_dcpl_216 | mul_loop_mul_if_land_9_lpi_1_dfm_st_6 | (cfg_precision!=2'b10);
  assign and_dcpl_389 = (else_mux_29_tmp[4]) & (else_mux_29_tmp[1]);
  assign and_dcpl_390 = (cfg_precision[1]) & (~ IsNaN_5U_23U_nor_9_tmp);
  assign and_dcpl_393 = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_loop_mul_if_land_10_lpi_1_dfm_st_5);
  assign and_dcpl_394 = and_dcpl_393 & (~ (cfg_precision[0]));
  assign or_dcpl_298 = IsNaN_5U_10U_nor_9_tmp | (~ cfg_nan_to_zero);
  assign and_dcpl_397 = or_309_cse & or_dcpl_298 & and_dcpl_394 & and_dcpl_390 &
      and_dcpl_389 & (else_mux_29_tmp[3]) & (else_mux_29_tmp[2]) & (else_mux_29_tmp[0]);
  assign and_dcpl_398 = and_dcpl_393 & and_dcpl_85;
  assign or_dcpl_304 = ((~ IsNaN_5U_10U_nor_9_tmp) & cfg_nan_to_zero) | IsNaN_5U_23U_nor_9_tmp
      | (else_mux_29_tmp!=5'b11111);
  assign and_dcpl_401 = or_dcpl_304 & or_309_cse & and_dcpl_398;
  assign or_dcpl_307 = or_dcpl_216 | mul_loop_mul_if_land_10_lpi_1_dfm_st_6 | (cfg_precision!=2'b10);
  assign and_dcpl_404 = (else_mux_32_tmp[3:2]==2'b11);
  assign and_dcpl_405 = (cfg_precision[1]) & (~ IsNaN_5U_23U_nor_10_tmp);
  assign and_dcpl_408 = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_loop_mul_if_land_11_lpi_1_dfm_st_5);
  assign and_dcpl_409 = and_dcpl_408 & (~ (cfg_precision[0]));
  assign or_dcpl_308 = IsNaN_5U_10U_nor_10_tmp | (~ cfg_nan_to_zero);
  assign and_dcpl_412 = or_309_cse & or_dcpl_308 & and_dcpl_409 & and_dcpl_405 &
      and_dcpl_404 & (else_mux_32_tmp[1]) & (else_mux_32_tmp[0]) & (else_mux_32_tmp[4]);
  assign and_dcpl_413 = and_dcpl_408 & and_dcpl_85;
  assign or_dcpl_314 = ((~ IsNaN_5U_10U_nor_10_tmp) & cfg_nan_to_zero) | IsNaN_5U_23U_nor_10_tmp
      | (else_mux_32_tmp!=5'b11111);
  assign and_dcpl_416 = or_dcpl_314 & or_309_cse & and_dcpl_413;
  assign or_dcpl_317 = or_dcpl_216 | mul_loop_mul_if_land_11_lpi_1_dfm_st_6 | (cfg_precision!=2'b10);
  assign and_dcpl_419 = (else_mux_35_tmp[2]) & (else_mux_35_tmp[4]);
  assign and_dcpl_420 = (cfg_precision[1]) & (~ IsNaN_5U_23U_nor_11_tmp);
  assign and_dcpl_423 = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_loop_mul_if_land_12_lpi_1_dfm_st_5);
  assign and_dcpl_424 = and_dcpl_423 & (~ (cfg_precision[0]));
  assign or_dcpl_318 = IsNaN_5U_10U_nor_11_tmp | (~ cfg_nan_to_zero);
  assign and_dcpl_427 = or_309_cse & or_dcpl_318 & and_dcpl_424 & and_dcpl_420 &
      and_dcpl_419 & (else_mux_35_tmp[3]) & (else_mux_35_tmp[1]) & (else_mux_35_tmp[0]);
  assign and_dcpl_428 = and_dcpl_423 & and_dcpl_85;
  assign or_dcpl_324 = ((~ IsNaN_5U_10U_nor_11_tmp) & cfg_nan_to_zero) | IsNaN_5U_23U_nor_11_tmp
      | (else_mux_35_tmp!=5'b11111);
  assign and_dcpl_431 = or_dcpl_324 & or_309_cse & and_dcpl_428;
  assign or_dcpl_327 = or_dcpl_216 | mul_loop_mul_if_land_12_lpi_1_dfm_st_6 | (cfg_precision!=2'b10);
  assign and_dcpl_434 = (else_mux_38_tmp[4:3]==2'b11);
  assign and_dcpl_435 = (cfg_precision[1]) & (~ IsNaN_5U_23U_nor_12_tmp);
  assign and_dcpl_438 = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_loop_mul_if_land_13_lpi_1_dfm_st_5);
  assign and_dcpl_439 = and_dcpl_438 & (~ (cfg_precision[0]));
  assign or_dcpl_328 = IsNaN_5U_10U_nor_12_tmp | (~ cfg_nan_to_zero);
  assign and_dcpl_442 = or_309_cse & or_dcpl_328 & and_dcpl_439 & and_dcpl_435 &
      and_dcpl_434 & (else_mux_38_tmp[2:0]==3'b111);
  assign and_dcpl_443 = and_dcpl_438 & and_dcpl_85;
  assign or_dcpl_334 = ((~ IsNaN_5U_10U_nor_12_tmp) & cfg_nan_to_zero) | IsNaN_5U_23U_nor_12_tmp
      | (else_mux_38_tmp!=5'b11111);
  assign and_dcpl_446 = or_dcpl_334 & or_309_cse & and_dcpl_443;
  assign or_dcpl_337 = or_dcpl_216 | mul_loop_mul_if_land_13_lpi_1_dfm_st_6 | (cfg_precision!=2'b10);
  assign and_dcpl_449 = (else_mux_41_tmp[4]) & (else_mux_41_tmp[1]);
  assign and_dcpl_450 = (cfg_precision[1]) & (~ IsNaN_5U_23U_nor_13_tmp);
  assign and_dcpl_453 = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_loop_mul_if_land_14_lpi_1_dfm_st_5);
  assign and_dcpl_454 = and_dcpl_453 & (~ (cfg_precision[0]));
  assign or_dcpl_338 = IsNaN_5U_10U_nor_13_tmp | (~ cfg_nan_to_zero);
  assign and_dcpl_457 = or_309_cse & or_dcpl_338 & and_dcpl_454 & and_dcpl_450 &
      and_dcpl_449 & (else_mux_41_tmp[3]) & (else_mux_41_tmp[2]) & (else_mux_41_tmp[0]);
  assign and_dcpl_458 = and_dcpl_453 & and_dcpl_85;
  assign or_dcpl_344 = ((~ IsNaN_5U_10U_nor_13_tmp) & cfg_nan_to_zero) | IsNaN_5U_23U_nor_13_tmp
      | (else_mux_41_tmp!=5'b11111);
  assign and_dcpl_461 = or_dcpl_344 & or_309_cse & and_dcpl_458;
  assign or_dcpl_347 = or_dcpl_216 | mul_loop_mul_if_land_14_lpi_1_dfm_st_6 | (cfg_precision!=2'b10);
  assign and_dcpl_464 = (else_mux_44_tmp[3:2]==2'b11);
  assign and_dcpl_465 = (cfg_precision[1]) & (~ IsNaN_5U_23U_nor_14_tmp);
  assign and_dcpl_468 = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_loop_mul_if_land_15_lpi_1_dfm_st_5);
  assign and_dcpl_469 = and_dcpl_468 & (~ (cfg_precision[0]));
  assign or_dcpl_348 = IsNaN_5U_10U_nor_14_tmp | (~ cfg_nan_to_zero);
  assign and_dcpl_472 = or_309_cse & or_dcpl_348 & and_dcpl_469 & and_dcpl_465 &
      and_dcpl_464 & (else_mux_44_tmp[1]) & (else_mux_44_tmp[0]) & (else_mux_44_tmp[4]);
  assign and_dcpl_473 = and_dcpl_468 & and_dcpl_85;
  assign or_dcpl_354 = ((~ IsNaN_5U_10U_nor_14_tmp) & cfg_nan_to_zero) | IsNaN_5U_23U_nor_14_tmp
      | (else_mux_44_tmp!=5'b11111);
  assign and_dcpl_476 = or_dcpl_354 & or_309_cse & and_dcpl_473;
  assign or_dcpl_357 = or_dcpl_216 | mul_loop_mul_if_land_15_lpi_1_dfm_st_6 | (cfg_precision!=2'b10);
  assign and_dcpl_479 = (else_mux_47_tmp[2]) & (else_mux_47_tmp[4]);
  assign and_dcpl_480 = (cfg_precision[1]) & (~ IsNaN_5U_23U_nor_15_tmp);
  assign and_dcpl_483 = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_loop_mul_if_land_lpi_1_dfm_st_5);
  assign and_dcpl_484 = and_dcpl_483 & (~ (cfg_precision[0]));
  assign or_dcpl_358 = IsNaN_5U_10U_nor_15_tmp | (~ cfg_nan_to_zero);
  assign and_dcpl_487 = or_309_cse & or_dcpl_358 & and_dcpl_484 & and_dcpl_480 &
      and_dcpl_479 & (else_mux_47_tmp[3]) & (else_mux_47_tmp[1]) & (else_mux_47_tmp[0]);
  assign and_dcpl_488 = and_dcpl_483 & and_dcpl_85;
  assign or_dcpl_364 = ((~ IsNaN_5U_10U_nor_15_tmp) & cfg_nan_to_zero) | IsNaN_5U_23U_nor_15_tmp
      | (else_mux_47_tmp!=5'b11111);
  assign and_dcpl_491 = or_dcpl_364 & or_309_cse & and_dcpl_488;
  assign or_dcpl_367 = or_dcpl_216 | mul_loop_mul_if_land_lpi_1_dfm_st_6 | (cfg_precision!=2'b10);
  assign and_dcpl_492 = (~ chn_mul_op_rsci_bawt) & cfg_mul_src_1_sva_st_1;
  assign or_dcpl_369 = and_dcpl_492 | and_dcpl_50 | or_90_cse;
  assign or_dcpl_373 = or_dcpl_27 | or_tmp_10 | mul_loop_mul_if_land_1_lpi_1_dfm_st_5
      | or_dcpl_369;
  assign or_dcpl_382 = and_dcpl_50 | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign or_dcpl_385 = or_dcpl_27 | and_dcpl_492 | (~ main_stage_v_1);
  assign and_dcpl_494 = (~ cfg_mul_bypass_rsci_d) & (cfg_precision==2'b10);
  assign and_1042_nl = (nor_21_cse | cfg_mul_bypass_rsci_d) & or_dcpl_4;
  assign mux_1632_nl = MUX_s_1_2_2((and_1042_nl), or_dcpl_4, or_90_cse);
  assign and_dcpl_497 = (mux_1632_nl) & or_309_cse;
  assign and_1046_nl = (nor_23_cse | cfg_mul_bypass_rsci_d) & or_dcpl_4;
  assign mux_1633_nl = MUX_s_1_2_2((and_1046_nl), or_dcpl_4, or_90_cse);
  assign and_dcpl_500 = (mux_1633_nl) & or_309_cse;
  assign and_1050_nl = (nor_25_cse | cfg_mul_bypass_rsci_d) & or_dcpl_4;
  assign mux_1634_nl = MUX_s_1_2_2((and_1050_nl), or_dcpl_4, or_90_cse);
  assign and_dcpl_503 = (mux_1634_nl) & or_309_cse;
  assign and_1054_nl = (nor_26_cse | cfg_mul_bypass_rsci_d) & or_dcpl_4;
  assign mux_1635_nl = MUX_s_1_2_2((and_1054_nl), or_dcpl_4, or_90_cse);
  assign and_dcpl_506 = (mux_1635_nl) & or_309_cse;
  assign and_1058_nl = (nor_28_cse | cfg_mul_bypass_rsci_d) & or_dcpl_4;
  assign mux_1636_nl = MUX_s_1_2_2((and_1058_nl), or_dcpl_4, or_90_cse);
  assign and_dcpl_509 = (mux_1636_nl) & or_309_cse;
  assign and_1062_nl = (nor_29_cse | cfg_mul_bypass_rsci_d) & or_dcpl_4;
  assign mux_1637_nl = MUX_s_1_2_2((and_1062_nl), or_dcpl_4, or_90_cse);
  assign and_dcpl_512 = (mux_1637_nl) & or_309_cse;
  assign and_1066_nl = (nor_30_cse | cfg_mul_bypass_rsci_d) & or_dcpl_4;
  assign mux_1638_nl = MUX_s_1_2_2((and_1066_nl), or_dcpl_4, or_90_cse);
  assign and_dcpl_515 = (mux_1638_nl) & or_309_cse;
  assign and_1070_nl = (nor_32_cse | cfg_mul_bypass_rsci_d) & or_dcpl_4;
  assign mux_1639_nl = MUX_s_1_2_2((and_1070_nl), or_dcpl_4, or_90_cse);
  assign and_dcpl_518 = (mux_1639_nl) & or_309_cse;
  assign and_1074_nl = (nor_34_cse | cfg_mul_bypass_rsci_d) & or_dcpl_4;
  assign mux_1640_nl = MUX_s_1_2_2((and_1074_nl), or_dcpl_4, or_90_cse);
  assign and_dcpl_521 = (mux_1640_nl) & or_309_cse;
  assign and_1078_nl = (nor_35_cse | cfg_mul_bypass_rsci_d) & or_dcpl_4;
  assign mux_1641_nl = MUX_s_1_2_2((and_1078_nl), or_dcpl_4, or_90_cse);
  assign and_dcpl_524 = (mux_1641_nl) & or_309_cse;
  assign and_1082_nl = (nor_36_cse | cfg_mul_bypass_rsci_d) & or_dcpl_4;
  assign mux_1642_nl = MUX_s_1_2_2((and_1082_nl), or_dcpl_4, or_90_cse);
  assign and_dcpl_527 = (mux_1642_nl) & or_309_cse;
  assign and_1086_nl = (nor_37_cse | cfg_mul_bypass_rsci_d) & or_dcpl_4;
  assign mux_1643_nl = MUX_s_1_2_2((and_1086_nl), or_dcpl_4, or_90_cse);
  assign and_dcpl_530 = (mux_1643_nl) & or_309_cse;
  assign and_1090_nl = (nor_39_cse | cfg_mul_bypass_rsci_d) & or_dcpl_4;
  assign mux_1644_nl = MUX_s_1_2_2((and_1090_nl), or_dcpl_4, or_90_cse);
  assign and_dcpl_533 = (mux_1644_nl) & or_309_cse;
  assign and_1094_nl = (nor_40_cse | cfg_mul_bypass_rsci_d) & or_dcpl_4;
  assign mux_1645_nl = MUX_s_1_2_2((and_1094_nl), or_dcpl_4, or_90_cse);
  assign and_dcpl_536 = (mux_1645_nl) & or_309_cse;
  assign and_1098_nl = (nor_42_cse | cfg_mul_bypass_rsci_d) & or_dcpl_4;
  assign mux_1646_nl = MUX_s_1_2_2((and_1098_nl), or_dcpl_4, or_90_cse);
  assign and_dcpl_539 = (mux_1646_nl) & or_309_cse;
  assign and_1102_nl = (nor_44_cse | cfg_mul_bypass_rsci_d) & or_dcpl_4;
  assign mux_1647_nl = MUX_s_1_2_2((and_1102_nl), or_dcpl_4, or_90_cse);
  assign and_dcpl_542 = (mux_1647_nl) & or_309_cse;
  assign and_dcpl_546 = (~ io_read_cfg_mul_bypass_rsc_svs_st_5) & (~ mul_loop_mul_if_land_lpi_1_dfm_st_6)
      & or_309_cse;
  assign and_dcpl_555 = (~ io_read_cfg_mul_bypass_rsc_svs_st_5) & (~ mul_loop_mul_if_land_15_lpi_1_dfm_st_6)
      & or_309_cse;
  assign and_dcpl_564 = (~ io_read_cfg_mul_bypass_rsc_svs_st_5) & (~ mul_loop_mul_if_land_14_lpi_1_dfm_st_6)
      & or_309_cse;
  assign and_dcpl_573 = (~ io_read_cfg_mul_bypass_rsc_svs_st_5) & (~ mul_loop_mul_if_land_13_lpi_1_dfm_st_6)
      & or_309_cse;
  assign and_dcpl_582 = (~ io_read_cfg_mul_bypass_rsc_svs_st_5) & (~ mul_loop_mul_if_land_12_lpi_1_dfm_st_6)
      & or_309_cse;
  assign and_dcpl_591 = (~ io_read_cfg_mul_bypass_rsc_svs_st_5) & (~ mul_loop_mul_if_land_11_lpi_1_dfm_st_6)
      & or_309_cse;
  assign and_dcpl_600 = (~ io_read_cfg_mul_bypass_rsc_svs_st_5) & (~ mul_loop_mul_if_land_10_lpi_1_dfm_st_6)
      & or_309_cse;
  assign and_dcpl_609 = (~ io_read_cfg_mul_bypass_rsc_svs_st_5) & (~ mul_loop_mul_if_land_9_lpi_1_dfm_st_6)
      & or_309_cse;
  assign and_dcpl_618 = (~ io_read_cfg_mul_bypass_rsc_svs_st_5) & (~ mul_loop_mul_if_land_8_lpi_1_dfm_st_6)
      & or_309_cse;
  assign and_dcpl_627 = (~ io_read_cfg_mul_bypass_rsc_svs_st_5) & (~ mul_loop_mul_if_land_7_lpi_1_dfm_st_6)
      & or_309_cse;
  assign and_dcpl_636 = (~ io_read_cfg_mul_bypass_rsc_svs_st_5) & (~ mul_loop_mul_if_land_6_lpi_1_dfm_st_6)
      & or_309_cse;
  assign and_dcpl_645 = (~ io_read_cfg_mul_bypass_rsc_svs_st_5) & (~ mul_loop_mul_if_land_5_lpi_1_dfm_st_6)
      & or_309_cse;
  assign and_dcpl_654 = (~ io_read_cfg_mul_bypass_rsc_svs_st_5) & (~ mul_loop_mul_if_land_4_lpi_1_dfm_st_6)
      & or_309_cse;
  assign and_dcpl_663 = (~ io_read_cfg_mul_bypass_rsc_svs_st_5) & (~ mul_loop_mul_if_land_3_lpi_1_dfm_st_6)
      & or_309_cse;
  assign and_dcpl_672 = (~ io_read_cfg_mul_bypass_rsc_svs_st_5) & (~ mul_loop_mul_if_land_2_lpi_1_dfm_st_6)
      & or_309_cse;
  assign and_dcpl_681 = (~ io_read_cfg_mul_bypass_rsc_svs_st_5) & (~ mul_loop_mul_if_land_1_lpi_1_dfm_st_6)
      & or_309_cse;
  assign and_dcpl_770 = main_stage_v_2 & (~ io_read_cfg_mul_bypass_rsc_svs_st_5)
      & or_309_cse;
  assign and_dcpl_873 = or_2575_cse & cfg_mul_op_rsc_triosy_obj_bawt & or_309_cse
      & cfg_mul_bypass_rsc_triosy_obj_bawt;
  assign and_dcpl_879 = or_dcpl_212 & or_2575_cse & or_309_cse & nor_tmp_568 & and_dcpl_263;
  assign and_dcpl_891 = or_dcpl_224 & or_2575_cse & or_309_cse & nor_tmp_568 & and_dcpl_278;
  assign and_dcpl_903 = or_dcpl_234 & or_2575_cse & or_309_cse & nor_tmp_568 & and_dcpl_293;
  assign and_dcpl_915 = or_dcpl_244 & or_2575_cse & or_309_cse & nor_tmp_568 & and_dcpl_308;
  assign and_dcpl_927 = or_dcpl_254 & or_2575_cse & or_309_cse & nor_tmp_568 & and_dcpl_323;
  assign and_dcpl_939 = or_dcpl_264 & or_2575_cse & or_309_cse & nor_tmp_568 & and_dcpl_338;
  assign and_dcpl_951 = or_dcpl_274 & or_2575_cse & or_309_cse & nor_tmp_568 & and_dcpl_353;
  assign and_dcpl_963 = or_dcpl_284 & or_2575_cse & or_309_cse & nor_tmp_568 & and_dcpl_368;
  assign and_dcpl_975 = or_dcpl_294 & or_2575_cse & or_309_cse & nor_tmp_568 & and_dcpl_383;
  assign and_dcpl_987 = or_dcpl_304 & or_2575_cse & or_309_cse & nor_tmp_568 & and_dcpl_398;
  assign and_dcpl_999 = or_dcpl_314 & or_2575_cse & or_309_cse & nor_tmp_568 & and_dcpl_413;
  assign and_dcpl_1011 = or_dcpl_324 & or_2575_cse & or_309_cse & nor_tmp_568 & and_dcpl_428;
  assign and_dcpl_1023 = or_dcpl_334 & or_2575_cse & or_309_cse & nor_tmp_568 & and_dcpl_443;
  assign and_dcpl_1035 = or_dcpl_344 & or_2575_cse & or_309_cse & nor_tmp_568 & and_dcpl_458;
  assign and_dcpl_1047 = or_dcpl_354 & or_2575_cse & or_309_cse & nor_tmp_568 & and_dcpl_473;
  assign and_dcpl_1059 = or_dcpl_364 & or_2575_cse & or_309_cse & nor_tmp_568 & and_dcpl_488;
  assign or_dcpl_665 = cfg_mul_bypass_rsci_d | (cfg_precision!=2'b10) | (~ chn_mul_in_rsci_bawt);
  assign or_tmp_3606 = and_dcpl_7 & chn_mul_in_rsci_bawt & (fsm_output[1]);
  assign and_1647_cse = and_dcpl_7 & and_dcpl_59 & cfg_mul_src_rsci_d & (fsm_output[1]);
  assign chn_mul_in_rsci_ld_core_psct_mx0c0 = main_stage_en_1 | (fsm_output[0]);
  assign chn_mul_op_rsci_ld_core_psct_mx0c1 = and_dcpl_5 & or_309_cse & main_stage_v_1
      & and_dcpl_67 & (or_dcpl_31 | (~ cfg_mul_src_rsci_d));
  assign main_stage_v_1_mx0c1 = or_4649_cse & or_309_cse & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & main_stage_v_1 & (~ chn_mul_in_rsci_bawt);
  assign cfg_mul_src_1_sva_st_1_mx0c1 = (and_dcpl_7 & and_dcpl_91 & (fsm_output[1]))
      | (or_dcpl_4 & and_dcpl_47 & and_dcpl_91);
  assign main_stage_v_2_mx0c1 = (or_dcpl_27 | and_dcpl_52 | (~ main_stage_v_1)) &
      and_dcpl_95;
  assign main_stage_v_3_mx0c1 = main_stage_v_3 & (~ main_stage_v_2) & or_309_cse;
  assign main_stage_v_4_mx0c1 = (~ main_stage_v_3) & main_stage_v_4 & or_309_cse;
  assign FpMul_8U_23U_mux_12_itm_mx0c1 = and_dcpl_770 & (~(mul_loop_mul_if_land_1_lpi_1_dfm_st_6
      | IsNaN_8U_23U_land_1_lpi_1_dfm_9)) & and_dcpl_85;
  assign FpMul_8U_23U_mux_28_itm_mx0c1 = and_dcpl_770 & (~(mul_loop_mul_if_land_2_lpi_1_dfm_st_6
      | IsNaN_8U_23U_land_2_lpi_1_dfm_9)) & and_dcpl_85;
  assign FpMul_8U_23U_mux_44_itm_mx0c1 = and_dcpl_770 & (~(mul_loop_mul_if_land_3_lpi_1_dfm_st_6
      | IsNaN_8U_23U_land_3_lpi_1_dfm_9)) & and_dcpl_85;
  assign FpMul_8U_23U_mux_60_itm_mx0c1 = and_dcpl_770 & (~(mul_loop_mul_if_land_4_lpi_1_dfm_st_6
      | IsNaN_8U_23U_land_4_lpi_1_dfm_9)) & and_dcpl_85;
  assign FpMul_8U_23U_mux_76_itm_mx0c1 = and_dcpl_770 & (~(mul_loop_mul_if_land_5_lpi_1_dfm_st_6
      | IsNaN_8U_23U_land_5_lpi_1_dfm_9)) & and_dcpl_85;
  assign FpMul_8U_23U_mux_92_itm_mx0c1 = and_dcpl_770 & (~(mul_loop_mul_if_land_6_lpi_1_dfm_st_6
      | IsNaN_8U_23U_land_6_lpi_1_dfm_9)) & and_dcpl_85;
  assign FpMul_8U_23U_mux_108_itm_mx0c1 = and_dcpl_770 & (~(mul_loop_mul_if_land_7_lpi_1_dfm_st_6
      | IsNaN_8U_23U_land_7_lpi_1_dfm_9)) & and_dcpl_85;
  assign FpMul_8U_23U_mux_124_itm_mx0c1 = and_dcpl_770 & (~(mul_loop_mul_if_land_8_lpi_1_dfm_st_6
      | IsNaN_8U_23U_land_8_lpi_1_dfm_9)) & and_dcpl_85;
  assign FpMul_8U_23U_mux_140_itm_mx0c1 = and_dcpl_770 & (~(mul_loop_mul_if_land_9_lpi_1_dfm_st_6
      | IsNaN_8U_23U_land_9_lpi_1_dfm_9)) & and_dcpl_85;
  assign FpMul_8U_23U_mux_156_itm_mx0c1 = and_dcpl_770 & (~(mul_loop_mul_if_land_10_lpi_1_dfm_st_6
      | IsNaN_8U_23U_land_10_lpi_1_dfm_9)) & and_dcpl_85;
  assign FpMul_8U_23U_mux_172_itm_mx0c1 = and_dcpl_770 & (~(mul_loop_mul_if_land_11_lpi_1_dfm_st_6
      | IsNaN_8U_23U_land_11_lpi_1_dfm_9)) & and_dcpl_85;
  assign FpMul_8U_23U_mux_188_itm_mx0c1 = and_dcpl_770 & (~(mul_loop_mul_if_land_12_lpi_1_dfm_st_6
      | IsNaN_8U_23U_land_12_lpi_1_dfm_9)) & and_dcpl_85;
  assign FpMul_8U_23U_mux_204_itm_mx0c1 = and_dcpl_770 & (~(mul_loop_mul_if_land_13_lpi_1_dfm_st_6
      | IsNaN_8U_23U_land_13_lpi_1_dfm_9)) & and_dcpl_85;
  assign FpMul_8U_23U_mux_220_itm_mx0c1 = and_dcpl_770 & (~(mul_loop_mul_if_land_14_lpi_1_dfm_st_6
      | IsNaN_8U_23U_land_14_lpi_1_dfm_9)) & and_dcpl_85;
  assign FpMul_8U_23U_mux_236_itm_mx0c1 = and_dcpl_770 & (~(mul_loop_mul_if_land_15_lpi_1_dfm_st_6
      | IsNaN_8U_23U_land_15_lpi_1_dfm_9)) & and_dcpl_85;
  assign FpMul_8U_23U_mux_252_itm_mx0c1 = and_dcpl_770 & (~(mul_loop_mul_if_land_lpi_1_dfm_st_6
      | IsNaN_8U_23U_land_lpi_1_dfm_9)) & and_dcpl_85;
  assign chn_mul_in_rsci_oswt_unreg = or_tmp_3606;
  assign chn_mul_op_rsci_oswt_unreg = nor_tmp_568 & and_dcpl_67 & or_309_cse;
  assign chn_mul_out_rsci_oswt_unreg = and_dcpl_47;
  assign cfg_mul_op_rsc_triosy_obj_oswt_unreg_pff = and_dcpl_75;
  assign not_tmp_1326 = ~(mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & mux_1690_cse);
  assign not_tmp_1344 = ~(mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & mux_1695_cse);
  assign not_tmp_1362 = ~(mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & mux_1700_cse);
  assign not_tmp_1380 = ~(mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & mux_1705_cse);
  assign not_tmp_1398 = ~(mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & mux_1710_cse);
  assign not_tmp_1416 = ~(mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & mux_1715_cse);
  assign not_tmp_1434 = ~(mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & mux_1720_cse);
  assign not_tmp_1452 = ~(mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & mux_1725_cse);
  assign not_tmp_1470 = ~(mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & mux_1730_cse);
  assign not_tmp_1488 = ~(mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & mux_1735_cse);
  assign not_tmp_1506 = ~(mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & mux_1741_cse);
  assign not_tmp_1524 = ~(mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & mux_1747_cse);
  assign not_tmp_1542 = ~(mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & mux_1752_cse);
  assign not_tmp_1578 = ~(mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & mux_1764_cse);
  assign not_tmp_1596 = ~(mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & mux_1769_cse);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_in_rsci_iswt0 <= 1'b0;
      reg_cfg_mul_src_rsc_triosy_obj_ld_core_psct_cse <= 1'b0;
      chn_mul_out_rsci_iswt0 <= 1'b0;
      chn_mul_op_rsci_iswt0 <= 1'b0;
    end
    else if ( core_wen ) begin
      chn_mul_in_rsci_iswt0 <= ~((~ main_stage_en_1) & (fsm_output[1]));
      reg_cfg_mul_src_rsc_triosy_obj_ld_core_psct_cse <= or_tmp_3606;
      chn_mul_out_rsci_iswt0 <= and_dcpl_56;
      chn_mul_op_rsci_iswt0 <= and_1647_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_in_rsci_ld_core_psct <= 1'b0;
    end
    else if ( core_wen & chn_mul_in_rsci_ld_core_psct_mx0c0 ) begin
      chn_mul_in_rsci_ld_core_psct <= chn_mul_in_rsci_ld_core_psct_mx0c0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_out_rsci_d_9_0 <= 10'b0;
      chn_mul_out_rsci_d_12_10 <= 3'b0;
      chn_mul_out_rsci_d_22_13 <= 10'b0;
      chn_mul_out_rsci_d_26_23 <= 4'b0;
      chn_mul_out_rsci_d_28_27 <= 2'b0;
      chn_mul_out_rsci_d_30_29 <= 2'b0;
      chn_mul_out_rsci_d_48_31 <= 18'b0;
      chn_mul_out_rsci_d_58_49 <= 10'b0;
      chn_mul_out_rsci_d_61_59 <= 3'b0;
      chn_mul_out_rsci_d_71_62 <= 10'b0;
      chn_mul_out_rsci_d_75_72 <= 4'b0;
      chn_mul_out_rsci_d_77_76 <= 2'b0;
      chn_mul_out_rsci_d_79_78 <= 2'b0;
      chn_mul_out_rsci_d_97_80 <= 18'b0;
      chn_mul_out_rsci_d_107_98 <= 10'b0;
      chn_mul_out_rsci_d_110_108 <= 3'b0;
      chn_mul_out_rsci_d_120_111 <= 10'b0;
      chn_mul_out_rsci_d_124_121 <= 4'b0;
      chn_mul_out_rsci_d_126_125 <= 2'b0;
      chn_mul_out_rsci_d_128_127 <= 2'b0;
      chn_mul_out_rsci_d_146_129 <= 18'b0;
      chn_mul_out_rsci_d_156_147 <= 10'b0;
      chn_mul_out_rsci_d_159_157 <= 3'b0;
      chn_mul_out_rsci_d_169_160 <= 10'b0;
      chn_mul_out_rsci_d_173_170 <= 4'b0;
      chn_mul_out_rsci_d_175_174 <= 2'b0;
      chn_mul_out_rsci_d_177_176 <= 2'b0;
      chn_mul_out_rsci_d_195_178 <= 18'b0;
      chn_mul_out_rsci_d_205_196 <= 10'b0;
      chn_mul_out_rsci_d_208_206 <= 3'b0;
      chn_mul_out_rsci_d_218_209 <= 10'b0;
      chn_mul_out_rsci_d_222_219 <= 4'b0;
      chn_mul_out_rsci_d_224_223 <= 2'b0;
      chn_mul_out_rsci_d_226_225 <= 2'b0;
      chn_mul_out_rsci_d_244_227 <= 18'b0;
      chn_mul_out_rsci_d_254_245 <= 10'b0;
      chn_mul_out_rsci_d_257_255 <= 3'b0;
      chn_mul_out_rsci_d_267_258 <= 10'b0;
      chn_mul_out_rsci_d_271_268 <= 4'b0;
      chn_mul_out_rsci_d_273_272 <= 2'b0;
      chn_mul_out_rsci_d_275_274 <= 2'b0;
      chn_mul_out_rsci_d_293_276 <= 18'b0;
      chn_mul_out_rsci_d_303_294 <= 10'b0;
      chn_mul_out_rsci_d_306_304 <= 3'b0;
      chn_mul_out_rsci_d_316_307 <= 10'b0;
      chn_mul_out_rsci_d_320_317 <= 4'b0;
      chn_mul_out_rsci_d_322_321 <= 2'b0;
      chn_mul_out_rsci_d_324_323 <= 2'b0;
      chn_mul_out_rsci_d_342_325 <= 18'b0;
      chn_mul_out_rsci_d_352_343 <= 10'b0;
      chn_mul_out_rsci_d_355_353 <= 3'b0;
      chn_mul_out_rsci_d_365_356 <= 10'b0;
      chn_mul_out_rsci_d_369_366 <= 4'b0;
      chn_mul_out_rsci_d_371_370 <= 2'b0;
      chn_mul_out_rsci_d_373_372 <= 2'b0;
      chn_mul_out_rsci_d_391_374 <= 18'b0;
      chn_mul_out_rsci_d_401_392 <= 10'b0;
      chn_mul_out_rsci_d_404_402 <= 3'b0;
      chn_mul_out_rsci_d_414_405 <= 10'b0;
      chn_mul_out_rsci_d_418_415 <= 4'b0;
      chn_mul_out_rsci_d_420_419 <= 2'b0;
      chn_mul_out_rsci_d_422_421 <= 2'b0;
      chn_mul_out_rsci_d_440_423 <= 18'b0;
      chn_mul_out_rsci_d_450_441 <= 10'b0;
      chn_mul_out_rsci_d_453_451 <= 3'b0;
      chn_mul_out_rsci_d_463_454 <= 10'b0;
      chn_mul_out_rsci_d_467_464 <= 4'b0;
      chn_mul_out_rsci_d_469_468 <= 2'b0;
      chn_mul_out_rsci_d_471_470 <= 2'b0;
      chn_mul_out_rsci_d_489_472 <= 18'b0;
      chn_mul_out_rsci_d_499_490 <= 10'b0;
      chn_mul_out_rsci_d_502_500 <= 3'b0;
      chn_mul_out_rsci_d_512_503 <= 10'b0;
      chn_mul_out_rsci_d_516_513 <= 4'b0;
      chn_mul_out_rsci_d_518_517 <= 2'b0;
      chn_mul_out_rsci_d_520_519 <= 2'b0;
      chn_mul_out_rsci_d_538_521 <= 18'b0;
      chn_mul_out_rsci_d_548_539 <= 10'b0;
      chn_mul_out_rsci_d_551_549 <= 3'b0;
      chn_mul_out_rsci_d_561_552 <= 10'b0;
      chn_mul_out_rsci_d_565_562 <= 4'b0;
      chn_mul_out_rsci_d_567_566 <= 2'b0;
      chn_mul_out_rsci_d_569_568 <= 2'b0;
      chn_mul_out_rsci_d_587_570 <= 18'b0;
      chn_mul_out_rsci_d_597_588 <= 10'b0;
      chn_mul_out_rsci_d_600_598 <= 3'b0;
      chn_mul_out_rsci_d_610_601 <= 10'b0;
      chn_mul_out_rsci_d_614_611 <= 4'b0;
      chn_mul_out_rsci_d_616_615 <= 2'b0;
      chn_mul_out_rsci_d_618_617 <= 2'b0;
      chn_mul_out_rsci_d_636_619 <= 18'b0;
      chn_mul_out_rsci_d_646_637 <= 10'b0;
      chn_mul_out_rsci_d_649_647 <= 3'b0;
      chn_mul_out_rsci_d_659_650 <= 10'b0;
      chn_mul_out_rsci_d_663_660 <= 4'b0;
      chn_mul_out_rsci_d_665_664 <= 2'b0;
      chn_mul_out_rsci_d_667_666 <= 2'b0;
      chn_mul_out_rsci_d_685_668 <= 18'b0;
      chn_mul_out_rsci_d_695_686 <= 10'b0;
      chn_mul_out_rsci_d_698_696 <= 3'b0;
      chn_mul_out_rsci_d_708_699 <= 10'b0;
      chn_mul_out_rsci_d_712_709 <= 4'b0;
      chn_mul_out_rsci_d_714_713 <= 2'b0;
      chn_mul_out_rsci_d_716_715 <= 2'b0;
      chn_mul_out_rsci_d_734_717 <= 18'b0;
      chn_mul_out_rsci_d_744_735 <= 10'b0;
      chn_mul_out_rsci_d_747_745 <= 3'b0;
      chn_mul_out_rsci_d_757_748 <= 10'b0;
      chn_mul_out_rsci_d_761_758 <= 4'b0;
      chn_mul_out_rsci_d_763_762 <= 2'b0;
      chn_mul_out_rsci_d_765_764 <= 2'b0;
      chn_mul_out_rsci_d_783_766 <= 18'b0;
      chn_mul_out_rsci_d_784 <= 1'b0;
      chn_mul_out_rsci_d_785 <= 1'b0;
      chn_mul_out_rsci_d_786 <= 1'b0;
      chn_mul_out_rsci_d_787 <= 1'b0;
      chn_mul_out_rsci_d_788 <= 1'b0;
      chn_mul_out_rsci_d_789 <= 1'b0;
      chn_mul_out_rsci_d_790 <= 1'b0;
      chn_mul_out_rsci_d_791 <= 1'b0;
      chn_mul_out_rsci_d_792 <= 1'b0;
      chn_mul_out_rsci_d_793 <= 1'b0;
      chn_mul_out_rsci_d_794 <= 1'b0;
      chn_mul_out_rsci_d_795 <= 1'b0;
      chn_mul_out_rsci_d_796 <= 1'b0;
      chn_mul_out_rsci_d_797 <= 1'b0;
      chn_mul_out_rsci_d_798 <= 1'b0;
      chn_mul_out_rsci_d_799 <= 1'b0;
    end
    else if ( chn_mul_out_and_cse ) begin
      chn_mul_out_rsci_d_9_0 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_33_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_9_9_0_1, (MulIn_data_sva_536[9:0]),
          (MulOut_data_0_sva_10[9:0]), {and_2496_cse , and_2497_cse , or_4733_cse
          , asn_1163});
      chn_mul_out_rsci_d_12_10 <= MUX1HOT_v_3_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_32_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_9_12_10_1, (MulIn_data_sva_536[12:10]),
          (MulOut_data_0_sva_10[12:10]), {and_2496_cse , and_2497_cse , or_4733_cse
          , asn_1163});
      chn_mul_out_rsci_d_22_13 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_16_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_9_22_13_1, (MulIn_data_sva_536[22:13]),
          (MulOut_data_0_sva_10[22:13]), {and_2496_cse , and_2497_cse , or_4733_cse
          , asn_1163});
      chn_mul_out_rsci_d_26_23 <= MUX1HOT_v_4_4_2((FpMul_8U_23U_FpMul_8U_23U_and_95_nl),
          reg_FpMul_8U_23U_p_expo_1_2_itm, (MulIn_data_sva_536[26:23]), (MulOut_data_0_sva_10[26:23]),
          {and_2488_cse , and_2489_cse , or_4733_cse , asn_1163});
      chn_mul_out_rsci_d_28_27 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_97_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_9_1_0_1, (MulIn_data_sva_536[28:27]),
          (MulOut_data_0_sva_10[28:27]), {and_2488_cse , and_2489_cse , or_4733_cse
          , asn_1163});
      chn_mul_out_rsci_d_30_29 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_96_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_9_3_2_1, (MulIn_data_sva_536[30:29]),
          (MulOut_data_0_sva_10[30:29]), {and_2488_cse , and_2489_cse , or_4733_cse
          , asn_1163});
      chn_mul_out_rsci_d_48_31 <= MUX1HOT_v_18_3_2(({{17{FpMul_8U_23U_mux_12_itm_4}},
          FpMul_8U_23U_mux_12_itm_4}), (signext_18_2(MulIn_data_sva_536[32:31])),
          (MulOut_data_0_sva_10[48:31]), {and_116_ssc , or_17_ssc , asn_1163});
      chn_mul_out_rsci_d_58_49 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_35_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_9_9_0_1, (MulIn_data_sva_536[42:33]),
          (MulOut_data_1_sva_10[9:0]), {and_2481_cse , and_2482_cse , or_4729_cse
          , asn_1173});
      chn_mul_out_rsci_d_61_59 <= MUX1HOT_v_3_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_34_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_9_12_10_1, (MulIn_data_sva_536[45:43]),
          (MulOut_data_1_sva_10[12:10]), {and_2481_cse , and_2482_cse , or_4729_cse
          , asn_1173});
      chn_mul_out_rsci_d_71_62 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_17_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_9_22_13_1, (MulIn_data_sva_536[55:46]),
          (MulOut_data_1_sva_10[22:13]), {and_2481_cse , and_2482_cse , or_4729_cse
          , asn_1173});
      chn_mul_out_rsci_d_75_72 <= MUX1HOT_v_4_4_2((FpMul_8U_23U_FpMul_8U_23U_and_98_nl),
          reg_FpMul_8U_23U_p_expo_2_2_itm, (MulIn_data_sva_536[59:56]), (MulOut_data_1_sva_10[26:23]),
          {and_2473_cse , and_2474_cse , or_4729_cse , asn_1173});
      chn_mul_out_rsci_d_77_76 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_100_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_9_1_0_1, (MulIn_data_sva_536[61:60]),
          (MulOut_data_1_sva_10[28:27]), {and_2473_cse , and_2474_cse , or_4729_cse
          , asn_1173});
      chn_mul_out_rsci_d_79_78 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_99_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_9_3_2_1, (MulIn_data_sva_536[63:62]),
          (MulOut_data_1_sva_10[30:29]), {and_2473_cse , and_2474_cse , or_4729_cse
          , asn_1173});
      chn_mul_out_rsci_d_97_80 <= MUX1HOT_v_18_3_2(({{17{FpMul_8U_23U_mux_28_itm_4}},
          FpMul_8U_23U_mux_28_itm_4}), (signext_18_2(MulIn_data_sva_536[65:64])),
          (MulOut_data_1_sva_10[48:31]), {and_51_ssc , or_1_ssc , asn_1173});
      chn_mul_out_rsci_d_107_98 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_37_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_9_9_0_1, (MulIn_data_sva_536[75:66]),
          (MulOut_data_2_sva_10[9:0]), {and_2466_cse , and_2467_cse , or_4725_cse
          , asn_1183});
      chn_mul_out_rsci_d_110_108 <= MUX1HOT_v_3_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_36_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_9_12_10_1, (MulIn_data_sva_536[78:76]),
          (MulOut_data_2_sva_10[12:10]), {and_2466_cse , and_2467_cse , or_4725_cse
          , asn_1183});
      chn_mul_out_rsci_d_120_111 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_18_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_9_22_13_1, (MulIn_data_sva_536[88:79]),
          (MulOut_data_2_sva_10[22:13]), {and_2466_cse , and_2467_cse , or_4725_cse
          , asn_1183});
      chn_mul_out_rsci_d_124_121 <= MUX1HOT_v_4_4_2((FpMul_8U_23U_FpMul_8U_23U_and_101_nl),
          reg_FpMul_8U_23U_p_expo_3_2_itm, (MulIn_data_sva_536[92:89]), (MulOut_data_2_sva_10[26:23]),
          {and_2458_cse , and_2459_cse , or_4725_cse , asn_1183});
      chn_mul_out_rsci_d_126_125 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_103_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_9_1_0_1, (MulIn_data_sva_536[94:93]),
          (MulOut_data_2_sva_10[28:27]), {and_2458_cse , and_2459_cse , or_4725_cse
          , asn_1183});
      chn_mul_out_rsci_d_128_127 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_102_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_9_3_2_1, (MulIn_data_sva_536[96:95]),
          (MulOut_data_2_sva_10[30:29]), {and_2458_cse , and_2459_cse , or_4725_cse
          , asn_1183});
      chn_mul_out_rsci_d_146_129 <= MUX1HOT_v_18_3_2(({{17{FpMul_8U_23U_mux_44_itm_4}},
          FpMul_8U_23U_mux_44_itm_4}), (signext_18_2(MulIn_data_sva_536[98:97])),
          (MulOut_data_2_sva_10[48:31]), {and_55_ssc , or_2_ssc , asn_1183});
      chn_mul_out_rsci_d_156_147 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_39_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_9_9_0_1, (MulIn_data_sva_536[108:99]),
          (MulOut_data_3_sva_10[9:0]), {and_2451_cse , and_2452_cse , or_4721_cse
          , asn_1193});
      chn_mul_out_rsci_d_159_157 <= MUX1HOT_v_3_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_38_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_9_12_10_1, (MulIn_data_sva_536[111:109]),
          (MulOut_data_3_sva_10[12:10]), {and_2451_cse , and_2452_cse , or_4721_cse
          , asn_1193});
      chn_mul_out_rsci_d_169_160 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_19_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_9_22_13_1, (MulIn_data_sva_536[121:112]),
          (MulOut_data_3_sva_10[22:13]), {and_2451_cse , and_2452_cse , or_4721_cse
          , asn_1193});
      chn_mul_out_rsci_d_173_170 <= MUX1HOT_v_4_4_2((FpMul_8U_23U_FpMul_8U_23U_and_104_nl),
          reg_FpMul_8U_23U_p_expo_4_2_itm, (MulIn_data_sva_536[125:122]), (MulOut_data_3_sva_10[26:23]),
          {and_2443_cse , and_2444_cse , or_4721_cse , asn_1193});
      chn_mul_out_rsci_d_175_174 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_106_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_9_1_0_1, (MulIn_data_sva_536[127:126]),
          (MulOut_data_3_sva_10[28:27]), {and_2443_cse , and_2444_cse , or_4721_cse
          , asn_1193});
      chn_mul_out_rsci_d_177_176 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_105_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_9_3_2_1, (MulIn_data_sva_536[129:128]),
          (MulOut_data_3_sva_10[30:29]), {and_2443_cse , and_2444_cse , or_4721_cse
          , asn_1193});
      chn_mul_out_rsci_d_195_178 <= MUX1HOT_v_18_3_2(({{17{FpMul_8U_23U_mux_60_itm_4}},
          FpMul_8U_23U_mux_60_itm_4}), (signext_18_2(MulIn_data_sva_536[131:130])),
          (MulOut_data_3_sva_10[48:31]), {and_59_ssc , or_3_ssc , asn_1193});
      chn_mul_out_rsci_d_205_196 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_41_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_9_9_0_1, (MulIn_data_sva_536[141:132]),
          (MulOut_data_4_sva_10[9:0]), {and_2436_cse , and_2437_cse , or_4717_cse
          , asn_1203});
      chn_mul_out_rsci_d_208_206 <= MUX1HOT_v_3_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_40_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_9_12_10_1, (MulIn_data_sva_536[144:142]),
          (MulOut_data_4_sva_10[12:10]), {and_2436_cse , and_2437_cse , or_4717_cse
          , asn_1203});
      chn_mul_out_rsci_d_218_209 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_20_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_9_22_13_1, (MulIn_data_sva_536[154:145]),
          (MulOut_data_4_sva_10[22:13]), {and_2436_cse , and_2437_cse , or_4717_cse
          , asn_1203});
      chn_mul_out_rsci_d_222_219 <= MUX1HOT_v_4_4_2((FpMul_8U_23U_FpMul_8U_23U_and_107_nl),
          reg_FpMul_8U_23U_p_expo_5_2_itm, (MulIn_data_sva_536[158:155]), (MulOut_data_4_sva_10[26:23]),
          {and_2428_cse , and_2429_cse , or_4717_cse , asn_1203});
      chn_mul_out_rsci_d_224_223 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_109_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_9_1_0_1, (MulIn_data_sva_536[160:159]),
          (MulOut_data_4_sva_10[28:27]), {and_2428_cse , and_2429_cse , or_4717_cse
          , asn_1203});
      chn_mul_out_rsci_d_226_225 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_108_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_9_3_2_1, (MulIn_data_sva_536[162:161]),
          (MulOut_data_4_sva_10[30:29]), {and_2428_cse , and_2429_cse , or_4717_cse
          , asn_1203});
      chn_mul_out_rsci_d_244_227 <= MUX1HOT_v_18_3_2(({{17{FpMul_8U_23U_mux_76_itm_4}},
          FpMul_8U_23U_mux_76_itm_4}), (signext_18_2(MulIn_data_sva_536[164:163])),
          (MulOut_data_4_sva_10[48:31]), {and_63_ssc , or_4_ssc , asn_1203});
      chn_mul_out_rsci_d_254_245 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_43_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_9_9_0_1, (MulIn_data_sva_536[174:165]),
          (MulOut_data_5_sva_10[9:0]), {and_2421_cse , and_2422_cse , or_4713_cse
          , asn_1213});
      chn_mul_out_rsci_d_257_255 <= MUX1HOT_v_3_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_42_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_9_12_10_1, (MulIn_data_sva_536[177:175]),
          (MulOut_data_5_sva_10[12:10]), {and_2421_cse , and_2422_cse , or_4713_cse
          , asn_1213});
      chn_mul_out_rsci_d_267_258 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_21_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_9_22_13_1, (MulIn_data_sva_536[187:178]),
          (MulOut_data_5_sva_10[22:13]), {and_2421_cse , and_2422_cse , or_4713_cse
          , asn_1213});
      chn_mul_out_rsci_d_271_268 <= MUX1HOT_v_4_4_2((FpMul_8U_23U_FpMul_8U_23U_and_110_nl),
          reg_FpMul_8U_23U_p_expo_6_2_itm, (MulIn_data_sva_536[191:188]), (MulOut_data_5_sva_10[26:23]),
          {and_2413_cse , and_2414_cse , or_4713_cse , asn_1213});
      chn_mul_out_rsci_d_273_272 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_112_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_9_1_0_1, (MulIn_data_sva_536[193:192]),
          (MulOut_data_5_sva_10[28:27]), {and_2413_cse , and_2414_cse , or_4713_cse
          , asn_1213});
      chn_mul_out_rsci_d_275_274 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_111_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_9_3_2_1, (MulIn_data_sva_536[195:194]),
          (MulOut_data_5_sva_10[30:29]), {and_2413_cse , and_2414_cse , or_4713_cse
          , asn_1213});
      chn_mul_out_rsci_d_293_276 <= MUX1HOT_v_18_3_2(({{17{FpMul_8U_23U_mux_92_itm_4}},
          FpMul_8U_23U_mux_92_itm_4}), (signext_18_2(MulIn_data_sva_536[197:196])),
          (MulOut_data_5_sva_10[48:31]), {and_67_ssc , or_5_ssc , asn_1213});
      chn_mul_out_rsci_d_303_294 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_45_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_9_9_0_1, (MulIn_data_sva_536[207:198]),
          (MulOut_data_6_sva_10[9:0]), {and_2406_cse , and_2407_cse , or_4709_cse
          , asn_1223});
      chn_mul_out_rsci_d_306_304 <= MUX1HOT_v_3_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_44_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_9_12_10_1, (MulIn_data_sva_536[210:208]),
          (MulOut_data_6_sva_10[12:10]), {and_2406_cse , and_2407_cse , or_4709_cse
          , asn_1223});
      chn_mul_out_rsci_d_316_307 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_22_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_9_22_13_1, (MulIn_data_sva_536[220:211]),
          (MulOut_data_6_sva_10[22:13]), {and_2406_cse , and_2407_cse , or_4709_cse
          , asn_1223});
      chn_mul_out_rsci_d_320_317 <= MUX1HOT_v_4_4_2((FpMul_8U_23U_FpMul_8U_23U_and_113_nl),
          reg_FpMul_8U_23U_p_expo_7_2_itm, (MulIn_data_sva_536[224:221]), (MulOut_data_6_sva_10[26:23]),
          {and_2398_cse , and_2399_cse , or_4709_cse , asn_1223});
      chn_mul_out_rsci_d_322_321 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_115_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_9_1_0_1, (MulIn_data_sva_536[226:225]),
          (MulOut_data_6_sva_10[28:27]), {and_2398_cse , and_2399_cse , or_4709_cse
          , asn_1223});
      chn_mul_out_rsci_d_324_323 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_114_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_9_3_2_1, (MulIn_data_sva_536[228:227]),
          (MulOut_data_6_sva_10[30:29]), {and_2398_cse , and_2399_cse , or_4709_cse
          , asn_1223});
      chn_mul_out_rsci_d_342_325 <= MUX1HOT_v_18_3_2(({{17{FpMul_8U_23U_mux_108_itm_4}},
          FpMul_8U_23U_mux_108_itm_4}), (signext_18_2(MulIn_data_sva_536[230:229])),
          (MulOut_data_6_sva_10[48:31]), {and_71_ssc , or_6_ssc , asn_1223});
      chn_mul_out_rsci_d_352_343 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_47_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_9_9_0_1, (MulIn_data_sva_536[240:231]),
          (MulOut_data_7_sva_10[9:0]), {and_2391_cse , and_2392_cse , or_4705_cse
          , asn_1233});
      chn_mul_out_rsci_d_355_353 <= MUX1HOT_v_3_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_46_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_9_12_10_1, (MulIn_data_sva_536[243:241]),
          (MulOut_data_7_sva_10[12:10]), {and_2391_cse , and_2392_cse , or_4705_cse
          , asn_1233});
      chn_mul_out_rsci_d_365_356 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_23_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_9_22_13_1, (MulIn_data_sva_536[253:244]),
          (MulOut_data_7_sva_10[22:13]), {and_2391_cse , and_2392_cse , or_4705_cse
          , asn_1233});
      chn_mul_out_rsci_d_369_366 <= MUX1HOT_v_4_4_2((FpMul_8U_23U_FpMul_8U_23U_and_116_nl),
          reg_FpMul_8U_23U_p_expo_8_2_itm, (MulIn_data_sva_536[257:254]), (MulOut_data_7_sva_10[26:23]),
          {and_2383_cse , and_2384_cse , or_4705_cse , asn_1233});
      chn_mul_out_rsci_d_371_370 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_118_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_9_1_0_1, (MulIn_data_sva_536[259:258]),
          (MulOut_data_7_sva_10[28:27]), {and_2383_cse , and_2384_cse , or_4705_cse
          , asn_1233});
      chn_mul_out_rsci_d_373_372 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_117_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_9_3_2_1, (MulIn_data_sva_536[261:260]),
          (MulOut_data_7_sva_10[30:29]), {and_2383_cse , and_2384_cse , or_4705_cse
          , asn_1233});
      chn_mul_out_rsci_d_391_374 <= MUX1HOT_v_18_3_2(({{17{FpMul_8U_23U_mux_124_itm_4}},
          FpMul_8U_23U_mux_124_itm_4}), (signext_18_2(MulIn_data_sva_536[263:262])),
          (MulOut_data_7_sva_10[48:31]), {and_75_ssc , or_7_ssc , asn_1233});
      chn_mul_out_rsci_d_401_392 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_49_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_9_9_0_1, (MulIn_data_sva_536[273:264]),
          (MulOut_data_8_sva_10[9:0]), {and_2376_cse , and_2377_cse , or_4701_cse
          , asn_1243});
      chn_mul_out_rsci_d_404_402 <= MUX1HOT_v_3_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_48_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_9_12_10_1, (MulIn_data_sva_536[276:274]),
          (MulOut_data_8_sva_10[12:10]), {and_2376_cse , and_2377_cse , or_4701_cse
          , asn_1243});
      chn_mul_out_rsci_d_414_405 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_24_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_9_22_13_1, (MulIn_data_sva_536[286:277]),
          (MulOut_data_8_sva_10[22:13]), {and_2376_cse , and_2377_cse , or_4701_cse
          , asn_1243});
      chn_mul_out_rsci_d_418_415 <= MUX1HOT_v_4_4_2((FpMul_8U_23U_FpMul_8U_23U_and_119_nl),
          reg_FpMul_8U_23U_p_expo_9_2_itm, (MulIn_data_sva_536[290:287]), (MulOut_data_8_sva_10[26:23]),
          {and_2368_cse , and_2369_cse , or_4701_cse , asn_1243});
      chn_mul_out_rsci_d_420_419 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_121_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_9_1_0_1, (MulIn_data_sva_536[292:291]),
          (MulOut_data_8_sva_10[28:27]), {and_2368_cse , and_2369_cse , or_4701_cse
          , asn_1243});
      chn_mul_out_rsci_d_422_421 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_120_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_9_3_2_1, (MulIn_data_sva_536[294:293]),
          (MulOut_data_8_sva_10[30:29]), {and_2368_cse , and_2369_cse , or_4701_cse
          , asn_1243});
      chn_mul_out_rsci_d_440_423 <= MUX1HOT_v_18_3_2(({{17{FpMul_8U_23U_mux_140_itm_4}},
          FpMul_8U_23U_mux_140_itm_4}), (signext_18_2(MulIn_data_sva_536[296:295])),
          (MulOut_data_8_sva_10[48:31]), {and_79_ssc , or_8_ssc , asn_1243});
      chn_mul_out_rsci_d_450_441 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_51_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_9_9_0_1, (MulIn_data_sva_536[306:297]),
          (MulOut_data_9_sva_10[9:0]), {and_2361_cse , and_2362_cse , or_4697_cse
          , asn_1253});
      chn_mul_out_rsci_d_453_451 <= MUX1HOT_v_3_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_50_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_9_12_10_1, (MulIn_data_sva_536[309:307]),
          (MulOut_data_9_sva_10[12:10]), {and_2361_cse , and_2362_cse , or_4697_cse
          , asn_1253});
      chn_mul_out_rsci_d_463_454 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_25_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_9_22_13_1, (MulIn_data_sva_536[319:310]),
          (MulOut_data_9_sva_10[22:13]), {and_2361_cse , and_2362_cse , or_4697_cse
          , asn_1253});
      chn_mul_out_rsci_d_467_464 <= MUX1HOT_v_4_4_2((FpMul_8U_23U_FpMul_8U_23U_and_122_nl),
          reg_FpMul_8U_23U_p_expo_10_2_itm, (MulIn_data_sva_536[323:320]), (MulOut_data_9_sva_10[26:23]),
          {and_2353_cse , and_2354_cse , or_4697_cse , asn_1253});
      chn_mul_out_rsci_d_469_468 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_124_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_9_1_0_1, (MulIn_data_sva_536[325:324]),
          (MulOut_data_9_sva_10[28:27]), {and_2353_cse , and_2354_cse , or_4697_cse
          , asn_1253});
      chn_mul_out_rsci_d_471_470 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_123_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_9_3_2_1, (MulIn_data_sva_536[327:326]),
          (MulOut_data_9_sva_10[30:29]), {and_2353_cse , and_2354_cse , or_4697_cse
          , asn_1253});
      chn_mul_out_rsci_d_489_472 <= MUX1HOT_v_18_3_2(({{17{FpMul_8U_23U_mux_156_itm_4}},
          FpMul_8U_23U_mux_156_itm_4}), (signext_18_2(MulIn_data_sva_536[329:328])),
          (MulOut_data_9_sva_10[48:31]), {and_83_ssc , or_9_ssc , asn_1253});
      chn_mul_out_rsci_d_499_490 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_53_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_9_9_0_1, (MulIn_data_sva_536[339:330]),
          (MulOut_data_10_sva_10[9:0]), {and_2346_cse , and_2347_cse , or_4693_cse
          , asn_1263});
      chn_mul_out_rsci_d_502_500 <= MUX1HOT_v_3_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_52_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_9_12_10_1, (MulIn_data_sva_536[342:340]),
          (MulOut_data_10_sva_10[12:10]), {and_2346_cse , and_2347_cse , or_4693_cse
          , asn_1263});
      chn_mul_out_rsci_d_512_503 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_26_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_9_22_13_1, (MulIn_data_sva_536[352:343]),
          (MulOut_data_10_sva_10[22:13]), {and_2346_cse , and_2347_cse , or_4693_cse
          , asn_1263});
      chn_mul_out_rsci_d_516_513 <= MUX1HOT_v_4_4_2((FpMul_8U_23U_FpMul_8U_23U_and_125_nl),
          reg_FpMul_8U_23U_p_expo_11_2_itm, (MulIn_data_sva_536[356:353]), (MulOut_data_10_sva_10[26:23]),
          {and_2338_cse , and_2339_cse , or_4693_cse , asn_1263});
      chn_mul_out_rsci_d_518_517 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_127_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_9_1_0_1, (MulIn_data_sva_536[358:357]),
          (MulOut_data_10_sva_10[28:27]), {and_2338_cse , and_2339_cse , or_4693_cse
          , asn_1263});
      chn_mul_out_rsci_d_520_519 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_126_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_9_3_2_1, (MulIn_data_sva_536[360:359]),
          (MulOut_data_10_sva_10[30:29]), {and_2338_cse , and_2339_cse , or_4693_cse
          , asn_1263});
      chn_mul_out_rsci_d_538_521 <= MUX1HOT_v_18_3_2(({{17{FpMul_8U_23U_mux_172_itm_4}},
          FpMul_8U_23U_mux_172_itm_4}), (signext_18_2(MulIn_data_sva_536[362:361])),
          (MulOut_data_10_sva_10[48:31]), {and_87_ssc , or_10_ssc , asn_1263});
      chn_mul_out_rsci_d_548_539 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_55_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_9_9_0_1, (MulIn_data_sva_536[372:363]),
          (MulOut_data_11_sva_10[9:0]), {and_2331_cse , and_2332_cse , or_4689_cse
          , asn_1273});
      chn_mul_out_rsci_d_551_549 <= MUX1HOT_v_3_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_54_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_9_12_10_1, (MulIn_data_sva_536[375:373]),
          (MulOut_data_11_sva_10[12:10]), {and_2331_cse , and_2332_cse , or_4689_cse
          , asn_1273});
      chn_mul_out_rsci_d_561_552 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_27_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_9_22_13_1, (MulIn_data_sva_536[385:376]),
          (MulOut_data_11_sva_10[22:13]), {and_2331_cse , and_2332_cse , or_4689_cse
          , asn_1273});
      chn_mul_out_rsci_d_565_562 <= MUX1HOT_v_4_4_2((FpMul_8U_23U_FpMul_8U_23U_and_128_nl),
          reg_FpMul_8U_23U_p_expo_12_2_itm, (MulIn_data_sva_536[389:386]), (MulOut_data_11_sva_10[26:23]),
          {and_2323_cse , and_2324_cse , or_4689_cse , asn_1273});
      chn_mul_out_rsci_d_567_566 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_130_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_9_1_0_1, (MulIn_data_sva_536[391:390]),
          (MulOut_data_11_sva_10[28:27]), {and_2323_cse , and_2324_cse , or_4689_cse
          , asn_1273});
      chn_mul_out_rsci_d_569_568 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_129_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_9_3_2_1, (MulIn_data_sva_536[393:392]),
          (MulOut_data_11_sva_10[30:29]), {and_2323_cse , and_2324_cse , or_4689_cse
          , asn_1273});
      chn_mul_out_rsci_d_587_570 <= MUX1HOT_v_18_3_2(({{17{FpMul_8U_23U_mux_188_itm_4}},
          FpMul_8U_23U_mux_188_itm_4}), (signext_18_2(MulIn_data_sva_536[395:394])),
          (MulOut_data_11_sva_10[48:31]), {and_91_ssc , or_11_ssc , asn_1273});
      chn_mul_out_rsci_d_597_588 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_57_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_9_9_0_1, (MulIn_data_sva_536[405:396]),
          (MulOut_data_12_sva_10[9:0]), {and_2316_cse , and_2317_cse , or_4685_cse
          , asn_1283});
      chn_mul_out_rsci_d_600_598 <= MUX1HOT_v_3_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_56_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_9_12_10_1, (MulIn_data_sva_536[408:406]),
          (MulOut_data_12_sva_10[12:10]), {and_2316_cse , and_2317_cse , or_4685_cse
          , asn_1283});
      chn_mul_out_rsci_d_610_601 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_28_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_9_22_13_1, (MulIn_data_sva_536[418:409]),
          (MulOut_data_12_sva_10[22:13]), {and_2316_cse , and_2317_cse , or_4685_cse
          , asn_1283});
      chn_mul_out_rsci_d_614_611 <= MUX1HOT_v_4_4_2((FpMul_8U_23U_FpMul_8U_23U_and_131_nl),
          reg_FpMul_8U_23U_p_expo_13_2_itm, (MulIn_data_sva_536[422:419]), (MulOut_data_12_sva_10[26:23]),
          {and_2308_cse , and_2309_cse , or_4685_cse , asn_1283});
      chn_mul_out_rsci_d_616_615 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_133_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_9_1_0_1, (MulIn_data_sva_536[424:423]),
          (MulOut_data_12_sva_10[28:27]), {and_2308_cse , and_2309_cse , or_4685_cse
          , asn_1283});
      chn_mul_out_rsci_d_618_617 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_132_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_9_3_2_1, (MulIn_data_sva_536[426:425]),
          (MulOut_data_12_sva_10[30:29]), {and_2308_cse , and_2309_cse , or_4685_cse
          , asn_1283});
      chn_mul_out_rsci_d_636_619 <= MUX1HOT_v_18_3_2(({{17{FpMul_8U_23U_mux_204_itm_4}},
          FpMul_8U_23U_mux_204_itm_4}), (signext_18_2(MulIn_data_sva_536[428:427])),
          (MulOut_data_12_sva_10[48:31]), {and_95_ssc , or_12_ssc , asn_1283});
      chn_mul_out_rsci_d_646_637 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_59_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_9_9_0_1, (MulIn_data_sva_536[438:429]),
          (MulOut_data_13_sva_10[9:0]), {and_2301_cse , and_2302_cse , or_4681_cse
          , asn_1293});
      chn_mul_out_rsci_d_649_647 <= MUX1HOT_v_3_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_58_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_9_12_10_1, (MulIn_data_sva_536[441:439]),
          (MulOut_data_13_sva_10[12:10]), {and_2301_cse , and_2302_cse , or_4681_cse
          , asn_1293});
      chn_mul_out_rsci_d_659_650 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_29_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_9_22_13_1, (MulIn_data_sva_536[451:442]),
          (MulOut_data_13_sva_10[22:13]), {and_2301_cse , and_2302_cse , or_4681_cse
          , asn_1293});
      chn_mul_out_rsci_d_663_660 <= MUX1HOT_v_4_4_2((FpMul_8U_23U_FpMul_8U_23U_and_134_nl),
          reg_FpMul_8U_23U_p_expo_14_2_itm, (MulIn_data_sva_536[455:452]), (MulOut_data_13_sva_10[26:23]),
          {and_2293_cse , and_2294_cse , or_4681_cse , asn_1293});
      chn_mul_out_rsci_d_665_664 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_136_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_9_1_0_1, (MulIn_data_sva_536[457:456]),
          (MulOut_data_13_sva_10[28:27]), {and_2293_cse , and_2294_cse , or_4681_cse
          , asn_1293});
      chn_mul_out_rsci_d_667_666 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_135_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_9_3_2_1, (MulIn_data_sva_536[459:458]),
          (MulOut_data_13_sva_10[30:29]), {and_2293_cse , and_2294_cse , or_4681_cse
          , asn_1293});
      chn_mul_out_rsci_d_685_668 <= MUX1HOT_v_18_3_2(({{17{FpMul_8U_23U_mux_220_itm_4}},
          FpMul_8U_23U_mux_220_itm_4}), (signext_18_2(MulIn_data_sva_536[461:460])),
          (MulOut_data_13_sva_10[48:31]), {and_99_ssc , or_13_ssc , asn_1293});
      chn_mul_out_rsci_d_695_686 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_61_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_9_9_0_1, (MulIn_data_sva_536[471:462]),
          (MulOut_data_14_sva_10[9:0]), {and_2286_cse , and_2287_cse , or_4677_cse
          , asn_1303});
      chn_mul_out_rsci_d_698_696 <= MUX1HOT_v_3_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_60_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_9_12_10_1, (MulIn_data_sva_536[474:472]),
          (MulOut_data_14_sva_10[12:10]), {and_2286_cse , and_2287_cse , or_4677_cse
          , asn_1303});
      chn_mul_out_rsci_d_708_699 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_30_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_9_22_13_1, (MulIn_data_sva_536[484:475]),
          (MulOut_data_14_sva_10[22:13]), {and_2286_cse , and_2287_cse , or_4677_cse
          , asn_1303});
      chn_mul_out_rsci_d_712_709 <= MUX1HOT_v_4_4_2((FpMul_8U_23U_FpMul_8U_23U_and_137_nl),
          reg_FpMul_8U_23U_p_expo_15_2_itm, (MulIn_data_sva_536[488:485]), (MulOut_data_14_sva_10[26:23]),
          {and_2278_cse , and_2279_cse , or_4677_cse , asn_1303});
      chn_mul_out_rsci_d_714_713 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_139_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_9_1_0_1, (MulIn_data_sva_536[490:489]),
          (MulOut_data_14_sva_10[28:27]), {and_2278_cse , and_2279_cse , or_4677_cse
          , asn_1303});
      chn_mul_out_rsci_d_716_715 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_138_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_9_3_2_1, (MulIn_data_sva_536[492:491]),
          (MulOut_data_14_sva_10[30:29]), {and_2278_cse , and_2279_cse , or_4677_cse
          , asn_1303});
      chn_mul_out_rsci_d_734_717 <= MUX1HOT_v_18_3_2(({{17{FpMul_8U_23U_mux_236_itm_4}},
          FpMul_8U_23U_mux_236_itm_4}), (signext_18_2(MulIn_data_sva_536[494:493])),
          (MulOut_data_14_sva_10[48:31]), {and_103_ssc , or_14_ssc , asn_1303});
      chn_mul_out_rsci_d_744_735 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_63_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_9_9_0_1, (MulIn_data_sva_536[504:495]),
          (MulOut_data_15_sva_10[9:0]), {and_2271_cse , and_2272_cse , or_4673_cse
          , asn_1313});
      chn_mul_out_rsci_d_747_745 <= MUX1HOT_v_3_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_62_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_9_12_10_1, (MulIn_data_sva_536[507:505]),
          (MulOut_data_15_sva_10[12:10]), {and_2271_cse , and_2272_cse , or_4673_cse
          , asn_1313});
      chn_mul_out_rsci_d_757_748 <= MUX1HOT_v_10_4_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_31_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_9_22_13_1, (MulIn_data_sva_536[517:508]),
          (MulOut_data_15_sva_10[22:13]), {and_2271_cse , and_2272_cse , or_4673_cse
          , asn_1313});
      chn_mul_out_rsci_d_761_758 <= MUX1HOT_v_4_4_2((FpMul_8U_23U_FpMul_8U_23U_and_140_nl),
          reg_FpMul_8U_23U_p_expo_2_itm_1, (MulIn_data_sva_536[521:518]), (MulOut_data_15_sva_10[26:23]),
          {and_2263_cse , and_2264_cse , or_4673_cse , asn_1313});
      chn_mul_out_rsci_d_763_762 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_142_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_9_1_0_1, (MulIn_data_sva_536[523:522]),
          (MulOut_data_15_sva_10[28:27]), {and_2263_cse , and_2264_cse , or_4673_cse
          , asn_1313});
      chn_mul_out_rsci_d_765_764 <= MUX1HOT_v_2_4_2((FpMul_8U_23U_FpMul_8U_23U_and_141_nl),
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_9_3_2_1, (MulIn_data_sva_536[525:524]),
          (MulOut_data_15_sva_10[30:29]), {and_2263_cse , and_2264_cse , or_4673_cse
          , asn_1313});
      chn_mul_out_rsci_d_783_766 <= MUX1HOT_v_18_3_2(({{17{FpMul_8U_23U_mux_252_itm_4}},
          FpMul_8U_23U_mux_252_itm_4}), (signext_18_2(MulIn_data_sva_536[527:526])),
          (MulOut_data_15_sva_10[48:31]), {and_107_ssc , or_15_ssc , asn_1313});
      chn_mul_out_rsci_d_784 <= mul_loop_mul_else_land_1_lpi_1_dfm_10 & (~ io_read_cfg_mul_bypass_rsc_svs_8);
      chn_mul_out_rsci_d_785 <= mul_loop_mul_else_land_2_lpi_1_dfm_10 & (~ io_read_cfg_mul_bypass_rsc_svs_8);
      chn_mul_out_rsci_d_786 <= mul_loop_mul_else_land_3_lpi_1_dfm_10 & (~ io_read_cfg_mul_bypass_rsc_svs_8);
      chn_mul_out_rsci_d_787 <= mul_loop_mul_else_land_4_lpi_1_dfm_10 & (~ io_read_cfg_mul_bypass_rsc_svs_8);
      chn_mul_out_rsci_d_788 <= mul_loop_mul_else_land_5_lpi_1_dfm_10 & (~ io_read_cfg_mul_bypass_rsc_svs_8);
      chn_mul_out_rsci_d_789 <= mul_loop_mul_else_land_6_lpi_1_dfm_10 & (~ io_read_cfg_mul_bypass_rsc_svs_8);
      chn_mul_out_rsci_d_790 <= mul_loop_mul_else_land_7_lpi_1_dfm_10 & (~ io_read_cfg_mul_bypass_rsc_svs_8);
      chn_mul_out_rsci_d_791 <= mul_loop_mul_else_land_8_lpi_1_dfm_10 & (~ io_read_cfg_mul_bypass_rsc_svs_8);
      chn_mul_out_rsci_d_792 <= mul_loop_mul_else_land_9_lpi_1_dfm_10 & (~ io_read_cfg_mul_bypass_rsc_svs_8);
      chn_mul_out_rsci_d_793 <= mul_loop_mul_else_land_10_lpi_1_dfm_10 & (~ io_read_cfg_mul_bypass_rsc_svs_8);
      chn_mul_out_rsci_d_794 <= mul_loop_mul_else_land_11_lpi_1_dfm_10 & (~ io_read_cfg_mul_bypass_rsc_svs_8);
      chn_mul_out_rsci_d_795 <= mul_loop_mul_else_land_12_lpi_1_dfm_10 & (~ io_read_cfg_mul_bypass_rsc_svs_8);
      chn_mul_out_rsci_d_796 <= mul_loop_mul_else_land_13_lpi_1_dfm_10 & (~ io_read_cfg_mul_bypass_rsc_svs_8);
      chn_mul_out_rsci_d_797 <= mul_loop_mul_else_land_14_lpi_1_dfm_10 & (~ io_read_cfg_mul_bypass_rsc_svs_8);
      chn_mul_out_rsci_d_798 <= mul_loop_mul_else_land_15_lpi_1_dfm_10 & (~ io_read_cfg_mul_bypass_rsc_svs_8);
      chn_mul_out_rsci_d_799 <= mul_loop_mul_else_land_lpi_1_dfm_10 & (~ io_read_cfg_mul_bypass_rsc_svs_8);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_mul_out_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_56 | and_dcpl_58) ) begin
      reg_chn_mul_out_rsci_ld_core_psct_cse <= ~ and_dcpl_58;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_op_rsci_ld_core_psct <= 1'b0;
    end
    else if ( core_wen & (and_1647_cse | (or_dcpl_4 & and_dcpl_47 & (~ cfg_mul_bypass_rsci_d)
        & chn_mul_in_rsci_bawt & cfg_mul_src_rsci_d) | chn_mul_op_rsci_ld_core_psct_mx0c1)
        ) begin
      chn_mul_op_rsci_ld_core_psct <= ~ chn_mul_op_rsci_ld_core_psct_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_1 <= 1'b0;
    end
    else if ( core_wen & (or_tmp_3606 | main_stage_v_1_mx0c1) ) begin
      main_stage_v_1 <= ~ main_stage_v_1_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_5 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_31_cse & (~ (mux_19_nl))
        ) begin
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_5 <= MUX_s_1_2_2(IsNaN_8U_23U_land_1_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_1_lpi_1_dfm, and_dcpl_87);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_5 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_31_cse & (~ (mux_29_nl))
        ) begin
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_5 <= MUX_s_1_2_2(IsNaN_8U_23U_land_2_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_2_lpi_1_dfm, and_dcpl_87);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_5 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_31_cse & (~ (mux_39_nl))
        ) begin
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_5 <= MUX_s_1_2_2(IsNaN_8U_23U_land_3_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_3_lpi_1_dfm, and_dcpl_87);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_4_lpi_1_dfm_st_5 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_31_cse & (~ (mux_49_nl))
        ) begin
      IsNaN_8U_23U_land_4_lpi_1_dfm_st_5 <= MUX_s_1_2_2(IsNaN_8U_23U_land_4_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_4_lpi_1_dfm, and_dcpl_87);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_5_lpi_1_dfm_st_5 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_31_cse & (~ (mux_59_nl))
        ) begin
      IsNaN_8U_23U_land_5_lpi_1_dfm_st_5 <= MUX_s_1_2_2(IsNaN_8U_23U_land_5_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_5_lpi_1_dfm, and_dcpl_87);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_6_lpi_1_dfm_st_5 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_31_cse & (~ (mux_66_nl))
        ) begin
      IsNaN_8U_23U_land_6_lpi_1_dfm_st_5 <= MUX_s_1_2_2(IsNaN_8U_23U_land_6_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_6_lpi_1_dfm, and_dcpl_87);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_7_lpi_1_dfm_st_5 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_31_cse & (~ (mux_73_nl))
        ) begin
      IsNaN_8U_23U_land_7_lpi_1_dfm_st_5 <= MUX_s_1_2_2(IsNaN_8U_23U_land_7_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_7_lpi_1_dfm, and_dcpl_87);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_8_lpi_1_dfm_st_5 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_31_cse & (~ (mux_83_nl))
        ) begin
      IsNaN_8U_23U_land_8_lpi_1_dfm_st_5 <= MUX_s_1_2_2(IsNaN_8U_23U_land_8_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_8_lpi_1_dfm, and_dcpl_87);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_9_lpi_1_dfm_st_5 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_31_cse & (~ (mux_93_nl))
        ) begin
      IsNaN_8U_23U_land_9_lpi_1_dfm_st_5 <= MUX_s_1_2_2(IsNaN_8U_23U_land_9_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_9_lpi_1_dfm, and_dcpl_87);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_10_lpi_1_dfm_st_5 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_31_cse & (~ (mux_100_nl))
        ) begin
      IsNaN_8U_23U_land_10_lpi_1_dfm_st_5 <= MUX_s_1_2_2(IsNaN_8U_23U_land_10_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_10_lpi_1_dfm, and_dcpl_87);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_11_lpi_1_dfm_st_5 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_31_cse & (~ (mux_107_nl))
        ) begin
      IsNaN_8U_23U_land_11_lpi_1_dfm_st_5 <= MUX_s_1_2_2(IsNaN_8U_23U_land_11_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_11_lpi_1_dfm, and_dcpl_87);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_12_lpi_1_dfm_st_5 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_31_cse & (~ (mux_114_nl))
        ) begin
      IsNaN_8U_23U_land_12_lpi_1_dfm_st_5 <= MUX_s_1_2_2(IsNaN_8U_23U_land_12_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_12_lpi_1_dfm, and_dcpl_87);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_13_lpi_1_dfm_st_5 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_31_cse & (~ (mux_124_nl))
        ) begin
      IsNaN_8U_23U_land_13_lpi_1_dfm_st_5 <= MUX_s_1_2_2(IsNaN_8U_23U_land_13_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_13_lpi_1_dfm, and_dcpl_87);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_14_lpi_1_dfm_st_5 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_31_cse & (~ (mux_131_nl))
        ) begin
      IsNaN_8U_23U_land_14_lpi_1_dfm_st_5 <= MUX_s_1_2_2(IsNaN_8U_23U_land_14_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_14_lpi_1_dfm, and_dcpl_87);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_15_lpi_1_dfm_st_5 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_31_cse & (~ (mux_141_nl))
        ) begin
      IsNaN_8U_23U_land_15_lpi_1_dfm_st_5 <= MUX_s_1_2_2(IsNaN_8U_23U_land_15_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_15_lpi_1_dfm, and_dcpl_87);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_st_5 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_31_cse & (~ (mux_151_nl))
        ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_st_5 <= MUX_s_1_2_2(IsNaN_8U_23U_land_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_lpi_1_dfm, and_dcpl_87);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_if_land_lpi_1_dfm_st_5 <= 1'b0;
      mul_loop_mul_if_land_15_lpi_1_dfm_st_5 <= 1'b0;
      mul_loop_mul_if_land_14_lpi_1_dfm_st_5 <= 1'b0;
      mul_loop_mul_if_land_13_lpi_1_dfm_st_5 <= 1'b0;
      mul_loop_mul_if_land_12_lpi_1_dfm_st_5 <= 1'b0;
      mul_loop_mul_if_land_11_lpi_1_dfm_st_5 <= 1'b0;
      mul_loop_mul_if_land_10_lpi_1_dfm_st_5 <= 1'b0;
      mul_loop_mul_if_land_9_lpi_1_dfm_st_5 <= 1'b0;
      mul_loop_mul_if_land_8_lpi_1_dfm_st_5 <= 1'b0;
      mul_loop_mul_if_land_7_lpi_1_dfm_st_5 <= 1'b0;
      mul_loop_mul_if_land_6_lpi_1_dfm_st_5 <= 1'b0;
      mul_loop_mul_if_land_5_lpi_1_dfm_st_5 <= 1'b0;
      mul_loop_mul_if_land_4_lpi_1_dfm_st_5 <= 1'b0;
      mul_loop_mul_if_land_3_lpi_1_dfm_st_5 <= 1'b0;
      mul_loop_mul_if_land_2_lpi_1_dfm_st_5 <= 1'b0;
      mul_loop_mul_if_land_1_lpi_1_dfm_st_5 <= 1'b0;
    end
    else if ( mul_loop_mul_if_aelse_and_16_cse ) begin
      mul_loop_mul_if_land_lpi_1_dfm_st_5 <= MUX_s_1_2_2(nor_44_cse, mul_loop_mul_if_land_lpi_1_dfm_st,
          and_dcpl_87);
      mul_loop_mul_if_land_15_lpi_1_dfm_st_5 <= MUX_s_1_2_2(nor_42_cse, mul_loop_mul_if_land_15_lpi_1_dfm_st,
          and_dcpl_87);
      mul_loop_mul_if_land_14_lpi_1_dfm_st_5 <= MUX_s_1_2_2(nor_40_cse, mul_loop_mul_if_land_14_lpi_1_dfm_st,
          and_dcpl_87);
      mul_loop_mul_if_land_13_lpi_1_dfm_st_5 <= MUX_s_1_2_2(nor_39_cse, mul_loop_mul_if_land_13_lpi_1_dfm_st,
          and_dcpl_87);
      mul_loop_mul_if_land_12_lpi_1_dfm_st_5 <= MUX_s_1_2_2(nor_37_cse, mul_loop_mul_if_land_12_lpi_1_dfm_st,
          and_dcpl_87);
      mul_loop_mul_if_land_11_lpi_1_dfm_st_5 <= MUX_s_1_2_2(nor_36_cse, mul_loop_mul_if_land_11_lpi_1_dfm_st,
          and_dcpl_87);
      mul_loop_mul_if_land_10_lpi_1_dfm_st_5 <= MUX_s_1_2_2(nor_35_cse, mul_loop_mul_if_land_10_lpi_1_dfm_st,
          and_dcpl_87);
      mul_loop_mul_if_land_9_lpi_1_dfm_st_5 <= MUX_s_1_2_2(nor_34_cse, mul_loop_mul_if_land_9_lpi_1_dfm_st,
          and_dcpl_87);
      mul_loop_mul_if_land_8_lpi_1_dfm_st_5 <= MUX_s_1_2_2(nor_32_cse, mul_loop_mul_if_land_8_lpi_1_dfm_st,
          and_dcpl_87);
      mul_loop_mul_if_land_7_lpi_1_dfm_st_5 <= MUX_s_1_2_2(nor_30_cse, mul_loop_mul_if_land_7_lpi_1_dfm_st,
          and_dcpl_87);
      mul_loop_mul_if_land_6_lpi_1_dfm_st_5 <= MUX_s_1_2_2(nor_29_cse, mul_loop_mul_if_land_6_lpi_1_dfm_st,
          and_dcpl_87);
      mul_loop_mul_if_land_5_lpi_1_dfm_st_5 <= MUX_s_1_2_2(nor_28_cse, mul_loop_mul_if_land_5_lpi_1_dfm_st,
          and_dcpl_87);
      mul_loop_mul_if_land_4_lpi_1_dfm_st_5 <= MUX_s_1_2_2(nor_26_cse, mul_loop_mul_if_land_4_lpi_1_dfm_st,
          and_dcpl_87);
      mul_loop_mul_if_land_3_lpi_1_dfm_st_5 <= MUX_s_1_2_2(nor_25_cse, mul_loop_mul_if_land_3_lpi_1_dfm_st,
          and_dcpl_87);
      mul_loop_mul_if_land_2_lpi_1_dfm_st_5 <= MUX_s_1_2_2(nor_23_cse, mul_loop_mul_if_land_2_lpi_1_dfm_st,
          and_dcpl_87);
      mul_loop_mul_if_land_1_lpi_1_dfm_st_5 <= MUX_s_1_2_2(nor_21_cse, mul_loop_mul_if_land_1_lpi_1_dfm_st,
          and_dcpl_87);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_mul_op_1_sva_1 <= 16'b0;
      cfg_mul_src_1_sva_1 <= 1'b0;
    end
    else if ( cfg_mul_op_and_cse ) begin
      cfg_mul_op_1_sva_1 <= cfg_mul_op_rsci_d;
      cfg_mul_src_1_sva_1 <= cfg_mul_src_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_mul_src_1_sva_st_1 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_7 & and_dcpl_59 & (fsm_output[1])) | (or_dcpl_4
        & and_dcpl_47 & and_dcpl_59) | cfg_mul_src_1_sva_st_1_mx0c1) ) begin
      cfg_mul_src_1_sva_st_1 <= MUX_s_1_2_2(cfg_mul_src_rsci_d, cfg_mul_src_1_sva_st,
          cfg_mul_src_1_sva_st_1_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      io_read_cfg_mul_bypass_rsc_svs_st_1 <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_53 | and_dcpl_50 | (~ chn_mul_in_rsci_bawt)
        | (fsm_output[0]))) ) begin
      io_read_cfg_mul_bypass_rsc_svs_st_1 <= cfg_mul_bypass_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_75 | main_stage_v_2_mx0c1) ) begin
      main_stage_v_2 <= ~ main_stage_v_2_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_7_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_7_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_12_10_1 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_48_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_7_3_2_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_3_2_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_3_2, and_dcpl_102);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_7_1_0_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_1_0_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_1_0, and_dcpl_102);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3, and_dcpl_102);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_12_10_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_12_10, and_dcpl_102);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulIn_data_sva_534 <= 528'b0;
      io_read_cfg_mul_bypass_rsc_svs_st_5 <= 1'b0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_4_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_5_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_6_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_7_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_8_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_9_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_10_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_11_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_12_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_13_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_14_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_15_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_if_land_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_if_land_15_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_if_land_14_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_if_land_13_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_if_land_12_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_if_land_11_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_if_land_10_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_if_land_9_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_if_land_8_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_if_land_7_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_if_land_6_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_if_land_5_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_if_land_4_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_if_land_3_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_if_land_2_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_if_land_1_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_else_land_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_else_land_15_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_else_land_14_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_else_land_13_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_else_land_12_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_else_land_11_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_else_land_10_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_else_land_9_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_else_land_8_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_else_land_7_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_else_land_6_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_else_land_5_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_else_land_4_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_else_land_3_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_else_land_2_lpi_1_dfm_8 <= 1'b0;
      mul_loop_mul_else_land_1_lpi_1_dfm_8 <= 1'b0;
      io_read_cfg_mul_bypass_rsc_svs_6 <= 1'b0;
    end
    else if ( MulIn_data_and_cse ) begin
      MulIn_data_sva_534 <= MulIn_data_sva_533;
      io_read_cfg_mul_bypass_rsc_svs_st_5 <= io_read_cfg_mul_bypass_rsc_svs_st_1;
      IsNaN_8U_23U_land_1_lpi_1_dfm_9 <= IsNaN_8U_23U_land_1_lpi_1_dfm_8;
      IsNaN_8U_23U_land_2_lpi_1_dfm_9 <= IsNaN_8U_23U_land_2_lpi_1_dfm_8;
      IsNaN_8U_23U_land_3_lpi_1_dfm_9 <= IsNaN_8U_23U_land_3_lpi_1_dfm_8;
      IsNaN_8U_23U_land_4_lpi_1_dfm_9 <= IsNaN_8U_23U_land_4_lpi_1_dfm_8;
      IsNaN_8U_23U_land_5_lpi_1_dfm_9 <= IsNaN_8U_23U_land_5_lpi_1_dfm_8;
      IsNaN_8U_23U_land_6_lpi_1_dfm_9 <= IsNaN_8U_23U_land_6_lpi_1_dfm_8;
      IsNaN_8U_23U_land_7_lpi_1_dfm_9 <= IsNaN_8U_23U_land_7_lpi_1_dfm_8;
      IsNaN_8U_23U_land_8_lpi_1_dfm_9 <= IsNaN_8U_23U_land_8_lpi_1_dfm_8;
      IsNaN_8U_23U_land_9_lpi_1_dfm_9 <= IsNaN_8U_23U_land_9_lpi_1_dfm_8;
      IsNaN_8U_23U_land_10_lpi_1_dfm_9 <= IsNaN_8U_23U_land_10_lpi_1_dfm_8;
      IsNaN_8U_23U_land_11_lpi_1_dfm_9 <= IsNaN_8U_23U_land_11_lpi_1_dfm_8;
      IsNaN_8U_23U_land_12_lpi_1_dfm_9 <= IsNaN_8U_23U_land_12_lpi_1_dfm_8;
      IsNaN_8U_23U_land_13_lpi_1_dfm_9 <= IsNaN_8U_23U_land_13_lpi_1_dfm_8;
      IsNaN_8U_23U_land_14_lpi_1_dfm_9 <= IsNaN_8U_23U_land_14_lpi_1_dfm_8;
      IsNaN_8U_23U_land_15_lpi_1_dfm_9 <= IsNaN_8U_23U_land_15_lpi_1_dfm_8;
      IsNaN_8U_23U_land_lpi_1_dfm_9 <= IsNaN_8U_23U_land_lpi_1_dfm_8;
      mul_loop_mul_if_land_lpi_1_dfm_8 <= mul_loop_mul_if_land_lpi_1_dfm_7;
      mul_loop_mul_if_land_15_lpi_1_dfm_8 <= mul_loop_mul_if_land_15_lpi_1_dfm_7;
      mul_loop_mul_if_land_14_lpi_1_dfm_8 <= mul_loop_mul_if_land_14_lpi_1_dfm_7;
      mul_loop_mul_if_land_13_lpi_1_dfm_8 <= mul_loop_mul_if_land_13_lpi_1_dfm_7;
      mul_loop_mul_if_land_12_lpi_1_dfm_8 <= mul_loop_mul_if_land_12_lpi_1_dfm_7;
      mul_loop_mul_if_land_11_lpi_1_dfm_8 <= mul_loop_mul_if_land_11_lpi_1_dfm_7;
      mul_loop_mul_if_land_10_lpi_1_dfm_8 <= mul_loop_mul_if_land_10_lpi_1_dfm_7;
      mul_loop_mul_if_land_9_lpi_1_dfm_8 <= mul_loop_mul_if_land_9_lpi_1_dfm_7;
      mul_loop_mul_if_land_8_lpi_1_dfm_8 <= mul_loop_mul_if_land_8_lpi_1_dfm_7;
      mul_loop_mul_if_land_7_lpi_1_dfm_8 <= mul_loop_mul_if_land_7_lpi_1_dfm_7;
      mul_loop_mul_if_land_6_lpi_1_dfm_8 <= mul_loop_mul_if_land_6_lpi_1_dfm_7;
      mul_loop_mul_if_land_5_lpi_1_dfm_8 <= mul_loop_mul_if_land_5_lpi_1_dfm_7;
      mul_loop_mul_if_land_4_lpi_1_dfm_8 <= mul_loop_mul_if_land_4_lpi_1_dfm_7;
      mul_loop_mul_if_land_3_lpi_1_dfm_8 <= mul_loop_mul_if_land_3_lpi_1_dfm_7;
      mul_loop_mul_if_land_2_lpi_1_dfm_8 <= mul_loop_mul_if_land_2_lpi_1_dfm_7;
      mul_loop_mul_if_land_1_lpi_1_dfm_8 <= mul_loop_mul_if_land_1_lpi_1_dfm_7;
      mul_loop_mul_else_land_lpi_1_dfm_8 <= mul_loop_mul_else_land_lpi_1_dfm_7;
      mul_loop_mul_else_land_15_lpi_1_dfm_8 <= mul_loop_mul_else_land_15_lpi_1_dfm_7;
      mul_loop_mul_else_land_14_lpi_1_dfm_8 <= mul_loop_mul_else_land_14_lpi_1_dfm_7;
      mul_loop_mul_else_land_13_lpi_1_dfm_8 <= mul_loop_mul_else_land_13_lpi_1_dfm_7;
      mul_loop_mul_else_land_12_lpi_1_dfm_8 <= mul_loop_mul_else_land_12_lpi_1_dfm_7;
      mul_loop_mul_else_land_11_lpi_1_dfm_8 <= mul_loop_mul_else_land_11_lpi_1_dfm_7;
      mul_loop_mul_else_land_10_lpi_1_dfm_8 <= mul_loop_mul_else_land_10_lpi_1_dfm_7;
      mul_loop_mul_else_land_9_lpi_1_dfm_8 <= mul_loop_mul_else_land_9_lpi_1_dfm_7;
      mul_loop_mul_else_land_8_lpi_1_dfm_8 <= mul_loop_mul_else_land_8_lpi_1_dfm_7;
      mul_loop_mul_else_land_7_lpi_1_dfm_8 <= mul_loop_mul_else_land_7_lpi_1_dfm_7;
      mul_loop_mul_else_land_6_lpi_1_dfm_8 <= mul_loop_mul_else_land_6_lpi_1_dfm_7;
      mul_loop_mul_else_land_5_lpi_1_dfm_8 <= mul_loop_mul_else_land_5_lpi_1_dfm_7;
      mul_loop_mul_else_land_4_lpi_1_dfm_8 <= mul_loop_mul_else_land_4_lpi_1_dfm_7;
      mul_loop_mul_else_land_3_lpi_1_dfm_8 <= mul_loop_mul_else_land_3_lpi_1_dfm_7;
      mul_loop_mul_else_land_2_lpi_1_dfm_8 <= mul_loop_mul_else_land_2_lpi_1_dfm_7;
      mul_loop_mul_else_land_1_lpi_1_dfm_8 <= mul_loop_mul_else_land_1_lpi_1_dfm_7;
      io_read_cfg_mul_bypass_rsc_svs_6 <= io_read_cfg_mul_bypass_rsc_svs_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_lor_3_lpi_1_dfm_4_cse <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_156_itm)
        ) begin
      reg_FpMul_8U_23U_lor_3_lpi_1_dfm_4_cse <= MUX_s_1_2_2(FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_tmp,
          FpMul_8U_23U_lor_3_lpi_1_dfm_st, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_7_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_7_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_12_10_1 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_51_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_7_3_2_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_3_2_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_3_2, and_dcpl_108);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_7_1_0_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_1_0_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_1_0, and_dcpl_108);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3, and_dcpl_108);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_12_10_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_12_10, and_dcpl_108);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_lor_4_lpi_1_dfm_4_cse <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_157_itm)
        ) begin
      reg_FpMul_8U_23U_lor_4_lpi_1_dfm_4_cse <= MUX_s_1_2_2(FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_2_tmp,
          FpMul_8U_23U_lor_4_lpi_1_dfm_st, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_7_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_7_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_12_10_1 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_54_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_7_3_2_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_3_2_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_3_2, and_dcpl_112);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_7_1_0_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_1_0_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_1_0, and_dcpl_112);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3, and_dcpl_112);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_12_10_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_12_10, and_dcpl_112);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_lor_5_lpi_1_dfm_4_cse <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_158_itm)
        ) begin
      reg_FpMul_8U_23U_lor_5_lpi_1_dfm_4_cse <= MUX_s_1_2_2(FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_4_tmp,
          FpMul_8U_23U_lor_5_lpi_1_dfm_st, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_7_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_7_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_12_10_1 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_57_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_7_3_2_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_3_2_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_3_2, and_dcpl_116);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_7_1_0_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_1_0_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_1_0, and_dcpl_116);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3, and_dcpl_116);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_12_10_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_12_10, and_dcpl_116);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_lor_6_lpi_1_dfm_4_cse <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_159_itm)
        ) begin
      reg_FpMul_8U_23U_lor_6_lpi_1_dfm_4_cse <= MUX_s_1_2_2(FpMul_8U_23U_lor_6_lpi_1_dfm_mx0w0,
          FpMul_8U_23U_lor_6_lpi_1_dfm_st, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_7_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_7_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_12_10_1 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_60_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_7_3_2_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_3_2_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_3_2, and_dcpl_120);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_7_1_0_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_1_0_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_1_0, and_dcpl_120);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3, and_dcpl_120);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_12_10_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_12_10, and_dcpl_120);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_lor_7_lpi_1_dfm_4_cse <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_160_itm)
        ) begin
      reg_FpMul_8U_23U_lor_7_lpi_1_dfm_4_cse <= MUX_s_1_2_2(FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_8_tmp,
          FpMul_8U_23U_lor_7_lpi_1_dfm_st, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_7_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_7_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_12_10_1 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_63_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_7_3_2_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_3_2_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_3_2, and_dcpl_124);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_7_1_0_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_1_0_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_1_0, and_dcpl_124);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3, and_dcpl_124);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_12_10_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_12_10, and_dcpl_124);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_lor_8_lpi_1_dfm_4_cse <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_161_itm)
        ) begin
      reg_FpMul_8U_23U_lor_8_lpi_1_dfm_4_cse <= MUX_s_1_2_2(FpMul_8U_23U_lor_8_lpi_1_dfm_mx0w0,
          FpMul_8U_23U_lor_8_lpi_1_dfm_st, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_7_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_7_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_12_10_1 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_66_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_7_3_2_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_3_2_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_3_2, and_dcpl_128);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_7_1_0_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_1_0_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_1_0, and_dcpl_128);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3, and_dcpl_128);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_12_10_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_12_10, and_dcpl_128);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_lor_9_lpi_1_dfm_4_cse <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_162_itm)
        ) begin
      reg_FpMul_8U_23U_lor_9_lpi_1_dfm_4_cse <= MUX_s_1_2_2(FpMul_8U_23U_lor_9_lpi_1_dfm_mx0w0,
          FpMul_8U_23U_lor_9_lpi_1_dfm_st, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_7_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_7_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_12_10_1 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_69_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_7_3_2_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_3_2_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_3_2, and_dcpl_132);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_7_1_0_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_1_0_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_1_0, and_dcpl_132);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3, and_dcpl_132);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_12_10_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_12_10, and_dcpl_132);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_lor_10_lpi_1_dfm_4_cse <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_163_itm)
        ) begin
      reg_FpMul_8U_23U_lor_10_lpi_1_dfm_4_cse <= MUX_s_1_2_2(FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_14_tmp,
          FpMul_8U_23U_lor_10_lpi_1_dfm_st, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_7_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_7_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_12_10_1 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_72_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_7_3_2_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_3_2_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_3_2, and_dcpl_136);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_7_1_0_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_1_0_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_1_0, and_dcpl_136);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3, and_dcpl_136);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_12_10_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_12_10, and_dcpl_136);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_lor_11_lpi_1_dfm_4_cse <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_164_itm)
        ) begin
      reg_FpMul_8U_23U_lor_11_lpi_1_dfm_4_cse <= MUX_s_1_2_2(FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_16_tmp,
          FpMul_8U_23U_lor_11_lpi_1_dfm_st, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_7_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_7_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_12_10_1 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_75_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_7_3_2_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_3_2_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_3_2, and_dcpl_140);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_7_1_0_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_1_0_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_1_0, and_dcpl_140);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3, and_dcpl_140);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_12_10_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_12_10, and_dcpl_140);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_lor_12_lpi_1_dfm_4_cse <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_165_itm)
        ) begin
      reg_FpMul_8U_23U_lor_12_lpi_1_dfm_4_cse <= MUX_s_1_2_2(FpMul_8U_23U_lor_12_lpi_1_dfm_mx0w0,
          FpMul_8U_23U_lor_12_lpi_1_dfm_st, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_7_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_7_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_12_10_1 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_78_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_7_3_2_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_3_2_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_3_2, and_dcpl_144);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_7_1_0_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_1_0_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_1_0, and_dcpl_144);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3, and_dcpl_144);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_12_10_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_12_10, and_dcpl_144);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_lor_13_lpi_1_dfm_4_cse <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_166_itm)
        ) begin
      reg_FpMul_8U_23U_lor_13_lpi_1_dfm_4_cse <= MUX_s_1_2_2(FpMul_8U_23U_lor_13_lpi_1_dfm_mx0w0,
          FpMul_8U_23U_lor_13_lpi_1_dfm_st, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_7_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_7_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_12_10_1 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_81_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_7_3_2_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_3_2_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_3_2, and_dcpl_148);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_7_1_0_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_1_0_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_1_0, and_dcpl_148);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3, and_dcpl_148);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_12_10_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_12_10, and_dcpl_148);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_lor_14_lpi_1_dfm_4_cse <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_167_itm)
        ) begin
      reg_FpMul_8U_23U_lor_14_lpi_1_dfm_4_cse <= MUX_s_1_2_2(FpMul_8U_23U_lor_14_lpi_1_dfm_mx0w0,
          FpMul_8U_23U_lor_14_lpi_1_dfm_st, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_7_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_7_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_12_10_1 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_84_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_7_3_2_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_3_2_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_3_2, and_dcpl_152);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_7_1_0_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_1_0_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_1_0, and_dcpl_152);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3, and_dcpl_152);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_12_10_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_12_10, and_dcpl_152);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_lor_15_lpi_1_dfm_4_cse <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_168_itm)
        ) begin
      reg_FpMul_8U_23U_lor_15_lpi_1_dfm_4_cse <= MUX_s_1_2_2(FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_24_tmp,
          FpMul_8U_23U_lor_15_lpi_1_dfm_st, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_7_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_7_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_12_10_1 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_87_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_7_3_2_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_3_2_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_3_2, and_dcpl_156);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_7_1_0_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_1_0_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_1_0, and_dcpl_156);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3, and_dcpl_156);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_12_10_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_12_10, and_dcpl_156);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_lor_16_lpi_1_dfm_4_cse <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_169_itm)
        ) begin
      reg_FpMul_8U_23U_lor_16_lpi_1_dfm_4_cse <= MUX_s_1_2_2(FpMul_8U_23U_lor_16_lpi_1_dfm_mx0w0,
          FpMul_8U_23U_lor_16_lpi_1_dfm_st, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_7_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_7_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_12_10_1 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_90_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_7_3_2_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_3_2_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_3_2, and_dcpl_160);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_7_1_0_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_1_0_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_1_0, and_dcpl_160);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3, and_dcpl_160);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_12_10_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_12_10, and_dcpl_160);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_lor_17_lpi_1_dfm_4_cse <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_170_itm)
        ) begin
      reg_FpMul_8U_23U_lor_17_lpi_1_dfm_4_cse <= MUX_s_1_2_2(FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_28_tmp,
          FpMul_8U_23U_lor_17_lpi_1_dfm_st, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_7_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_7_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_9 <= 4'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_12_10_1 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_93_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_7_3_2_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_3_2_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_3_2, and_dcpl_164);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_7_1_0_1 <= MUX_v_2_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_1_0_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_1_0, and_dcpl_164);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3, and_dcpl_164);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_12_10_1 <= MUX_v_3_2_2(FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_12_10_mx0w0,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_12_10, and_dcpl_164);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_lor_lpi_1_dfm_4_cse <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_171_itm)
        ) begin
      reg_FpMul_8U_23U_lor_lpi_1_dfm_4_cse <= MUX_s_1_2_2(FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_30_tmp,
          FpMul_8U_23U_lor_lpi_1_dfm_st, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_if_land_lpi_1_dfm_st_6 <= 1'b0;
      mul_loop_mul_if_land_15_lpi_1_dfm_st_6 <= 1'b0;
      mul_loop_mul_if_land_14_lpi_1_dfm_st_6 <= 1'b0;
      mul_loop_mul_if_land_13_lpi_1_dfm_st_6 <= 1'b0;
      mul_loop_mul_if_land_12_lpi_1_dfm_st_6 <= 1'b0;
      mul_loop_mul_if_land_11_lpi_1_dfm_st_6 <= 1'b0;
      mul_loop_mul_if_land_10_lpi_1_dfm_st_6 <= 1'b0;
      mul_loop_mul_if_land_9_lpi_1_dfm_st_6 <= 1'b0;
      mul_loop_mul_if_land_8_lpi_1_dfm_st_6 <= 1'b0;
      mul_loop_mul_if_land_7_lpi_1_dfm_st_6 <= 1'b0;
      mul_loop_mul_if_land_6_lpi_1_dfm_st_6 <= 1'b0;
      mul_loop_mul_if_land_5_lpi_1_dfm_st_6 <= 1'b0;
      mul_loop_mul_if_land_4_lpi_1_dfm_st_6 <= 1'b0;
      mul_loop_mul_if_land_3_lpi_1_dfm_st_6 <= 1'b0;
      mul_loop_mul_if_land_2_lpi_1_dfm_st_6 <= 1'b0;
      mul_loop_mul_if_land_1_lpi_1_dfm_st_6 <= 1'b0;
    end
    else if ( mul_loop_mul_if_aelse_and_32_cse ) begin
      mul_loop_mul_if_land_lpi_1_dfm_st_6 <= mul_loop_mul_if_land_lpi_1_dfm_st_5;
      mul_loop_mul_if_land_15_lpi_1_dfm_st_6 <= mul_loop_mul_if_land_15_lpi_1_dfm_st_5;
      mul_loop_mul_if_land_14_lpi_1_dfm_st_6 <= mul_loop_mul_if_land_14_lpi_1_dfm_st_5;
      mul_loop_mul_if_land_13_lpi_1_dfm_st_6 <= mul_loop_mul_if_land_13_lpi_1_dfm_st_5;
      mul_loop_mul_if_land_12_lpi_1_dfm_st_6 <= mul_loop_mul_if_land_12_lpi_1_dfm_st_5;
      mul_loop_mul_if_land_11_lpi_1_dfm_st_6 <= mul_loop_mul_if_land_11_lpi_1_dfm_st_5;
      mul_loop_mul_if_land_10_lpi_1_dfm_st_6 <= mul_loop_mul_if_land_10_lpi_1_dfm_st_5;
      mul_loop_mul_if_land_9_lpi_1_dfm_st_6 <= mul_loop_mul_if_land_9_lpi_1_dfm_st_5;
      mul_loop_mul_if_land_8_lpi_1_dfm_st_6 <= mul_loop_mul_if_land_8_lpi_1_dfm_st_5;
      mul_loop_mul_if_land_7_lpi_1_dfm_st_6 <= mul_loop_mul_if_land_7_lpi_1_dfm_st_5;
      mul_loop_mul_if_land_6_lpi_1_dfm_st_6 <= mul_loop_mul_if_land_6_lpi_1_dfm_st_5;
      mul_loop_mul_if_land_5_lpi_1_dfm_st_6 <= mul_loop_mul_if_land_5_lpi_1_dfm_st_5;
      mul_loop_mul_if_land_4_lpi_1_dfm_st_6 <= mul_loop_mul_if_land_4_lpi_1_dfm_st_5;
      mul_loop_mul_if_land_3_lpi_1_dfm_st_6 <= mul_loop_mul_if_land_3_lpi_1_dfm_st_5;
      mul_loop_mul_if_land_2_lpi_1_dfm_st_6 <= mul_loop_mul_if_land_2_lpi_1_dfm_st_5;
      mul_loop_mul_if_land_1_lpi_1_dfm_st_6 <= mul_loop_mul_if_land_1_lpi_1_dfm_st_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_95 | main_stage_v_3_mx0c1) ) begin
      main_stage_v_3 <= ~ main_stage_v_3_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_1_lpi_1_dfm_8 <= 1'b0;
      IsZero_8U_23U_1_land_1_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_32_cse ) begin
      IsZero_8U_23U_land_1_lpi_1_dfm_8 <= IsZero_8U_23U_land_1_lpi_1_dfm_5;
      IsZero_8U_23U_1_land_1_lpi_1_dfm_7 <= IsZero_8U_23U_1_land_1_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulIn_data_sva_535 <= 528'b0;
      io_read_cfg_mul_bypass_rsc_svs_st_6 <= 1'b0;
      mul_loop_mul_if_land_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_if_land_15_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_if_land_14_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_if_land_13_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_if_land_12_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_if_land_11_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_if_land_10_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_if_land_9_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_if_land_8_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_if_land_7_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_if_land_6_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_if_land_5_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_if_land_4_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_if_land_3_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_if_land_2_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_if_land_1_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_else_land_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_else_land_15_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_else_land_14_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_else_land_13_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_else_land_12_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_else_land_11_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_else_land_10_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_else_land_9_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_else_land_8_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_else_land_7_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_else_land_6_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_else_land_5_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_else_land_4_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_else_land_3_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_else_land_2_lpi_1_dfm_9 <= 1'b0;
      mul_loop_mul_else_land_1_lpi_1_dfm_9 <= 1'b0;
      io_read_cfg_mul_bypass_rsc_svs_7 <= 1'b0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_4_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_5_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_6_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_7_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_8_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_9_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_10_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_11_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_12_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_13_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_14_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_15_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_10 <= 1'b0;
    end
    else if ( MulIn_data_and_1_cse ) begin
      MulIn_data_sva_535 <= MulIn_data_sva_534;
      io_read_cfg_mul_bypass_rsc_svs_st_6 <= io_read_cfg_mul_bypass_rsc_svs_st_5;
      mul_loop_mul_if_land_lpi_1_dfm_9 <= mul_loop_mul_if_land_lpi_1_dfm_8;
      mul_loop_mul_if_land_15_lpi_1_dfm_9 <= mul_loop_mul_if_land_15_lpi_1_dfm_8;
      mul_loop_mul_if_land_14_lpi_1_dfm_9 <= mul_loop_mul_if_land_14_lpi_1_dfm_8;
      mul_loop_mul_if_land_13_lpi_1_dfm_9 <= mul_loop_mul_if_land_13_lpi_1_dfm_8;
      mul_loop_mul_if_land_12_lpi_1_dfm_9 <= mul_loop_mul_if_land_12_lpi_1_dfm_8;
      mul_loop_mul_if_land_11_lpi_1_dfm_9 <= mul_loop_mul_if_land_11_lpi_1_dfm_8;
      mul_loop_mul_if_land_10_lpi_1_dfm_9 <= mul_loop_mul_if_land_10_lpi_1_dfm_8;
      mul_loop_mul_if_land_9_lpi_1_dfm_9 <= mul_loop_mul_if_land_9_lpi_1_dfm_8;
      mul_loop_mul_if_land_8_lpi_1_dfm_9 <= mul_loop_mul_if_land_8_lpi_1_dfm_8;
      mul_loop_mul_if_land_7_lpi_1_dfm_9 <= mul_loop_mul_if_land_7_lpi_1_dfm_8;
      mul_loop_mul_if_land_6_lpi_1_dfm_9 <= mul_loop_mul_if_land_6_lpi_1_dfm_8;
      mul_loop_mul_if_land_5_lpi_1_dfm_9 <= mul_loop_mul_if_land_5_lpi_1_dfm_8;
      mul_loop_mul_if_land_4_lpi_1_dfm_9 <= mul_loop_mul_if_land_4_lpi_1_dfm_8;
      mul_loop_mul_if_land_3_lpi_1_dfm_9 <= mul_loop_mul_if_land_3_lpi_1_dfm_8;
      mul_loop_mul_if_land_2_lpi_1_dfm_9 <= mul_loop_mul_if_land_2_lpi_1_dfm_8;
      mul_loop_mul_if_land_1_lpi_1_dfm_9 <= mul_loop_mul_if_land_1_lpi_1_dfm_8;
      mul_loop_mul_else_land_lpi_1_dfm_9 <= mul_loop_mul_else_land_lpi_1_dfm_8;
      mul_loop_mul_else_land_15_lpi_1_dfm_9 <= mul_loop_mul_else_land_15_lpi_1_dfm_8;
      mul_loop_mul_else_land_14_lpi_1_dfm_9 <= mul_loop_mul_else_land_14_lpi_1_dfm_8;
      mul_loop_mul_else_land_13_lpi_1_dfm_9 <= mul_loop_mul_else_land_13_lpi_1_dfm_8;
      mul_loop_mul_else_land_12_lpi_1_dfm_9 <= mul_loop_mul_else_land_12_lpi_1_dfm_8;
      mul_loop_mul_else_land_11_lpi_1_dfm_9 <= mul_loop_mul_else_land_11_lpi_1_dfm_8;
      mul_loop_mul_else_land_10_lpi_1_dfm_9 <= mul_loop_mul_else_land_10_lpi_1_dfm_8;
      mul_loop_mul_else_land_9_lpi_1_dfm_9 <= mul_loop_mul_else_land_9_lpi_1_dfm_8;
      mul_loop_mul_else_land_8_lpi_1_dfm_9 <= mul_loop_mul_else_land_8_lpi_1_dfm_8;
      mul_loop_mul_else_land_7_lpi_1_dfm_9 <= mul_loop_mul_else_land_7_lpi_1_dfm_8;
      mul_loop_mul_else_land_6_lpi_1_dfm_9 <= mul_loop_mul_else_land_6_lpi_1_dfm_8;
      mul_loop_mul_else_land_5_lpi_1_dfm_9 <= mul_loop_mul_else_land_5_lpi_1_dfm_8;
      mul_loop_mul_else_land_4_lpi_1_dfm_9 <= mul_loop_mul_else_land_4_lpi_1_dfm_8;
      mul_loop_mul_else_land_3_lpi_1_dfm_9 <= mul_loop_mul_else_land_3_lpi_1_dfm_8;
      mul_loop_mul_else_land_2_lpi_1_dfm_9 <= mul_loop_mul_else_land_2_lpi_1_dfm_8;
      mul_loop_mul_else_land_1_lpi_1_dfm_9 <= mul_loop_mul_else_land_1_lpi_1_dfm_8;
      io_read_cfg_mul_bypass_rsc_svs_7 <= io_read_cfg_mul_bypass_rsc_svs_6;
      IsNaN_8U_23U_land_1_lpi_1_dfm_10 <= IsNaN_8U_23U_land_1_lpi_1_dfm_9;
      IsNaN_8U_23U_land_2_lpi_1_dfm_10 <= IsNaN_8U_23U_land_2_lpi_1_dfm_9;
      IsNaN_8U_23U_land_3_lpi_1_dfm_10 <= IsNaN_8U_23U_land_3_lpi_1_dfm_9;
      IsNaN_8U_23U_land_4_lpi_1_dfm_10 <= IsNaN_8U_23U_land_4_lpi_1_dfm_9;
      IsNaN_8U_23U_land_5_lpi_1_dfm_10 <= IsNaN_8U_23U_land_5_lpi_1_dfm_9;
      IsNaN_8U_23U_land_6_lpi_1_dfm_10 <= IsNaN_8U_23U_land_6_lpi_1_dfm_9;
      IsNaN_8U_23U_land_7_lpi_1_dfm_10 <= IsNaN_8U_23U_land_7_lpi_1_dfm_9;
      IsNaN_8U_23U_land_8_lpi_1_dfm_10 <= IsNaN_8U_23U_land_8_lpi_1_dfm_9;
      IsNaN_8U_23U_land_9_lpi_1_dfm_10 <= IsNaN_8U_23U_land_9_lpi_1_dfm_9;
      IsNaN_8U_23U_land_10_lpi_1_dfm_10 <= IsNaN_8U_23U_land_10_lpi_1_dfm_9;
      IsNaN_8U_23U_land_11_lpi_1_dfm_10 <= IsNaN_8U_23U_land_11_lpi_1_dfm_9;
      IsNaN_8U_23U_land_12_lpi_1_dfm_10 <= IsNaN_8U_23U_land_12_lpi_1_dfm_9;
      IsNaN_8U_23U_land_13_lpi_1_dfm_10 <= IsNaN_8U_23U_land_13_lpi_1_dfm_9;
      IsNaN_8U_23U_land_14_lpi_1_dfm_10 <= IsNaN_8U_23U_land_14_lpi_1_dfm_9;
      IsNaN_8U_23U_land_15_lpi_1_dfm_10 <= IsNaN_8U_23U_land_15_lpi_1_dfm_9;
      IsNaN_8U_23U_land_lpi_1_dfm_10 <= IsNaN_8U_23U_land_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_48_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_22_13_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_9_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_186_nl)
        ) begin
      mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= MUX_s_1_2_2(mul_loop_mul_1_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st,
          and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_18_lpi_1_dfm_st_3 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_187_itm)
        ) begin
      FpMul_8U_23U_lor_18_lpi_1_dfm_st_3 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_31_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_2_lpi_1_dfm_8 <= 1'b0;
      IsZero_8U_23U_1_land_2_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_33_cse ) begin
      IsZero_8U_23U_land_2_lpi_1_dfm_8 <= IsZero_8U_23U_land_2_lpi_1_dfm_5;
      IsZero_8U_23U_1_land_2_lpi_1_dfm_7 <= IsZero_8U_23U_1_land_2_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_51_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_22_13_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_9_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_201_nl))
        ) begin
      mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= MUX_s_1_2_2(mul_loop_mul_2_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st,
          and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_19_lpi_1_dfm_st_3 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_202_itm)
        ) begin
      FpMul_8U_23U_lor_19_lpi_1_dfm_st_3 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_30_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_3_lpi_1_dfm_8 <= 1'b0;
      IsZero_8U_23U_1_land_3_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_34_cse ) begin
      IsZero_8U_23U_land_3_lpi_1_dfm_8 <= IsZero_8U_23U_land_3_lpi_1_dfm_5;
      IsZero_8U_23U_1_land_3_lpi_1_dfm_7 <= IsZero_8U_23U_1_land_3_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_54_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_22_13_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_9_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_215_nl)
        ) begin
      mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= MUX_s_1_2_2(mul_loop_mul_3_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st,
          and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_20_lpi_1_dfm_st_3 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_216_itm)
        ) begin
      FpMul_8U_23U_lor_20_lpi_1_dfm_st_3 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_29_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_4_lpi_1_dfm_8 <= 1'b0;
      IsZero_8U_23U_1_land_4_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_35_cse ) begin
      IsZero_8U_23U_land_4_lpi_1_dfm_8 <= IsZero_8U_23U_land_4_lpi_1_dfm_5;
      IsZero_8U_23U_1_land_4_lpi_1_dfm_6 <= IsZero_8U_23U_1_land_4_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_57_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_22_13_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_9_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_229_nl)
        ) begin
      mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= MUX_s_1_2_2(mul_loop_mul_4_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st,
          and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_21_lpi_1_dfm_st_3 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_230_itm)
        ) begin
      FpMul_8U_23U_lor_21_lpi_1_dfm_st_3 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_28_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_5_lpi_1_dfm_8 <= 1'b0;
      IsZero_8U_23U_1_land_5_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_36_cse ) begin
      IsZero_8U_23U_land_5_lpi_1_dfm_8 <= IsZero_8U_23U_land_5_lpi_1_dfm_5;
      IsZero_8U_23U_1_land_5_lpi_1_dfm_7 <= IsZero_8U_23U_1_land_5_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_60_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_22_13_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_9_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_244_nl))
        ) begin
      mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= MUX_s_1_2_2(mul_loop_mul_5_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st,
          and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_22_lpi_1_dfm_st_3 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_245_itm)
        ) begin
      FpMul_8U_23U_lor_22_lpi_1_dfm_st_3 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_27_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_6_lpi_1_dfm_8 <= 1'b0;
      IsZero_8U_23U_1_land_6_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_37_cse ) begin
      IsZero_8U_23U_land_6_lpi_1_dfm_8 <= IsZero_8U_23U_land_6_lpi_1_dfm_5;
      IsZero_8U_23U_1_land_6_lpi_1_dfm_6 <= IsZero_8U_23U_1_land_6_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_63_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_22_13_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_9_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_258_nl)
        ) begin
      mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= MUX_s_1_2_2(mul_loop_mul_6_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st,
          and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_23_lpi_1_dfm_st_3 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_259_itm)
        ) begin
      FpMul_8U_23U_lor_23_lpi_1_dfm_st_3 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_26_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_7_lpi_1_dfm_8 <= 1'b0;
      IsZero_8U_23U_1_land_7_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_38_cse ) begin
      IsZero_8U_23U_land_7_lpi_1_dfm_8 <= IsZero_8U_23U_land_7_lpi_1_dfm_5;
      IsZero_8U_23U_1_land_7_lpi_1_dfm_6 <= IsZero_8U_23U_1_land_7_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_66_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_22_13_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_9_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_272_nl)
        ) begin
      mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= MUX_s_1_2_2(mul_loop_mul_7_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st,
          and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_24_lpi_1_dfm_st_3 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_273_itm)
        ) begin
      FpMul_8U_23U_lor_24_lpi_1_dfm_st_3 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_25_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_8_lpi_1_dfm_8 <= 1'b0;
      IsZero_8U_23U_1_land_8_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_39_cse ) begin
      IsZero_8U_23U_land_8_lpi_1_dfm_8 <= IsZero_8U_23U_land_8_lpi_1_dfm_5;
      IsZero_8U_23U_1_land_8_lpi_1_dfm_7 <= IsZero_8U_23U_1_land_8_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_69_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_22_13_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_9_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_287_nl))
        ) begin
      mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= MUX_s_1_2_2(mul_loop_mul_8_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st,
          and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_25_lpi_1_dfm_st_3 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_288_itm)
        ) begin
      FpMul_8U_23U_lor_25_lpi_1_dfm_st_3 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_24_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_9_lpi_1_dfm_8 <= 1'b0;
      IsZero_8U_23U_1_land_9_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_40_cse ) begin
      IsZero_8U_23U_land_9_lpi_1_dfm_8 <= IsZero_8U_23U_land_9_lpi_1_dfm_5;
      IsZero_8U_23U_1_land_9_lpi_1_dfm_7 <= IsZero_8U_23U_1_land_9_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_72_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_22_13_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_9_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_302_nl))
        ) begin
      mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= MUX_s_1_2_2(mul_loop_mul_9_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st,
          and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_26_lpi_1_dfm_st_3 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_303_itm)
        ) begin
      FpMul_8U_23U_lor_26_lpi_1_dfm_st_3 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_23_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_10_lpi_1_dfm_8 <= 1'b0;
      IsZero_8U_23U_1_land_10_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_41_cse ) begin
      IsZero_8U_23U_land_10_lpi_1_dfm_8 <= IsZero_8U_23U_land_10_lpi_1_dfm_5;
      IsZero_8U_23U_1_land_10_lpi_1_dfm_6 <= IsZero_8U_23U_1_land_10_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_75_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_22_13_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_9_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_317_nl))
        ) begin
      mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= MUX_s_1_2_2(mul_loop_mul_10_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st,
          and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_27_lpi_1_dfm_st_3 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_318_itm)
        ) begin
      FpMul_8U_23U_lor_27_lpi_1_dfm_st_3 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_22_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_11_lpi_1_dfm_8 <= 1'b0;
      IsZero_8U_23U_1_land_11_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_42_cse ) begin
      IsZero_8U_23U_land_11_lpi_1_dfm_8 <= IsZero_8U_23U_land_11_lpi_1_dfm_5;
      IsZero_8U_23U_1_land_11_lpi_1_dfm_6 <= IsZero_8U_23U_1_land_11_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_78_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_22_13_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_9_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_331_nl)
        ) begin
      mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= MUX_s_1_2_2(mul_loop_mul_11_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st,
          and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_28_lpi_1_dfm_st_3 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_332_itm)
        ) begin
      FpMul_8U_23U_lor_28_lpi_1_dfm_st_3 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_21_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_12_lpi_1_dfm_8 <= 1'b0;
      IsZero_8U_23U_1_land_12_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_43_cse ) begin
      IsZero_8U_23U_land_12_lpi_1_dfm_8 <= IsZero_8U_23U_land_12_lpi_1_dfm_5;
      IsZero_8U_23U_1_land_12_lpi_1_dfm_6 <= IsZero_8U_23U_1_land_12_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_81_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_22_13_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_9_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_345_nl)
        ) begin
      mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= MUX_s_1_2_2(mul_loop_mul_12_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st,
          and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_29_lpi_1_dfm_st_3 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_346_itm)
        ) begin
      FpMul_8U_23U_lor_29_lpi_1_dfm_st_3 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_20_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_13_lpi_1_dfm_8 <= 1'b0;
      IsZero_8U_23U_1_land_13_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_44_cse ) begin
      IsZero_8U_23U_land_13_lpi_1_dfm_8 <= IsZero_8U_23U_land_13_lpi_1_dfm_5;
      IsZero_8U_23U_1_land_13_lpi_1_dfm_7 <= IsZero_8U_23U_1_land_13_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_84_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_22_13_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_9_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_359_nl)
        ) begin
      mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= MUX_s_1_2_2(mul_loop_mul_13_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st,
          and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_30_lpi_1_dfm_st_3 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_360_itm)
        ) begin
      FpMul_8U_23U_lor_30_lpi_1_dfm_st_3 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_19_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_14_lpi_1_dfm_8 <= 1'b0;
      IsZero_8U_23U_1_land_14_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_45_cse ) begin
      IsZero_8U_23U_land_14_lpi_1_dfm_8 <= IsZero_8U_23U_land_14_lpi_1_dfm_5;
      IsZero_8U_23U_1_land_14_lpi_1_dfm_6 <= IsZero_8U_23U_1_land_14_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_87_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_22_13_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_9_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_373_nl)
        ) begin
      mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= MUX_s_1_2_2(mul_loop_mul_14_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st,
          and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_31_lpi_1_dfm_st_3 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_374_itm)
        ) begin
      FpMul_8U_23U_lor_31_lpi_1_dfm_st_3 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_18_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_15_lpi_1_dfm_8 <= 1'b0;
      IsZero_8U_23U_1_land_15_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_46_cse ) begin
      IsZero_8U_23U_land_15_lpi_1_dfm_8 <= IsZero_8U_23U_land_15_lpi_1_dfm_5;
      IsZero_8U_23U_1_land_15_lpi_1_dfm_7 <= IsZero_8U_23U_1_land_15_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_90_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_22_13_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_9_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_387_nl)
        ) begin
      mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= MUX_s_1_2_2(mul_loop_mul_15_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st,
          and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_32_lpi_1_dfm_st_3 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_388_itm)
        ) begin
      FpMul_8U_23U_lor_32_lpi_1_dfm_st_3 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_17_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_lpi_1_dfm_8 <= 1'b0;
      IsZero_8U_23U_1_land_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_47_cse ) begin
      IsZero_8U_23U_land_lpi_1_dfm_8 <= IsZero_8U_23U_land_lpi_1_dfm_5;
      IsZero_8U_23U_1_land_lpi_1_dfm_7 <= IsZero_8U_23U_1_land_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_93_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_22_13_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_9_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_402_nl))
        ) begin
      mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= MUX_s_1_2_2(mul_loop_mul_16_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st,
          and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_403_itm)
        ) begin
      FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_16_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_if_land_lpi_1_dfm_st_7 <= 1'b0;
      mul_loop_mul_if_land_15_lpi_1_dfm_st_7 <= 1'b0;
      mul_loop_mul_if_land_14_lpi_1_dfm_st_7 <= 1'b0;
      mul_loop_mul_if_land_13_lpi_1_dfm_st_7 <= 1'b0;
      mul_loop_mul_if_land_12_lpi_1_dfm_st_7 <= 1'b0;
      mul_loop_mul_if_land_11_lpi_1_dfm_st_7 <= 1'b0;
      mul_loop_mul_if_land_10_lpi_1_dfm_st_7 <= 1'b0;
      mul_loop_mul_if_land_9_lpi_1_dfm_st_7 <= 1'b0;
      mul_loop_mul_if_land_8_lpi_1_dfm_st_7 <= 1'b0;
      mul_loop_mul_if_land_7_lpi_1_dfm_st_7 <= 1'b0;
      mul_loop_mul_if_land_6_lpi_1_dfm_st_7 <= 1'b0;
      mul_loop_mul_if_land_5_lpi_1_dfm_st_7 <= 1'b0;
      mul_loop_mul_if_land_4_lpi_1_dfm_st_7 <= 1'b0;
      mul_loop_mul_if_land_3_lpi_1_dfm_st_7 <= 1'b0;
      mul_loop_mul_if_land_2_lpi_1_dfm_st_7 <= 1'b0;
      mul_loop_mul_if_land_1_lpi_1_dfm_st_7 <= 1'b0;
    end
    else if ( mul_loop_mul_if_aelse_and_48_cse ) begin
      mul_loop_mul_if_land_lpi_1_dfm_st_7 <= mul_loop_mul_if_land_lpi_1_dfm_st_6;
      mul_loop_mul_if_land_15_lpi_1_dfm_st_7 <= mul_loop_mul_if_land_15_lpi_1_dfm_st_6;
      mul_loop_mul_if_land_14_lpi_1_dfm_st_7 <= mul_loop_mul_if_land_14_lpi_1_dfm_st_6;
      mul_loop_mul_if_land_13_lpi_1_dfm_st_7 <= mul_loop_mul_if_land_13_lpi_1_dfm_st_6;
      mul_loop_mul_if_land_12_lpi_1_dfm_st_7 <= mul_loop_mul_if_land_12_lpi_1_dfm_st_6;
      mul_loop_mul_if_land_11_lpi_1_dfm_st_7 <= mul_loop_mul_if_land_11_lpi_1_dfm_st_6;
      mul_loop_mul_if_land_10_lpi_1_dfm_st_7 <= mul_loop_mul_if_land_10_lpi_1_dfm_st_6;
      mul_loop_mul_if_land_9_lpi_1_dfm_st_7 <= mul_loop_mul_if_land_9_lpi_1_dfm_st_6;
      mul_loop_mul_if_land_8_lpi_1_dfm_st_7 <= mul_loop_mul_if_land_8_lpi_1_dfm_st_6;
      mul_loop_mul_if_land_7_lpi_1_dfm_st_7 <= mul_loop_mul_if_land_7_lpi_1_dfm_st_6;
      mul_loop_mul_if_land_6_lpi_1_dfm_st_7 <= mul_loop_mul_if_land_6_lpi_1_dfm_st_6;
      mul_loop_mul_if_land_5_lpi_1_dfm_st_7 <= mul_loop_mul_if_land_5_lpi_1_dfm_st_6;
      mul_loop_mul_if_land_4_lpi_1_dfm_st_7 <= mul_loop_mul_if_land_4_lpi_1_dfm_st_6;
      mul_loop_mul_if_land_3_lpi_1_dfm_st_7 <= mul_loop_mul_if_land_3_lpi_1_dfm_st_6;
      mul_loop_mul_if_land_2_lpi_1_dfm_st_7 <= mul_loop_mul_if_land_2_lpi_1_dfm_st_6;
      mul_loop_mul_if_land_1_lpi_1_dfm_st_7 <= mul_loop_mul_if_land_1_lpi_1_dfm_st_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_4 <= 1'b0;
    end
    else if ( core_wen & ((or_309_cse & main_stage_v_3) | main_stage_v_4_mx0c1) )
        begin
      main_stage_v_4 <= ~ main_stage_v_4_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulIn_data_sva_536 <= 528'b0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_11 <= 1'b0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_11 <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_11 <= 1'b0;
      IsNaN_8U_23U_land_4_lpi_1_dfm_11 <= 1'b0;
      IsNaN_8U_23U_land_5_lpi_1_dfm_11 <= 1'b0;
      IsNaN_8U_23U_land_6_lpi_1_dfm_11 <= 1'b0;
      IsNaN_8U_23U_land_7_lpi_1_dfm_11 <= 1'b0;
      IsNaN_8U_23U_land_8_lpi_1_dfm_11 <= 1'b0;
      IsNaN_8U_23U_land_9_lpi_1_dfm_11 <= 1'b0;
      IsNaN_8U_23U_land_10_lpi_1_dfm_11 <= 1'b0;
      IsNaN_8U_23U_land_11_lpi_1_dfm_11 <= 1'b0;
      IsNaN_8U_23U_land_12_lpi_1_dfm_11 <= 1'b0;
      IsNaN_8U_23U_land_13_lpi_1_dfm_11 <= 1'b0;
      IsNaN_8U_23U_land_14_lpi_1_dfm_11 <= 1'b0;
      IsNaN_8U_23U_land_15_lpi_1_dfm_11 <= 1'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_11 <= 1'b0;
      mul_loop_mul_else_land_lpi_1_dfm_10 <= 1'b0;
      io_read_cfg_mul_bypass_rsc_svs_8 <= 1'b0;
      mul_loop_mul_else_land_1_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_if_land_1_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_else_land_15_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_else_land_2_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_if_land_2_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_else_land_14_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_else_land_3_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_if_land_3_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_else_land_13_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_else_land_4_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_if_land_4_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_else_land_12_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_else_land_5_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_if_land_5_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_else_land_11_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_else_land_6_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_if_land_6_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_else_land_10_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_else_land_7_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_if_land_7_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_else_land_9_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_else_land_8_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_if_land_8_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_if_land_9_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_if_land_10_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_if_land_11_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_if_land_12_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_if_land_13_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_if_land_14_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_if_land_15_lpi_1_dfm_10 <= 1'b0;
      mul_loop_mul_if_land_lpi_1_dfm_10 <= 1'b0;
      io_read_cfg_mul_bypass_rsc_svs_st_7 <= 1'b0;
    end
    else if ( MulIn_data_and_2_cse ) begin
      MulIn_data_sva_536 <= MulIn_data_sva_535;
      IsNaN_8U_23U_land_1_lpi_1_dfm_11 <= IsNaN_8U_23U_land_1_lpi_1_dfm_10;
      IsNaN_8U_23U_land_2_lpi_1_dfm_11 <= IsNaN_8U_23U_land_2_lpi_1_dfm_10;
      IsNaN_8U_23U_land_3_lpi_1_dfm_11 <= IsNaN_8U_23U_land_3_lpi_1_dfm_10;
      IsNaN_8U_23U_land_4_lpi_1_dfm_11 <= IsNaN_8U_23U_land_4_lpi_1_dfm_10;
      IsNaN_8U_23U_land_5_lpi_1_dfm_11 <= IsNaN_8U_23U_land_5_lpi_1_dfm_10;
      IsNaN_8U_23U_land_6_lpi_1_dfm_11 <= IsNaN_8U_23U_land_6_lpi_1_dfm_10;
      IsNaN_8U_23U_land_7_lpi_1_dfm_11 <= IsNaN_8U_23U_land_7_lpi_1_dfm_10;
      IsNaN_8U_23U_land_8_lpi_1_dfm_11 <= IsNaN_8U_23U_land_8_lpi_1_dfm_10;
      IsNaN_8U_23U_land_9_lpi_1_dfm_11 <= IsNaN_8U_23U_land_9_lpi_1_dfm_10;
      IsNaN_8U_23U_land_10_lpi_1_dfm_11 <= IsNaN_8U_23U_land_10_lpi_1_dfm_10;
      IsNaN_8U_23U_land_11_lpi_1_dfm_11 <= IsNaN_8U_23U_land_11_lpi_1_dfm_10;
      IsNaN_8U_23U_land_12_lpi_1_dfm_11 <= IsNaN_8U_23U_land_12_lpi_1_dfm_10;
      IsNaN_8U_23U_land_13_lpi_1_dfm_11 <= IsNaN_8U_23U_land_13_lpi_1_dfm_10;
      IsNaN_8U_23U_land_14_lpi_1_dfm_11 <= IsNaN_8U_23U_land_14_lpi_1_dfm_10;
      IsNaN_8U_23U_land_15_lpi_1_dfm_11 <= IsNaN_8U_23U_land_15_lpi_1_dfm_10;
      IsNaN_8U_23U_land_lpi_1_dfm_11 <= IsNaN_8U_23U_land_lpi_1_dfm_10;
      mul_loop_mul_else_land_lpi_1_dfm_10 <= mul_loop_mul_else_land_lpi_1_dfm_9;
      io_read_cfg_mul_bypass_rsc_svs_8 <= io_read_cfg_mul_bypass_rsc_svs_7;
      mul_loop_mul_else_land_1_lpi_1_dfm_10 <= mul_loop_mul_else_land_1_lpi_1_dfm_9;
      mul_loop_mul_if_land_1_lpi_1_dfm_10 <= mul_loop_mul_if_land_1_lpi_1_dfm_9;
      mul_loop_mul_else_land_15_lpi_1_dfm_10 <= mul_loop_mul_else_land_15_lpi_1_dfm_9;
      mul_loop_mul_else_land_2_lpi_1_dfm_10 <= mul_loop_mul_else_land_2_lpi_1_dfm_9;
      mul_loop_mul_if_land_2_lpi_1_dfm_10 <= mul_loop_mul_if_land_2_lpi_1_dfm_9;
      mul_loop_mul_else_land_14_lpi_1_dfm_10 <= mul_loop_mul_else_land_14_lpi_1_dfm_9;
      mul_loop_mul_else_land_3_lpi_1_dfm_10 <= mul_loop_mul_else_land_3_lpi_1_dfm_9;
      mul_loop_mul_if_land_3_lpi_1_dfm_10 <= mul_loop_mul_if_land_3_lpi_1_dfm_9;
      mul_loop_mul_else_land_13_lpi_1_dfm_10 <= mul_loop_mul_else_land_13_lpi_1_dfm_9;
      mul_loop_mul_else_land_4_lpi_1_dfm_10 <= mul_loop_mul_else_land_4_lpi_1_dfm_9;
      mul_loop_mul_if_land_4_lpi_1_dfm_10 <= mul_loop_mul_if_land_4_lpi_1_dfm_9;
      mul_loop_mul_else_land_12_lpi_1_dfm_10 <= mul_loop_mul_else_land_12_lpi_1_dfm_9;
      mul_loop_mul_else_land_5_lpi_1_dfm_10 <= mul_loop_mul_else_land_5_lpi_1_dfm_9;
      mul_loop_mul_if_land_5_lpi_1_dfm_10 <= mul_loop_mul_if_land_5_lpi_1_dfm_9;
      mul_loop_mul_else_land_11_lpi_1_dfm_10 <= mul_loop_mul_else_land_11_lpi_1_dfm_9;
      mul_loop_mul_else_land_6_lpi_1_dfm_10 <= mul_loop_mul_else_land_6_lpi_1_dfm_9;
      mul_loop_mul_if_land_6_lpi_1_dfm_10 <= mul_loop_mul_if_land_6_lpi_1_dfm_9;
      mul_loop_mul_else_land_10_lpi_1_dfm_10 <= mul_loop_mul_else_land_10_lpi_1_dfm_9;
      mul_loop_mul_else_land_7_lpi_1_dfm_10 <= mul_loop_mul_else_land_7_lpi_1_dfm_9;
      mul_loop_mul_if_land_7_lpi_1_dfm_10 <= mul_loop_mul_if_land_7_lpi_1_dfm_9;
      mul_loop_mul_else_land_9_lpi_1_dfm_10 <= mul_loop_mul_else_land_9_lpi_1_dfm_9;
      mul_loop_mul_else_land_8_lpi_1_dfm_10 <= mul_loop_mul_else_land_8_lpi_1_dfm_9;
      mul_loop_mul_if_land_8_lpi_1_dfm_10 <= mul_loop_mul_if_land_8_lpi_1_dfm_9;
      mul_loop_mul_if_land_9_lpi_1_dfm_10 <= mul_loop_mul_if_land_9_lpi_1_dfm_9;
      mul_loop_mul_if_land_10_lpi_1_dfm_10 <= mul_loop_mul_if_land_10_lpi_1_dfm_9;
      mul_loop_mul_if_land_11_lpi_1_dfm_10 <= mul_loop_mul_if_land_11_lpi_1_dfm_9;
      mul_loop_mul_if_land_12_lpi_1_dfm_10 <= mul_loop_mul_if_land_12_lpi_1_dfm_9;
      mul_loop_mul_if_land_13_lpi_1_dfm_10 <= mul_loop_mul_if_land_13_lpi_1_dfm_9;
      mul_loop_mul_if_land_14_lpi_1_dfm_10 <= mul_loop_mul_if_land_14_lpi_1_dfm_9;
      mul_loop_mul_if_land_15_lpi_1_dfm_10 <= mul_loop_mul_if_land_15_lpi_1_dfm_9;
      mul_loop_mul_if_land_lpi_1_dfm_10 <= mul_loop_mul_if_land_lpi_1_dfm_9;
      io_read_cfg_mul_bypass_rsc_svs_st_7 <= io_read_cfg_mul_bypass_rsc_svs_st_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_12_itm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_408_nl)) ) begin
      FpMul_8U_23U_mux_12_itm_4 <= FpMul_8U_23U_mux_12_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_0_sva_10 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_412_nl)) ) begin
      MulOut_data_0_sva_10 <= MulOut_data_0_sva_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_28_itm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_415_nl)) ) begin
      FpMul_8U_23U_mux_28_itm_4 <= FpMul_8U_23U_mux_28_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_1_sva_10 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_418_nl)) ) begin
      MulOut_data_1_sva_10 <= MulOut_data_1_sva_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_44_itm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_421_nl)) ) begin
      FpMul_8U_23U_mux_44_itm_4 <= FpMul_8U_23U_mux_44_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_2_sva_10 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_424_nl)) ) begin
      MulOut_data_2_sva_10 <= MulOut_data_2_sva_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_60_itm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_427_nl)) ) begin
      FpMul_8U_23U_mux_60_itm_4 <= FpMul_8U_23U_mux_60_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_3_sva_10 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_430_nl)) ) begin
      MulOut_data_3_sva_10 <= MulOut_data_3_sva_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_76_itm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_433_nl)) ) begin
      FpMul_8U_23U_mux_76_itm_4 <= FpMul_8U_23U_mux_76_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_4_sva_10 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_436_nl)) ) begin
      MulOut_data_4_sva_10 <= MulOut_data_4_sva_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_92_itm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_439_nl)) ) begin
      FpMul_8U_23U_mux_92_itm_4 <= FpMul_8U_23U_mux_92_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_5_sva_10 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_442_nl)) ) begin
      MulOut_data_5_sva_10 <= MulOut_data_5_sva_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_108_itm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_445_nl)) ) begin
      FpMul_8U_23U_mux_108_itm_4 <= FpMul_8U_23U_mux_108_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_6_sva_10 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_448_nl)) ) begin
      MulOut_data_6_sva_10 <= MulOut_data_6_sva_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_124_itm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_451_nl)) ) begin
      FpMul_8U_23U_mux_124_itm_4 <= FpMul_8U_23U_mux_124_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_7_sva_10 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_454_nl)) ) begin
      MulOut_data_7_sva_10 <= MulOut_data_7_sva_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_140_itm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_457_nl)) ) begin
      FpMul_8U_23U_mux_140_itm_4 <= FpMul_8U_23U_mux_140_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_8_sva_10 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_460_nl)) ) begin
      MulOut_data_8_sva_10 <= MulOut_data_8_sva_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_156_itm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_463_nl)) ) begin
      FpMul_8U_23U_mux_156_itm_4 <= FpMul_8U_23U_mux_156_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_9_sva_10 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_466_nl)) ) begin
      MulOut_data_9_sva_10 <= MulOut_data_9_sva_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_172_itm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_469_nl)) ) begin
      FpMul_8U_23U_mux_172_itm_4 <= FpMul_8U_23U_mux_172_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_10_sva_10 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_472_nl)) ) begin
      MulOut_data_10_sva_10 <= MulOut_data_10_sva_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_188_itm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_475_nl)) ) begin
      FpMul_8U_23U_mux_188_itm_4 <= FpMul_8U_23U_mux_188_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_11_sva_10 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_478_nl)) ) begin
      MulOut_data_11_sva_10 <= MulOut_data_11_sva_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_204_itm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_481_nl)) ) begin
      FpMul_8U_23U_mux_204_itm_4 <= FpMul_8U_23U_mux_204_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_12_sva_10 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_484_nl)) ) begin
      MulOut_data_12_sva_10 <= MulOut_data_12_sva_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_220_itm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_487_nl)) ) begin
      FpMul_8U_23U_mux_220_itm_4 <= FpMul_8U_23U_mux_220_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_13_sva_10 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_490_nl)) ) begin
      MulOut_data_13_sva_10 <= MulOut_data_13_sva_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_236_itm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_493_nl)) ) begin
      FpMul_8U_23U_mux_236_itm_4 <= FpMul_8U_23U_mux_236_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_14_sva_10 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_496_nl)) ) begin
      MulOut_data_14_sva_10 <= MulOut_data_14_sva_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_252_itm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_499_nl)) ) begin
      FpMul_8U_23U_mux_252_itm_4 <= FpMul_8U_23U_mux_252_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_15_sva_10 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_502_nl)) ) begin
      MulOut_data_15_sva_10 <= MulOut_data_15_sva_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_1_itm <= 4'b0;
    end
    else if ( mux_1690_cse & core_wen & (~(mul_loop_mul_if_land_1_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
        | IsNaN_8U_23U_land_1_lpi_1_dfm_10)) & (~(mul_loop_mul_if_land_1_lpi_1_dfm_st_7
        | io_read_cfg_mul_bypass_rsc_svs_st_6)) & main_stage_v_3 & mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        & (~ FpMul_8U_23U_lor_18_lpi_1_dfm_st_3) & (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_8)
        & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_1_itm <= FpMul_8U_23U_p_expo_mux1h_1_itm[7:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_1_2_itm <= 4'b0;
    end
    else if ( (mux_1693_nl) & core_wen & (~ mul_loop_mul_if_land_1_lpi_1_dfm_9) &
        (~ io_read_cfg_mul_bypass_rsc_svs_7) & (~(IsNaN_8U_23U_land_1_lpi_1_dfm_10
        | mul_loop_mul_if_land_1_lpi_1_dfm_st_7)) & (~ io_read_cfg_mul_bypass_rsc_svs_st_6)
        & main_stage_v_3 & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_1_2_itm <= FpMul_8U_23U_p_expo_mux1h_1_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_512_nl)
        ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_mx0w0,
          FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_514_nl) ) begin
      mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_515_nl)) ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_9_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_9_1_0_1 <= 2'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_96_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_9_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_8_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_9_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_8_1_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_520_nl)
        ) begin
      mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_31_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_9_9_0_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_9_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_9_22_13_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_96_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_9_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_9_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_9_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_9_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_8_22_13_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_8 <= 1'b0;
      FpMul_8U_23U_lor_18_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_48_cse ) begin
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_8 <= IsNaN_8U_23U_land_1_lpi_1_dfm_st_7;
      FpMul_8U_23U_lor_18_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_18_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_18_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_523_itm) ) begin
      FpMul_8U_23U_lor_18_lpi_1_dfm_7 <= FpMul_8U_23U_lor_18_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_522_itm)
        ) begin
      mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs_st_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_31_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_1_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= 23'b0;
      FpMantRNE_48U_24U_else_carry_1_sva_2 <= 1'b0;
    end
    else if ( FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_cse ) begin
      mul_loop_mul_1_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= MUX_v_23_2_2((FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[45:23]), mul_loop_mul_1_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2,
          and_dcpl_104);
      FpMantRNE_48U_24U_else_carry_1_sva_2 <= MUX_s_1_2_2(FpMantRNE_48U_24U_else_carry_1_sva_mx0w0,
          FpMantRNE_48U_24U_else_carry_1_sva, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_523_itm)
        ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_itm_mx0w0,
          FpMul_8U_23U_FpMul_8U_23U_and_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_2_itm <= 4'b0;
    end
    else if ( mux_1695_cse & core_wen & (~(mul_loop_mul_if_land_2_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
        | IsNaN_8U_23U_land_2_lpi_1_dfm_10)) & (~(mul_loop_mul_if_land_2_lpi_1_dfm_st_7
        | io_read_cfg_mul_bypass_rsc_svs_st_6)) & main_stage_v_3 & mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        & (~ FpMul_8U_23U_lor_19_lpi_1_dfm_st_3) & (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_8)
        & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_2_itm <= FpMul_8U_23U_p_expo_mux1h_3_itm[7:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_2_2_itm <= 4'b0;
    end
    else if ( (mux_1698_nl) & core_wen & (~ mul_loop_mul_if_land_2_lpi_1_dfm_9) &
        (~ io_read_cfg_mul_bypass_rsc_svs_7) & (~(IsNaN_8U_23U_land_2_lpi_1_dfm_10
        | mul_loop_mul_if_land_2_lpi_1_dfm_st_7)) & (~ io_read_cfg_mul_bypass_rsc_svs_st_6)
        & main_stage_v_3 & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_2_2_itm <= FpMul_8U_23U_p_expo_mux1h_3_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_536_nl)
        ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_mx0w0,
          FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_538_nl)) ) begin
      mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_539_nl)) ) begin
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_9_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_9_1_0_1 <= 2'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_98_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_9_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_8_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_9_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_8_1_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_544_nl)
        ) begin
      mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_29_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_9_9_0_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_9_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_9_22_13_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_99_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_9_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_9_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_9_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_9_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_8_22_13_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_8 <= 1'b0;
      FpMul_8U_23U_lor_19_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_50_cse ) begin
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_8 <= IsNaN_8U_23U_land_2_lpi_1_dfm_st_7;
      FpMul_8U_23U_lor_19_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_19_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_19_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_547_itm) ) begin
      FpMul_8U_23U_lor_19_lpi_1_dfm_7 <= FpMul_8U_23U_lor_19_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_546_itm)
        ) begin
      mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs_st_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_29_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_2_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= 23'b0;
      FpMantRNE_48U_24U_else_carry_2_sva_2 <= 1'b0;
    end
    else if ( FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_1_cse ) begin
      mul_loop_mul_2_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= MUX_v_23_2_2((FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[45:23]), mul_loop_mul_2_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2,
          and_dcpl_104);
      FpMantRNE_48U_24U_else_carry_2_sva_2 <= MUX_s_1_2_2(FpMantRNE_48U_24U_else_carry_2_sva_mx0w0,
          FpMantRNE_48U_24U_else_carry_2_sva, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_64_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_547_itm)
        ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_64_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_64_itm_mx0w0,
          FpMul_8U_23U_FpMul_8U_23U_and_64_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_3_itm <= 4'b0;
    end
    else if ( mux_1700_cse & core_wen & (~(mul_loop_mul_if_land_3_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
        | IsNaN_8U_23U_land_3_lpi_1_dfm_10)) & (~(mul_loop_mul_if_land_3_lpi_1_dfm_st_7
        | io_read_cfg_mul_bypass_rsc_svs_st_6)) & main_stage_v_3 & mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        & (~ FpMul_8U_23U_lor_20_lpi_1_dfm_st_3) & (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_8)
        & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_3_itm <= FpMul_8U_23U_p_expo_mux1h_5_itm[7:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_3_2_itm <= 4'b0;
    end
    else if ( (mux_1703_nl) & core_wen & (~ mul_loop_mul_if_land_3_lpi_1_dfm_9) &
        (~ io_read_cfg_mul_bypass_rsc_svs_7) & (~(IsNaN_8U_23U_land_3_lpi_1_dfm_10
        | mul_loop_mul_if_land_3_lpi_1_dfm_st_7)) & (~ io_read_cfg_mul_bypass_rsc_svs_st_6)
        & main_stage_v_3 & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_3_2_itm <= FpMul_8U_23U_p_expo_mux1h_5_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_560_nl)
        ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_mx0w0,
          FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_562_nl) ) begin
      mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_563_nl)) ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_9_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_9_1_0_1 <= 2'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_100_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_9_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_8_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_9_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_8_1_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_568_nl)
        ) begin
      mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_27_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_9_9_0_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_9_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_9_22_13_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_102_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_9_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_9_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_9_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_9_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_8_22_13_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_8 <= 1'b0;
      FpMul_8U_23U_lor_20_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_52_cse ) begin
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_8 <= IsNaN_8U_23U_land_3_lpi_1_dfm_st_7;
      FpMul_8U_23U_lor_20_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_20_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_20_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_571_itm) ) begin
      FpMul_8U_23U_lor_20_lpi_1_dfm_7 <= FpMul_8U_23U_lor_20_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_570_itm)
        ) begin
      mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs_st_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_27_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_3_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= 23'b0;
      FpMantRNE_48U_24U_else_carry_3_sva_2 <= 1'b0;
    end
    else if ( FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_2_cse ) begin
      mul_loop_mul_3_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= MUX_v_23_2_2((FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[45:23]), mul_loop_mul_3_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2,
          and_dcpl_104);
      FpMantRNE_48U_24U_else_carry_3_sva_2 <= MUX_s_1_2_2(FpMantRNE_48U_24U_else_carry_3_sva_mx0w0,
          FpMantRNE_48U_24U_else_carry_3_sva, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_65_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_571_itm)
        ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_65_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_65_itm_mx0w0,
          FpMul_8U_23U_FpMul_8U_23U_and_65_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_4_itm <= 4'b0;
    end
    else if ( mux_1705_cse & core_wen & (~(mul_loop_mul_if_land_4_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
        | IsNaN_8U_23U_land_4_lpi_1_dfm_10)) & (~(mul_loop_mul_if_land_4_lpi_1_dfm_st_7
        | io_read_cfg_mul_bypass_rsc_svs_st_6)) & main_stage_v_3 & mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        & (~ FpMul_8U_23U_lor_21_lpi_1_dfm_st_3) & (~ IsNaN_8U_23U_1_land_4_lpi_1_dfm_8)
        & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_4_itm <= FpMul_8U_23U_p_expo_mux1h_7_itm[7:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_4_2_itm <= 4'b0;
    end
    else if ( (mux_1708_nl) & core_wen & (~ mul_loop_mul_if_land_4_lpi_1_dfm_9) &
        (~ io_read_cfg_mul_bypass_rsc_svs_7) & (~(IsNaN_8U_23U_land_4_lpi_1_dfm_10
        | mul_loop_mul_if_land_4_lpi_1_dfm_st_7)) & (~ io_read_cfg_mul_bypass_rsc_svs_st_6)
        & main_stage_v_3 & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_4_2_itm <= FpMul_8U_23U_p_expo_mux1h_7_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_584_nl)
        ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_mx0w0,
          FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_588_nl)) ) begin
      mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_4_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_589_nl)) ) begin
      IsNaN_8U_23U_1_land_4_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_4_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_9_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_9_1_0_1 <= 2'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_102_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_9_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_8_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_9_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_8_1_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_594_nl)
        ) begin
      mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_25_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_9_9_0_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_9_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_9_22_13_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_105_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_9_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_9_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_9_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_9_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_8_22_13_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_4_lpi_1_dfm_st_8 <= 1'b0;
      FpMul_8U_23U_lor_21_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_54_cse ) begin
      IsNaN_8U_23U_land_4_lpi_1_dfm_st_8 <= IsNaN_8U_23U_land_4_lpi_1_dfm_st_7;
      FpMul_8U_23U_lor_21_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_21_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_21_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_597_itm) ) begin
      FpMul_8U_23U_lor_21_lpi_1_dfm_7 <= FpMul_8U_23U_lor_21_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_596_itm)
        ) begin
      mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs_st_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_25_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_4_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= 23'b0;
      FpMantRNE_48U_24U_else_carry_4_sva_2 <= 1'b0;
    end
    else if ( FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_3_cse ) begin
      mul_loop_mul_4_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= MUX_v_23_2_2((FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[45:23]), mul_loop_mul_4_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2,
          and_dcpl_104);
      FpMantRNE_48U_24U_else_carry_4_sva_2 <= MUX_s_1_2_2(FpMantRNE_48U_24U_else_carry_4_sva_mx0w0,
          FpMantRNE_48U_24U_else_carry_4_sva, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_66_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_597_itm)
        ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_66_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_66_itm_mx0w0,
          FpMul_8U_23U_FpMul_8U_23U_and_66_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_5_itm <= 4'b0;
    end
    else if ( mux_1710_cse & core_wen & (~(mul_loop_mul_if_land_5_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
        | IsNaN_8U_23U_land_5_lpi_1_dfm_10)) & (~(mul_loop_mul_if_land_5_lpi_1_dfm_st_7
        | io_read_cfg_mul_bypass_rsc_svs_st_6)) & main_stage_v_3 & mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        & (~ FpMul_8U_23U_lor_22_lpi_1_dfm_st_3) & (~ IsNaN_8U_23U_1_land_5_lpi_1_dfm_8)
        & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_5_itm <= FpMul_8U_23U_p_expo_mux1h_9_itm[7:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_5_2_itm <= 4'b0;
    end
    else if ( (mux_1713_nl) & core_wen & (~ mul_loop_mul_if_land_5_lpi_1_dfm_9) &
        (~ io_read_cfg_mul_bypass_rsc_svs_7) & (~(IsNaN_8U_23U_land_5_lpi_1_dfm_10
        | mul_loop_mul_if_land_5_lpi_1_dfm_st_7)) & (~ io_read_cfg_mul_bypass_rsc_svs_st_6)
        & main_stage_v_3 & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_5_2_itm <= FpMul_8U_23U_p_expo_mux1h_9_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_4_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_610_nl)
        ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_4_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_4_itm_mx0w0,
          FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_4_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_612_nl)) ) begin
      mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_5_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_613_nl)) ) begin
      IsNaN_8U_23U_1_land_5_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_5_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_9_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_9_1_0_1 <= 2'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_104_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_9_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_8_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_9_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_8_1_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_618_nl)
        ) begin
      mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_23_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_9_9_0_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_9_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_9_22_13_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_108_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_9_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_9_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_9_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_9_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_8_22_13_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_5_lpi_1_dfm_st_8 <= 1'b0;
      FpMul_8U_23U_lor_22_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_56_cse ) begin
      IsNaN_8U_23U_land_5_lpi_1_dfm_st_8 <= IsNaN_8U_23U_land_5_lpi_1_dfm_st_7;
      FpMul_8U_23U_lor_22_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_22_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_22_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_621_itm) ) begin
      FpMul_8U_23U_lor_22_lpi_1_dfm_7 <= FpMul_8U_23U_lor_22_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_620_itm)
        ) begin
      mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs_st_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_23_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_5_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= 23'b0;
      FpMantRNE_48U_24U_else_carry_5_sva_2 <= 1'b0;
    end
    else if ( FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_4_cse ) begin
      mul_loop_mul_5_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= MUX_v_23_2_2((FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[45:23]), mul_loop_mul_5_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2,
          and_dcpl_104);
      FpMantRNE_48U_24U_else_carry_5_sva_2 <= MUX_s_1_2_2(FpMantRNE_48U_24U_else_carry_5_sva_mx0w0,
          FpMantRNE_48U_24U_else_carry_5_sva, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_67_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_621_itm)
        ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_67_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_67_itm_mx0w0,
          FpMul_8U_23U_FpMul_8U_23U_and_67_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_6_itm <= 4'b0;
    end
    else if ( mux_1715_cse & core_wen & (~(mul_loop_mul_if_land_6_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
        | IsNaN_8U_23U_land_6_lpi_1_dfm_10)) & (~(mul_loop_mul_if_land_6_lpi_1_dfm_st_7
        | io_read_cfg_mul_bypass_rsc_svs_st_6)) & main_stage_v_3 & mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        & (~ FpMul_8U_23U_lor_23_lpi_1_dfm_st_3) & (~ IsNaN_8U_23U_1_land_6_lpi_1_dfm_8)
        & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_6_itm <= FpMul_8U_23U_p_expo_mux1h_11_itm[7:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_6_2_itm <= 4'b0;
    end
    else if ( (mux_1718_nl) & core_wen & (~ mul_loop_mul_if_land_6_lpi_1_dfm_9) &
        (~ io_read_cfg_mul_bypass_rsc_svs_7) & (~(IsNaN_8U_23U_land_6_lpi_1_dfm_10
        | mul_loop_mul_if_land_6_lpi_1_dfm_st_7)) & (~ io_read_cfg_mul_bypass_rsc_svs_st_6)
        & main_stage_v_3 & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_6_2_itm <= FpMul_8U_23U_p_expo_mux1h_11_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_5_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_634_nl)
        ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_5_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_5_itm_mx0w0,
          FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_5_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_636_nl) ) begin
      mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_6_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_637_nl)) ) begin
      IsNaN_8U_23U_1_land_6_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_6_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_9_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_9_1_0_1 <= 2'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_106_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_9_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_8_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_9_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_8_1_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_642_nl)
        ) begin
      mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_21_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_9_9_0_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_9_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_9_22_13_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_111_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_9_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_9_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_9_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_9_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_8_22_13_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_6_lpi_1_dfm_st_8 <= 1'b0;
      FpMul_8U_23U_lor_23_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_58_cse ) begin
      IsNaN_8U_23U_land_6_lpi_1_dfm_st_8 <= IsNaN_8U_23U_land_6_lpi_1_dfm_st_7;
      FpMul_8U_23U_lor_23_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_23_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_23_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_645_itm) ) begin
      FpMul_8U_23U_lor_23_lpi_1_dfm_7 <= FpMul_8U_23U_lor_23_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_644_itm)
        ) begin
      mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs_st_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_21_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_6_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= 23'b0;
      FpMantRNE_48U_24U_else_carry_6_sva_2 <= 1'b0;
    end
    else if ( FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_5_cse ) begin
      mul_loop_mul_6_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= MUX_v_23_2_2((FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[45:23]), mul_loop_mul_6_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2,
          and_dcpl_104);
      FpMantRNE_48U_24U_else_carry_6_sva_2 <= MUX_s_1_2_2(FpMantRNE_48U_24U_else_carry_6_sva_mx0w0,
          FpMantRNE_48U_24U_else_carry_6_sva, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_68_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_645_itm)
        ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_68_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_68_itm_mx0w0,
          FpMul_8U_23U_FpMul_8U_23U_and_68_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_7_itm <= 4'b0;
    end
    else if ( mux_1720_cse & core_wen & (~(mul_loop_mul_if_land_7_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
        | IsNaN_8U_23U_land_7_lpi_1_dfm_10)) & (~(mul_loop_mul_if_land_7_lpi_1_dfm_st_7
        | io_read_cfg_mul_bypass_rsc_svs_st_6)) & main_stage_v_3 & mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        & (~ FpMul_8U_23U_lor_24_lpi_1_dfm_st_3) & (~ IsNaN_8U_23U_1_land_7_lpi_1_dfm_8)
        & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_7_itm <= FpMul_8U_23U_p_expo_mux1h_13_itm[7:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_7_2_itm <= 4'b0;
    end
    else if ( (mux_1723_nl) & core_wen & (~ mul_loop_mul_if_land_7_lpi_1_dfm_9) &
        (~ io_read_cfg_mul_bypass_rsc_svs_7) & (~(IsNaN_8U_23U_land_7_lpi_1_dfm_10
        | mul_loop_mul_if_land_7_lpi_1_dfm_st_7)) & (~ io_read_cfg_mul_bypass_rsc_svs_st_6)
        & main_stage_v_3 & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_7_2_itm <= FpMul_8U_23U_p_expo_mux1h_13_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_6_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_658_nl)
        ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_6_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_6_itm_mx0w0,
          FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_6_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_660_nl) ) begin
      mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_7_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_661_nl)) ) begin
      IsNaN_8U_23U_1_land_7_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_7_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_9_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_9_1_0_1 <= 2'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_108_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_9_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_8_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_9_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_8_1_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_666_nl)
        ) begin
      mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_19_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_9_9_0_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_9_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_9_22_13_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_114_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_9_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_9_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_9_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_9_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_8_22_13_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_7_lpi_1_dfm_st_8 <= 1'b0;
      FpMul_8U_23U_lor_24_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_60_cse ) begin
      IsNaN_8U_23U_land_7_lpi_1_dfm_st_8 <= IsNaN_8U_23U_land_7_lpi_1_dfm_st_7;
      FpMul_8U_23U_lor_24_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_24_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_24_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_669_itm) ) begin
      FpMul_8U_23U_lor_24_lpi_1_dfm_7 <= FpMul_8U_23U_lor_24_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_668_itm)
        ) begin
      mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs_st_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_19_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_7_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= 23'b0;
      FpMantRNE_48U_24U_else_carry_7_sva_2 <= 1'b0;
    end
    else if ( FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_6_cse ) begin
      mul_loop_mul_7_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= MUX_v_23_2_2((FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[45:23]), mul_loop_mul_7_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2,
          and_dcpl_104);
      FpMantRNE_48U_24U_else_carry_7_sva_2 <= MUX_s_1_2_2(FpMantRNE_48U_24U_else_carry_7_sva_mx0w0,
          FpMantRNE_48U_24U_else_carry_7_sva, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_69_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_669_itm)
        ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_69_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_69_itm_mx0w0,
          FpMul_8U_23U_FpMul_8U_23U_and_69_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_8_itm <= 4'b0;
    end
    else if ( mux_1725_cse & core_wen & (~(mul_loop_mul_if_land_8_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
        | IsNaN_8U_23U_land_8_lpi_1_dfm_10)) & (~(mul_loop_mul_if_land_8_lpi_1_dfm_st_7
        | io_read_cfg_mul_bypass_rsc_svs_st_6)) & main_stage_v_3 & mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        & (~ FpMul_8U_23U_lor_25_lpi_1_dfm_st_3) & (~ IsNaN_8U_23U_1_land_8_lpi_1_dfm_8)
        & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_8_itm <= FpMul_8U_23U_p_expo_mux1h_15_itm[7:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_8_2_itm <= 4'b0;
    end
    else if ( (mux_1728_nl) & core_wen & (~ mul_loop_mul_if_land_8_lpi_1_dfm_9) &
        (~ io_read_cfg_mul_bypass_rsc_svs_7) & (~(IsNaN_8U_23U_land_8_lpi_1_dfm_10
        | mul_loop_mul_if_land_8_lpi_1_dfm_st_7)) & (~ io_read_cfg_mul_bypass_rsc_svs_st_6)
        & main_stage_v_3 & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_8_2_itm <= FpMul_8U_23U_p_expo_mux1h_15_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_7_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_682_nl)
        ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_7_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_7_itm_mx0w0,
          FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_7_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_684_nl)) ) begin
      mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_8_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_685_nl)) ) begin
      IsNaN_8U_23U_1_land_8_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_8_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_9_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_9_1_0_1 <= 2'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_110_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_9_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_8_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_9_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_8_1_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_690_nl)
        ) begin
      mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_17_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_9_9_0_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_9_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_9_22_13_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_117_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_9_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_9_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_9_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_9_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_8_22_13_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_8_lpi_1_dfm_st_8 <= 1'b0;
      FpMul_8U_23U_lor_25_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_62_cse ) begin
      IsNaN_8U_23U_land_8_lpi_1_dfm_st_8 <= IsNaN_8U_23U_land_8_lpi_1_dfm_st_7;
      FpMul_8U_23U_lor_25_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_25_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_25_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_693_itm) ) begin
      FpMul_8U_23U_lor_25_lpi_1_dfm_7 <= FpMul_8U_23U_lor_25_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_692_itm)
        ) begin
      mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs_st_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_17_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_8_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= 23'b0;
      FpMantRNE_48U_24U_else_carry_8_sva_2 <= 1'b0;
    end
    else if ( FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_7_cse ) begin
      mul_loop_mul_8_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= MUX_v_23_2_2((FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[45:23]), mul_loop_mul_8_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2,
          and_dcpl_104);
      FpMantRNE_48U_24U_else_carry_8_sva_2 <= MUX_s_1_2_2(FpMantRNE_48U_24U_else_carry_8_sva_mx0w0,
          FpMantRNE_48U_24U_else_carry_8_sva, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_70_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_693_itm)
        ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_70_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_70_itm_mx0w0,
          FpMul_8U_23U_FpMul_8U_23U_and_70_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_9_itm <= 4'b0;
    end
    else if ( mux_1730_cse & core_wen & (~(mul_loop_mul_if_land_9_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
        | IsNaN_8U_23U_land_9_lpi_1_dfm_10)) & (~(mul_loop_mul_if_land_9_lpi_1_dfm_st_7
        | io_read_cfg_mul_bypass_rsc_svs_st_6)) & main_stage_v_3 & mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        & (~ FpMul_8U_23U_lor_26_lpi_1_dfm_st_3) & (~ IsNaN_8U_23U_1_land_9_lpi_1_dfm_8)
        & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_9_itm <= FpMul_8U_23U_p_expo_mux1h_17_itm[7:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_9_2_itm <= 4'b0;
    end
    else if ( (mux_1733_nl) & core_wen & (~ mul_loop_mul_if_land_9_lpi_1_dfm_9) &
        (~ io_read_cfg_mul_bypass_rsc_svs_7) & (~(IsNaN_8U_23U_land_9_lpi_1_dfm_10
        | mul_loop_mul_if_land_9_lpi_1_dfm_st_7)) & (~ io_read_cfg_mul_bypass_rsc_svs_st_6)
        & main_stage_v_3 & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_9_2_itm <= FpMul_8U_23U_p_expo_mux1h_17_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_8_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_706_nl)
        ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_8_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_8_itm_mx0w0,
          FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_8_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_708_nl)) ) begin
      mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_9_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_709_nl)) ) begin
      IsNaN_8U_23U_1_land_9_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_9_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_9_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_9_1_0_1 <= 2'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_112_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_9_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_8_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_9_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_8_1_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_714_nl)
        ) begin
      mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_15_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_9_9_0_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_9_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_9_22_13_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_120_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_9_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_9_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_9_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_9_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_8_22_13_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_9_lpi_1_dfm_st_8 <= 1'b0;
      FpMul_8U_23U_lor_26_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_64_cse ) begin
      IsNaN_8U_23U_land_9_lpi_1_dfm_st_8 <= IsNaN_8U_23U_land_9_lpi_1_dfm_st_7;
      FpMul_8U_23U_lor_26_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_26_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_26_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_717_itm) ) begin
      FpMul_8U_23U_lor_26_lpi_1_dfm_7 <= FpMul_8U_23U_lor_26_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_716_itm)
        ) begin
      mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs_st_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_15_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_9_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= 23'b0;
      FpMantRNE_48U_24U_else_carry_9_sva_2 <= 1'b0;
    end
    else if ( FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_8_cse ) begin
      mul_loop_mul_9_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= MUX_v_23_2_2((FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[45:23]), mul_loop_mul_9_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2,
          and_dcpl_104);
      FpMantRNE_48U_24U_else_carry_9_sva_2 <= MUX_s_1_2_2(FpMantRNE_48U_24U_else_carry_9_sva_mx0w0,
          FpMantRNE_48U_24U_else_carry_9_sva, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_71_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_717_itm)
        ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_71_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_71_itm_mx0w0,
          FpMul_8U_23U_FpMul_8U_23U_and_71_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_10_itm <= 4'b0;
    end
    else if ( mux_1735_cse & core_wen & (~(mul_loop_mul_if_land_10_lpi_1_dfm_9 |
        io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_land_10_lpi_1_dfm_10)) &
        (~(mul_loop_mul_if_land_10_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6))
        & main_stage_v_3 & mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        & (~ FpMul_8U_23U_lor_27_lpi_1_dfm_st_3) & (~ IsNaN_8U_23U_1_land_10_lpi_1_dfm_8)
        & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_10_itm <= FpMul_8U_23U_p_expo_mux1h_19_itm[7:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_10_2_itm <= 4'b0;
    end
    else if ( (mux_1738_nl) & core_wen & (~ mul_loop_mul_if_land_10_lpi_1_dfm_9)
        & (~ io_read_cfg_mul_bypass_rsc_svs_7) & (~(IsNaN_8U_23U_land_10_lpi_1_dfm_10
        | mul_loop_mul_if_land_10_lpi_1_dfm_st_7)) & (~ io_read_cfg_mul_bypass_rsc_svs_st_6)
        & main_stage_v_3 & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_10_2_itm <= FpMul_8U_23U_p_expo_mux1h_19_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_9_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_730_nl)
        ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_9_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_9_itm_mx0w0,
          FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_9_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_732_nl)) ) begin
      mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_10_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_733_nl)) ) begin
      IsNaN_8U_23U_1_land_10_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_10_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_9_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_9_1_0_1 <= 2'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_114_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_9_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_8_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_9_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_8_1_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_738_nl)
        ) begin
      mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_13_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_9_9_0_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_9_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_9_22_13_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_123_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_9_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_9_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_9_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_9_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_8_22_13_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_10_lpi_1_dfm_st_8 <= 1'b0;
      FpMul_8U_23U_lor_27_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_66_cse ) begin
      IsNaN_8U_23U_land_10_lpi_1_dfm_st_8 <= IsNaN_8U_23U_land_10_lpi_1_dfm_st_7;
      FpMul_8U_23U_lor_27_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_27_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_27_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_741_itm) ) begin
      FpMul_8U_23U_lor_27_lpi_1_dfm_7 <= FpMul_8U_23U_lor_27_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_740_itm)
        ) begin
      mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs_st_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_13_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_10_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= 23'b0;
      FpMantRNE_48U_24U_else_carry_10_sva_2 <= 1'b0;
    end
    else if ( FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_9_cse ) begin
      mul_loop_mul_10_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= MUX_v_23_2_2((FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[45:23]), mul_loop_mul_10_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2,
          and_dcpl_104);
      FpMantRNE_48U_24U_else_carry_10_sva_2 <= MUX_s_1_2_2(FpMantRNE_48U_24U_else_carry_10_sva_mx0w0,
          FpMantRNE_48U_24U_else_carry_10_sva, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_72_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_741_itm)
        ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_72_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_72_itm_mx0w0,
          FpMul_8U_23U_FpMul_8U_23U_and_72_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_11_itm <= 4'b0;
    end
    else if ( mux_1741_cse & core_wen & (~(io_read_cfg_mul_bypass_rsc_svs_7 | mul_loop_mul_if_land_11_lpi_1_dfm_9
        | IsNaN_8U_23U_land_11_lpi_1_dfm_10)) & main_stage_v_3 & (~ io_read_cfg_mul_bypass_rsc_svs_st_6)
        & (~ mul_loop_mul_if_land_11_lpi_1_dfm_st_7) & mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        & (~ FpMul_8U_23U_lor_28_lpi_1_dfm_st_3) & (~ IsNaN_8U_23U_1_land_11_lpi_1_dfm_8)
        & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_11_itm <= FpMul_8U_23U_p_expo_mux1h_21_itm[7:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_11_2_itm <= 4'b0;
    end
    else if ( (mux_1745_nl) & core_wen & (~ io_read_cfg_mul_bypass_rsc_svs_7) & (~
        mul_loop_mul_if_land_11_lpi_1_dfm_9) & (~ IsNaN_8U_23U_land_11_lpi_1_dfm_10)
        & main_stage_v_3 & (~(io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_11_lpi_1_dfm_st_7))
        & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_11_2_itm <= FpMul_8U_23U_p_expo_mux1h_21_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_10_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_754_nl)
        ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_10_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_10_itm_mx0w0,
          FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_10_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_759_nl)) ) begin
      mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_11_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_760_nl)) ) begin
      IsNaN_8U_23U_1_land_11_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_11_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_9_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_9_1_0_1 <= 2'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_116_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_9_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_8_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_9_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_8_1_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_765_nl)
        ) begin
      mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_11_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_9_9_0_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_9_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_9_22_13_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_126_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_9_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_9_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_9_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_9_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_8_22_13_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_11_lpi_1_dfm_st_8 <= 1'b0;
      FpMul_8U_23U_lor_28_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_68_cse ) begin
      IsNaN_8U_23U_land_11_lpi_1_dfm_st_8 <= IsNaN_8U_23U_land_11_lpi_1_dfm_st_7;
      FpMul_8U_23U_lor_28_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_28_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_28_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_767_itm) ) begin
      FpMul_8U_23U_lor_28_lpi_1_dfm_7 <= FpMul_8U_23U_lor_28_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_tmp_748)
        ) begin
      mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs_st_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_11_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_11_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= 23'b0;
      FpMantRNE_48U_24U_else_carry_11_sva_2 <= 1'b0;
    end
    else if ( FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_10_cse ) begin
      mul_loop_mul_11_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= MUX_v_23_2_2((FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[45:23]), mul_loop_mul_11_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2,
          and_dcpl_104);
      FpMantRNE_48U_24U_else_carry_11_sva_2 <= MUX_s_1_2_2(FpMantRNE_48U_24U_else_carry_11_sva_mx0w0,
          FpMantRNE_48U_24U_else_carry_11_sva, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_73_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_767_itm)
        ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_73_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_73_itm_mx0w0,
          FpMul_8U_23U_FpMul_8U_23U_and_73_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_12_itm <= 4'b0;
    end
    else if ( mux_1747_cse & core_wen & (~(mul_loop_mul_if_land_12_lpi_1_dfm_9 |
        io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_land_12_lpi_1_dfm_10)) &
        (~(mul_loop_mul_if_land_12_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6))
        & main_stage_v_3 & mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        & (~ FpMul_8U_23U_lor_29_lpi_1_dfm_st_3) & (~ IsNaN_8U_23U_1_land_12_lpi_1_dfm_8)
        & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_12_itm <= FpMul_8U_23U_p_expo_mux1h_23_itm[7:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_12_2_itm <= 4'b0;
    end
    else if ( (mux_1750_nl) & core_wen & (~ mul_loop_mul_if_land_12_lpi_1_dfm_9)
        & (~ io_read_cfg_mul_bypass_rsc_svs_7) & (~(IsNaN_8U_23U_land_12_lpi_1_dfm_10
        | mul_loop_mul_if_land_12_lpi_1_dfm_st_7)) & (~ io_read_cfg_mul_bypass_rsc_svs_st_6)
        & main_stage_v_3 & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_12_2_itm <= FpMul_8U_23U_p_expo_mux1h_23_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_11_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_781_nl)
        ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_11_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_11_itm_mx0w0,
          FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_11_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_785_nl)) ) begin
      mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_12_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_786_nl)) ) begin
      IsNaN_8U_23U_1_land_12_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_12_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_9_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_9_1_0_1 <= 2'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_118_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_9_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_8_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_9_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_8_1_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_791_nl)
        ) begin
      mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_9_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_9_9_0_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_9_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_9_22_13_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_129_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_9_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_9_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_9_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_9_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_8_22_13_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_12_lpi_1_dfm_st_8 <= 1'b0;
      FpMul_8U_23U_lor_29_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_70_cse ) begin
      IsNaN_8U_23U_land_12_lpi_1_dfm_st_8 <= IsNaN_8U_23U_land_12_lpi_1_dfm_st_7;
      FpMul_8U_23U_lor_29_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_29_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_29_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_794_itm) ) begin
      FpMul_8U_23U_lor_29_lpi_1_dfm_7 <= FpMul_8U_23U_lor_29_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_793_itm)
        ) begin
      mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs_st_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_9_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_12_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= 23'b0;
      FpMantRNE_48U_24U_else_carry_12_sva_2 <= 1'b0;
    end
    else if ( FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_11_cse ) begin
      mul_loop_mul_12_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= MUX_v_23_2_2((FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[45:23]), mul_loop_mul_12_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2,
          and_dcpl_104);
      FpMantRNE_48U_24U_else_carry_12_sva_2 <= MUX_s_1_2_2(FpMantRNE_48U_24U_else_carry_12_sva_mx0w0,
          FpMantRNE_48U_24U_else_carry_12_sva, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_74_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_794_itm)
        ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_74_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_74_itm_mx0w0,
          FpMul_8U_23U_FpMul_8U_23U_and_74_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_13_itm <= 4'b0;
    end
    else if ( mux_1752_cse & core_wen & (~(mul_loop_mul_if_land_13_lpi_1_dfm_9 |
        io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_land_13_lpi_1_dfm_10)) &
        (~(mul_loop_mul_if_land_13_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6))
        & main_stage_v_3 & mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        & (~ FpMul_8U_23U_lor_30_lpi_1_dfm_st_3) & (~ IsNaN_8U_23U_1_land_13_lpi_1_dfm_8)
        & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_13_itm <= FpMul_8U_23U_p_expo_mux1h_25_itm[7:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_13_2_itm <= 4'b0;
    end
    else if ( (mux_1755_nl) & core_wen & (~ mul_loop_mul_if_land_13_lpi_1_dfm_9)
        & (~ io_read_cfg_mul_bypass_rsc_svs_7) & (~(IsNaN_8U_23U_land_13_lpi_1_dfm_10
        | mul_loop_mul_if_land_13_lpi_1_dfm_st_7)) & (~ io_read_cfg_mul_bypass_rsc_svs_st_6)
        & main_stage_v_3 & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_13_2_itm <= FpMul_8U_23U_p_expo_mux1h_25_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_12_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_808_nl)
        ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_12_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_12_itm_mx0w0,
          FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_12_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_812_nl)) ) begin
      mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_13_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_813_nl)) ) begin
      IsNaN_8U_23U_1_land_13_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_13_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_9_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_9_1_0_1 <= 2'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_120_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_9_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_8_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_9_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_8_1_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_818_nl)
        ) begin
      mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_7_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_9_9_0_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_9_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_9_22_13_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_132_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_9_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_9_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_9_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_9_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_8_22_13_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_13_lpi_1_dfm_st_8 <= 1'b0;
      FpMul_8U_23U_lor_30_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_72_cse ) begin
      IsNaN_8U_23U_land_13_lpi_1_dfm_st_8 <= IsNaN_8U_23U_land_13_lpi_1_dfm_st_7;
      FpMul_8U_23U_lor_30_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_30_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_30_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_821_itm) ) begin
      FpMul_8U_23U_lor_30_lpi_1_dfm_7 <= FpMul_8U_23U_lor_30_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_820_itm)
        ) begin
      mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs_st_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_7_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_13_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= 23'b0;
      FpMantRNE_48U_24U_else_carry_13_sva_2 <= 1'b0;
    end
    else if ( FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_12_cse ) begin
      mul_loop_mul_13_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= MUX_v_23_2_2((FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[45:23]), mul_loop_mul_13_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2,
          and_dcpl_104);
      FpMantRNE_48U_24U_else_carry_13_sva_2 <= MUX_s_1_2_2(FpMantRNE_48U_24U_else_carry_13_sva_mx0w0,
          FpMantRNE_48U_24U_else_carry_13_sva, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_75_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_821_itm)
        ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_75_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_75_itm_mx0w0,
          FpMul_8U_23U_FpMul_8U_23U_and_75_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_14_itm <= 4'b0;
    end
    else if ( mux_1758_cse & core_wen & (~(io_read_cfg_mul_bypass_rsc_svs_st_6 |
        io_read_cfg_mul_bypass_rsc_svs_7 | mul_loop_mul_if_land_14_lpi_1_dfm_9))
        & (~(mul_loop_mul_if_land_14_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_14_lpi_1_dfm_10))
        & main_stage_v_3 & (~ FpMul_8U_23U_lor_31_lpi_1_dfm_st_3) & mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        & (~ IsNaN_8U_23U_1_land_14_lpi_1_dfm_8) & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_14_itm <= FpMul_8U_23U_p_expo_mux1h_27_itm[7:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_14_2_itm <= 4'b0;
    end
    else if ( (mux_1762_nl) & core_wen & (~ io_read_cfg_mul_bypass_rsc_svs_st_6)
        & (~ io_read_cfg_mul_bypass_rsc_svs_7) & (~(mul_loop_mul_if_land_14_lpi_1_dfm_9
        | mul_loop_mul_if_land_14_lpi_1_dfm_st_7)) & (~ IsNaN_8U_23U_land_14_lpi_1_dfm_10)
        & main_stage_v_3 & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_14_2_itm <= FpMul_8U_23U_p_expo_mux1h_27_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_13_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_835_nl)
        ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_13_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_13_itm_mx0w0,
          FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_13_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_837_nl) ) begin
      mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_14_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_838_nl)) ) begin
      IsNaN_8U_23U_1_land_14_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_14_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_9_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_9_1_0_1 <= 2'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_122_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_9_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_8_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_9_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_8_1_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_843_nl)
        ) begin
      mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_5_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_9_9_0_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_9_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_9_22_13_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_135_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_9_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_9_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_9_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_9_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_8_22_13_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_14_lpi_1_dfm_st_8 <= 1'b0;
      FpMul_8U_23U_lor_31_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_74_cse ) begin
      IsNaN_8U_23U_land_14_lpi_1_dfm_st_8 <= IsNaN_8U_23U_land_14_lpi_1_dfm_st_7;
      FpMul_8U_23U_lor_31_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_31_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_31_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_846_itm) ) begin
      FpMul_8U_23U_lor_31_lpi_1_dfm_7 <= FpMul_8U_23U_lor_31_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_845_itm)
        ) begin
      mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs_st_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_5_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_14_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= 23'b0;
      FpMantRNE_48U_24U_else_carry_14_sva_2 <= 1'b0;
    end
    else if ( FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_13_cse ) begin
      mul_loop_mul_14_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= MUX_v_23_2_2((FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[45:23]), mul_loop_mul_14_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2,
          and_dcpl_104);
      FpMantRNE_48U_24U_else_carry_14_sva_2 <= MUX_s_1_2_2(FpMantRNE_48U_24U_else_carry_14_sva_mx0w0,
          FpMantRNE_48U_24U_else_carry_14_sva, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_76_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_846_itm)
        ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_76_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_76_itm_mx0w0,
          FpMul_8U_23U_FpMul_8U_23U_and_76_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_15_itm <= 4'b0;
    end
    else if ( mux_1764_cse & core_wen & (~(mul_loop_mul_if_land_15_lpi_1_dfm_9 |
        io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_land_15_lpi_1_dfm_10)) &
        (~(mul_loop_mul_if_land_15_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6))
        & main_stage_v_3 & mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        & (~ FpMul_8U_23U_lor_32_lpi_1_dfm_st_3) & (~ IsNaN_8U_23U_1_land_15_lpi_1_dfm_8)
        & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_15_itm <= FpMul_8U_23U_p_expo_mux1h_29_itm[7:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_15_2_itm <= 4'b0;
    end
    else if ( (mux_1767_nl) & core_wen & (~ mul_loop_mul_if_land_15_lpi_1_dfm_9)
        & (~ io_read_cfg_mul_bypass_rsc_svs_7) & (~(IsNaN_8U_23U_land_15_lpi_1_dfm_10
        | mul_loop_mul_if_land_15_lpi_1_dfm_st_7)) & (~ io_read_cfg_mul_bypass_rsc_svs_st_6)
        & main_stage_v_3 & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_15_2_itm <= FpMul_8U_23U_p_expo_mux1h_29_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_14_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_860_nl)
        ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_14_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_14_itm_mx0w0,
          FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_14_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_862_nl) ) begin
      mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_15_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_863_nl)) ) begin
      IsNaN_8U_23U_1_land_15_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_15_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_9_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_9_1_0_1 <= 2'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_124_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_9_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_8_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_9_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_8_1_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_868_nl)
        ) begin
      mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_3_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_9_9_0_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_9_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_9_22_13_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_138_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_9_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_9_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_9_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_9_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_8_22_13_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_15_lpi_1_dfm_st_8 <= 1'b0;
      FpMul_8U_23U_lor_32_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_76_cse ) begin
      IsNaN_8U_23U_land_15_lpi_1_dfm_st_8 <= IsNaN_8U_23U_land_15_lpi_1_dfm_st_7;
      FpMul_8U_23U_lor_32_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_32_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_32_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_871_itm) ) begin
      FpMul_8U_23U_lor_32_lpi_1_dfm_7 <= FpMul_8U_23U_lor_32_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_870_itm)
        ) begin
      mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs_st_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_3_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_15_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= 23'b0;
      FpMantRNE_48U_24U_else_carry_15_sva_2 <= 1'b0;
    end
    else if ( FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_14_cse ) begin
      mul_loop_mul_15_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= MUX_v_23_2_2((FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[45:23]), mul_loop_mul_15_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2,
          and_dcpl_104);
      FpMantRNE_48U_24U_else_carry_15_sva_2 <= MUX_s_1_2_2(FpMantRNE_48U_24U_else_carry_15_sva_mx0w0,
          FpMantRNE_48U_24U_else_carry_15_sva, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_77_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_871_itm)
        ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_77_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_77_itm_mx0w0,
          FpMul_8U_23U_FpMul_8U_23U_and_77_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_itm <= 4'b0;
    end
    else if ( mux_1769_cse & core_wen & (~(mul_loop_mul_if_land_lpi_1_dfm_9 | io_read_cfg_mul_bypass_rsc_svs_7
        | IsNaN_8U_23U_land_lpi_1_dfm_10)) & (~(mul_loop_mul_if_land_lpi_1_dfm_st_7
        | io_read_cfg_mul_bypass_rsc_svs_st_6)) & main_stage_v_3 & mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        & (~ FpMul_8U_23U_lor_1_lpi_1_dfm_st_3) & (~ IsNaN_8U_23U_1_land_lpi_1_dfm_8)
        & or_309_cse ) begin
      reg_FpMul_8U_23U_p_expo_itm <= FpMul_8U_23U_p_expo_mux1h_31_itm[7:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_8U_23U_p_expo_2_itm_1 <= 4'b0;
    end
    else if ( (mux_1772_nl) & core_wen & (~ mul_loop_mul_if_land_lpi_1_dfm_9) & (~
        io_read_cfg_mul_bypass_rsc_svs_7) & (~(IsNaN_8U_23U_land_lpi_1_dfm_10 | mul_loop_mul_if_land_lpi_1_dfm_st_7))
        & (~ io_read_cfg_mul_bypass_rsc_svs_st_6) & main_stage_v_3 & or_309_cse )
        begin
      reg_FpMul_8U_23U_p_expo_2_itm_1 <= FpMul_8U_23U_p_expo_mux1h_31_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_15_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_885_nl)
        ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_15_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_15_itm_mx0w0,
          FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_15_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_887_nl)) ) begin
      mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_888_nl)) ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_9_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_9_1_0_1 <= 2'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_126_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_9_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_8_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_9_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_8_1_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (mux_893_nl)
        ) begin
      mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_1_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_9_9_0_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_9_12_10_1 <= 3'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_9_22_13_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_141_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_9_9_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_9_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_9_12_10_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_12_10_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_9_22_13_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_8_22_13_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_st_8 <= 1'b0;
      FpMul_8U_23U_lor_1_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_78_cse ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_st_8 <= IsNaN_8U_23U_land_lpi_1_dfm_st_7;
      FpMul_8U_23U_lor_1_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_1_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_896_itm) ) begin
      FpMul_8U_23U_lor_1_lpi_1_dfm_7 <= FpMul_8U_23U_lor_1_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_895_itm)
        ) begin
      mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs_st_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_1_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_16_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= 23'b0;
      FpMantRNE_48U_24U_else_carry_sva_2 <= 1'b0;
    end
    else if ( FpMantWidthDec_8U_47U_23U_0U_0U_overflow_and_15_cse ) begin
      mul_loop_mul_16_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_3
          <= MUX_v_23_2_2((FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[45:23]), mul_loop_mul_16_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2,
          and_dcpl_104);
      FpMantRNE_48U_24U_else_carry_sva_2 <= MUX_s_1_2_2(FpMantRNE_48U_24U_else_carry_sva_mx0w0,
          FpMantRNE_48U_24U_else_carry_sva, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_78_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ mux_896_itm)
        ) begin
      FpMul_8U_23U_FpMul_8U_23U_and_78_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_78_itm_mx0w0,
          FpMul_8U_23U_FpMul_8U_23U_and_78_itm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_if_land_lpi_1_dfm_st_8 <= 1'b0;
      mul_loop_mul_if_land_15_lpi_1_dfm_st_8 <= 1'b0;
      mul_loop_mul_if_land_14_lpi_1_dfm_st_8 <= 1'b0;
      mul_loop_mul_if_land_13_lpi_1_dfm_st_8 <= 1'b0;
      mul_loop_mul_if_land_12_lpi_1_dfm_st_8 <= 1'b0;
      mul_loop_mul_if_land_11_lpi_1_dfm_st_8 <= 1'b0;
      mul_loop_mul_if_land_10_lpi_1_dfm_st_8 <= 1'b0;
      mul_loop_mul_if_land_9_lpi_1_dfm_st_8 <= 1'b0;
      mul_loop_mul_if_land_8_lpi_1_dfm_st_8 <= 1'b0;
      mul_loop_mul_if_land_7_lpi_1_dfm_st_8 <= 1'b0;
      mul_loop_mul_if_land_6_lpi_1_dfm_st_8 <= 1'b0;
      mul_loop_mul_if_land_5_lpi_1_dfm_st_8 <= 1'b0;
      mul_loop_mul_if_land_4_lpi_1_dfm_st_8 <= 1'b0;
      mul_loop_mul_if_land_3_lpi_1_dfm_st_8 <= 1'b0;
      mul_loop_mul_if_land_2_lpi_1_dfm_st_8 <= 1'b0;
      mul_loop_mul_if_land_1_lpi_1_dfm_st_8 <= 1'b0;
    end
    else if ( mul_loop_mul_if_aelse_and_64_cse ) begin
      mul_loop_mul_if_land_lpi_1_dfm_st_8 <= mul_loop_mul_if_land_lpi_1_dfm_st_7;
      mul_loop_mul_if_land_15_lpi_1_dfm_st_8 <= mul_loop_mul_if_land_15_lpi_1_dfm_st_7;
      mul_loop_mul_if_land_14_lpi_1_dfm_st_8 <= mul_loop_mul_if_land_14_lpi_1_dfm_st_7;
      mul_loop_mul_if_land_13_lpi_1_dfm_st_8 <= mul_loop_mul_if_land_13_lpi_1_dfm_st_7;
      mul_loop_mul_if_land_12_lpi_1_dfm_st_8 <= mul_loop_mul_if_land_12_lpi_1_dfm_st_7;
      mul_loop_mul_if_land_11_lpi_1_dfm_st_8 <= mul_loop_mul_if_land_11_lpi_1_dfm_st_7;
      mul_loop_mul_if_land_10_lpi_1_dfm_st_8 <= mul_loop_mul_if_land_10_lpi_1_dfm_st_7;
      mul_loop_mul_if_land_9_lpi_1_dfm_st_8 <= mul_loop_mul_if_land_9_lpi_1_dfm_st_7;
      mul_loop_mul_if_land_8_lpi_1_dfm_st_8 <= mul_loop_mul_if_land_8_lpi_1_dfm_st_7;
      mul_loop_mul_if_land_7_lpi_1_dfm_st_8 <= mul_loop_mul_if_land_7_lpi_1_dfm_st_7;
      mul_loop_mul_if_land_6_lpi_1_dfm_st_8 <= mul_loop_mul_if_land_6_lpi_1_dfm_st_7;
      mul_loop_mul_if_land_5_lpi_1_dfm_st_8 <= mul_loop_mul_if_land_5_lpi_1_dfm_st_7;
      mul_loop_mul_if_land_4_lpi_1_dfm_st_8 <= mul_loop_mul_if_land_4_lpi_1_dfm_st_7;
      mul_loop_mul_if_land_3_lpi_1_dfm_st_8 <= mul_loop_mul_if_land_3_lpi_1_dfm_st_7;
      mul_loop_mul_if_land_2_lpi_1_dfm_st_8 <= mul_loop_mul_if_land_2_lpi_1_dfm_st_7;
      mul_loop_mul_if_land_1_lpi_1_dfm_st_8 <= mul_loop_mul_if_land_1_lpi_1_dfm_st_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_92) & (mux_902_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_2
          <= mul_loop_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs <= 1'b0;
      FpMantRNE_48U_24U_else_carry_1_sva <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_itm <= 1'b0;
    end
    else if ( FpMantRNE_48U_24U_else_and_cse ) begin
      mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs <= mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs_mx0w0;
      FpMantRNE_48U_24U_else_carry_1_sva <= FpMantRNE_48U_24U_else_carry_1_sva_mx0w0;
      FpMul_8U_23U_FpMul_8U_23U_and_itm <= FpMul_8U_23U_FpMul_8U_23U_and_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_1_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= 23'b0;
    end
    else if ( core_wen & (~ or_dcpl_96) & (mux_905_nl) ) begin
      mul_loop_mul_1_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[45:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_1_sva_1 <= 8'b0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm <= 1'b0;
      mul_loop_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <=
          1'b0;
    end
    else if ( FpMul_8U_23U_p_expo_and_cse ) begin
      FpMul_8U_23U_p_expo_1_sva_1 <= FpMul_8U_23U_p_expo_1_sva_1_mx0w0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm <= FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_mx0w0;
      mul_loop_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <=
          mul_loop_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_100) & (mux_907_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_2
          <= mul_loop_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs <= 1'b0;
      FpMantRNE_48U_24U_else_carry_2_sva <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_64_itm <= 1'b0;
    end
    else if ( FpMantRNE_48U_24U_else_and_2_cse ) begin
      mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs <= mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs_mx0w0;
      FpMantRNE_48U_24U_else_carry_2_sva <= FpMantRNE_48U_24U_else_carry_2_sva_mx0w0;
      FpMul_8U_23U_FpMul_8U_23U_and_64_itm <= FpMul_8U_23U_FpMul_8U_23U_and_64_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_2_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= 23'b0;
    end
    else if ( core_wen & (~ or_dcpl_103) & (mux_910_nl) ) begin
      mul_loop_mul_2_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[45:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_2_sva_1 <= 8'b0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm <= 1'b0;
      mul_loop_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <=
          1'b0;
    end
    else if ( FpMul_8U_23U_p_expo_and_1_cse ) begin
      FpMul_8U_23U_p_expo_2_sva_1 <= FpMul_8U_23U_p_expo_2_sva_1_mx0w0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm <= FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_mx0w0;
      mul_loop_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <=
          mul_loop_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_107) & (mux_912_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_2
          <= mul_loop_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_3_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= 23'b0;
    end
    else if ( core_wen & (~ or_dcpl_110) & (mux_915_nl) ) begin
      mul_loop_mul_3_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[45:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_48U_24U_else_carry_3_sva <= 1'b0;
      mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_65_itm <= 1'b0;
    end
    else if ( FpMantRNE_48U_24U_else_carry_and_2_cse ) begin
      FpMantRNE_48U_24U_else_carry_3_sva <= FpMantRNE_48U_24U_else_carry_3_sva_mx0w0;
      mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs <= mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs_mx0w0;
      FpMul_8U_23U_FpMul_8U_23U_and_65_itm <= FpMul_8U_23U_FpMul_8U_23U_and_65_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_3_sva_1 <= 8'b0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm <= 1'b0;
      mul_loop_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <=
          1'b0;
    end
    else if ( FpMul_8U_23U_p_expo_and_2_cse ) begin
      FpMul_8U_23U_p_expo_3_sva_1 <= FpMul_8U_23U_p_expo_3_sva_1_mx0w0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm <= FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_mx0w0;
      mul_loop_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <=
          mul_loop_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_4_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_115) & (mux_917_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_4_sva_st_2
          <= mul_loop_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs <= 1'b0;
      FpMantRNE_48U_24U_else_carry_4_sva <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_66_itm <= 1'b0;
    end
    else if ( FpMantRNE_48U_24U_else_and_6_cse ) begin
      mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs <= mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs_mx0w0;
      FpMantRNE_48U_24U_else_carry_4_sva <= FpMantRNE_48U_24U_else_carry_4_sva_mx0w0;
      FpMul_8U_23U_FpMul_8U_23U_and_66_itm <= FpMul_8U_23U_FpMul_8U_23U_and_66_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_4_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= 23'b0;
    end
    else if ( core_wen & (~ or_dcpl_118) & (mux_920_nl) ) begin
      mul_loop_mul_4_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= FpMul_8U_23U_p_mant_46_1_4_lpi_1_dfm_3_mx0[45:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_4_sva_1 <= 8'b0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm <= 1'b0;
      mul_loop_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <=
          1'b0;
    end
    else if ( FpMul_8U_23U_p_expo_and_3_cse ) begin
      FpMul_8U_23U_p_expo_4_sva_1 <= FpMul_8U_23U_p_expo_4_sva_1_mx0w0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm <= FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_mx0w0;
      mul_loop_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <=
          mul_loop_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_5_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_122) & (mux_922_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_5_sva_st_2
          <= mul_loop_mul_5_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs <= 1'b0;
      FpMantRNE_48U_24U_else_carry_5_sva <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_67_itm <= 1'b0;
    end
    else if ( FpMantRNE_48U_24U_else_and_8_cse ) begin
      mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs <= mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs_mx0w0;
      FpMantRNE_48U_24U_else_carry_5_sva <= FpMantRNE_48U_24U_else_carry_5_sva_mx0w0;
      FpMul_8U_23U_FpMul_8U_23U_and_67_itm <= FpMul_8U_23U_FpMul_8U_23U_and_67_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_5_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= 23'b0;
    end
    else if ( core_wen & (~ or_dcpl_125) & (mux_925_nl) ) begin
      mul_loop_mul_5_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= FpMul_8U_23U_p_mant_46_1_5_lpi_1_dfm_3_mx0[45:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_5_sva_1 <= 8'b0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_4_itm <= 1'b0;
      mul_loop_mul_5_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <=
          1'b0;
    end
    else if ( FpMul_8U_23U_p_expo_and_4_cse ) begin
      FpMul_8U_23U_p_expo_5_sva_1 <= FpMul_8U_23U_p_expo_5_sva_1_mx0w0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_4_itm <= FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_4_itm_mx0w0;
      mul_loop_mul_5_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <=
          mul_loop_mul_5_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_6_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_129) & (mux_927_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_6_sva_st_2
          <= mul_loop_mul_6_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs <= 1'b0;
      FpMantRNE_48U_24U_else_carry_6_sva <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_68_itm <= 1'b0;
    end
    else if ( FpMantRNE_48U_24U_else_and_10_cse ) begin
      mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs <= mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs_mx0w0;
      FpMantRNE_48U_24U_else_carry_6_sva <= FpMantRNE_48U_24U_else_carry_6_sva_mx0w0;
      FpMul_8U_23U_FpMul_8U_23U_and_68_itm <= FpMul_8U_23U_FpMul_8U_23U_and_68_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_6_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= 23'b0;
    end
    else if ( core_wen & (~ or_dcpl_132) & (mux_932_nl) ) begin
      mul_loop_mul_6_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= FpMul_8U_23U_p_mant_46_1_6_lpi_1_dfm_3_mx0[45:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_6_sva_1 <= 8'b0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_5_itm <= 1'b0;
      mul_loop_mul_6_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <=
          1'b0;
    end
    else if ( FpMul_8U_23U_p_expo_and_5_cse ) begin
      FpMul_8U_23U_p_expo_6_sva_1 <= FpMul_8U_23U_p_expo_6_sva_1_mx0w0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_5_itm <= FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_5_itm_mx0w0;
      mul_loop_mul_6_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <=
          mul_loop_mul_6_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_7_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_136) & (mux_934_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_7_sva_st_2
          <= mul_loop_mul_7_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_7_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= 23'b0;
    end
    else if ( core_wen & (~ or_dcpl_139) & (mux_937_nl) ) begin
      mul_loop_mul_7_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= FpMul_8U_23U_p_mant_46_1_7_lpi_1_dfm_3_mx0[45:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_48U_24U_else_carry_7_sva <= 1'b0;
      mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_69_itm <= 1'b0;
    end
    else if ( FpMantRNE_48U_24U_else_carry_and_6_cse ) begin
      FpMantRNE_48U_24U_else_carry_7_sva <= FpMantRNE_48U_24U_else_carry_7_sva_mx0w0;
      mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs <= mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs_mx0w0;
      FpMul_8U_23U_FpMul_8U_23U_and_69_itm <= FpMul_8U_23U_FpMul_8U_23U_and_69_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_7_sva_1 <= 8'b0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_6_itm <= 1'b0;
      mul_loop_mul_7_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <=
          1'b0;
    end
    else if ( FpMul_8U_23U_p_expo_and_6_cse ) begin
      FpMul_8U_23U_p_expo_7_sva_1 <= FpMul_8U_23U_p_expo_7_sva_1_mx0w0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_6_itm <= FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_6_itm_mx0w0;
      mul_loop_mul_7_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <=
          mul_loop_mul_7_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_8_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_143) & (mux_939_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_8_sva_st_2
          <= mul_loop_mul_8_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs <= 1'b0;
      FpMantRNE_48U_24U_else_carry_8_sva <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_70_itm <= 1'b0;
    end
    else if ( FpMantRNE_48U_24U_else_and_14_cse ) begin
      mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs <= mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs_mx0w0;
      FpMantRNE_48U_24U_else_carry_8_sva <= FpMantRNE_48U_24U_else_carry_8_sva_mx0w0;
      FpMul_8U_23U_FpMul_8U_23U_and_70_itm <= FpMul_8U_23U_FpMul_8U_23U_and_70_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_8_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= 23'b0;
    end
    else if ( core_wen & (~ or_dcpl_146) & (mux_942_nl) ) begin
      mul_loop_mul_8_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= FpMul_8U_23U_p_mant_46_1_8_lpi_1_dfm_3_mx0[45:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_8_sva_1 <= 8'b0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_7_itm <= 1'b0;
      mul_loop_mul_8_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <=
          1'b0;
    end
    else if ( FpMul_8U_23U_p_expo_and_7_cse ) begin
      FpMul_8U_23U_p_expo_8_sva_1 <= FpMul_8U_23U_p_expo_8_sva_1_mx0w0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_7_itm <= FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_7_itm_mx0w0;
      mul_loop_mul_8_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <=
          mul_loop_mul_8_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_9_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_150) & (mux_944_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_9_sva_st_2
          <= mul_loop_mul_9_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs <= 1'b0;
      FpMantRNE_48U_24U_else_carry_9_sva <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_71_itm <= 1'b0;
    end
    else if ( FpMantRNE_48U_24U_else_and_16_cse ) begin
      mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs <= mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs_mx0w0;
      FpMantRNE_48U_24U_else_carry_9_sva <= FpMantRNE_48U_24U_else_carry_9_sva_mx0w0;
      FpMul_8U_23U_FpMul_8U_23U_and_71_itm <= FpMul_8U_23U_FpMul_8U_23U_and_71_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_9_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= 23'b0;
    end
    else if ( core_wen & (~ or_dcpl_153) & (mux_947_nl) ) begin
      mul_loop_mul_9_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= FpMul_8U_23U_p_mant_46_1_9_lpi_1_dfm_3_mx0[45:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_9_sva_1 <= 8'b0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_8_itm <= 1'b0;
      mul_loop_mul_9_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <=
          1'b0;
    end
    else if ( FpMul_8U_23U_p_expo_and_8_cse ) begin
      FpMul_8U_23U_p_expo_9_sva_1 <= FpMul_8U_23U_p_expo_9_sva_1_mx0w0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_8_itm <= FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_8_itm_mx0w0;
      mul_loop_mul_9_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <=
          mul_loop_mul_9_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_10_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_157) & (mux_949_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_10_sva_st_2
          <= mul_loop_mul_10_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs <= 1'b0;
      FpMantRNE_48U_24U_else_carry_10_sva <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_72_itm <= 1'b0;
    end
    else if ( FpMantRNE_48U_24U_else_and_18_cse ) begin
      mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs <= mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs_mx0w0;
      FpMantRNE_48U_24U_else_carry_10_sva <= FpMantRNE_48U_24U_else_carry_10_sva_mx0w0;
      FpMul_8U_23U_FpMul_8U_23U_and_72_itm <= FpMul_8U_23U_FpMul_8U_23U_and_72_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_10_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= 23'b0;
    end
    else if ( core_wen & (~ or_dcpl_160) & (mux_954_nl) ) begin
      mul_loop_mul_10_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= FpMul_8U_23U_p_mant_46_1_10_lpi_1_dfm_3_mx0[45:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_10_sva_1 <= 8'b0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_9_itm <= 1'b0;
      mul_loop_mul_10_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_p_expo_and_9_cse ) begin
      FpMul_8U_23U_p_expo_10_sva_1 <= FpMul_8U_23U_p_expo_10_sva_1_mx0w0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_9_itm <= FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_9_itm_mx0w0;
      mul_loop_mul_10_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
          <= mul_loop_mul_10_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_11_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_165) & (mux_956_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_11_sva_st_2
          <= mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs <= 1'b0;
      FpMantRNE_48U_24U_else_carry_11_sva <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_73_itm <= 1'b0;
    end
    else if ( FpMantRNE_48U_24U_else_and_20_cse ) begin
      mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs <= mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs_mx0w0;
      FpMantRNE_48U_24U_else_carry_11_sva <= FpMantRNE_48U_24U_else_carry_11_sva_mx0w0;
      FpMul_8U_23U_FpMul_8U_23U_and_73_itm <= FpMul_8U_23U_FpMul_8U_23U_and_73_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_11_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= 23'b0;
    end
    else if ( core_wen & (~ or_dcpl_168) & (mux_959_nl) ) begin
      mul_loop_mul_11_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= FpMul_8U_23U_p_mant_46_1_11_lpi_1_dfm_3_mx0[45:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_11_sva_1 <= 8'b0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_10_itm <= 1'b0;
      mul_loop_mul_11_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_p_expo_and_10_cse ) begin
      FpMul_8U_23U_p_expo_11_sva_1 <= FpMul_8U_23U_p_expo_11_sva_1_mx0w0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_10_itm <= FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_10_itm_mx0w0;
      mul_loop_mul_11_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
          <= mul_loop_mul_11_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_12_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_173) & (mux_961_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_12_sva_st_2
          <= mul_loop_mul_12_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs <= 1'b0;
      FpMantRNE_48U_24U_else_carry_12_sva <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_74_itm <= 1'b0;
    end
    else if ( FpMantRNE_48U_24U_else_and_22_cse ) begin
      mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs <= mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs_mx0w0;
      FpMantRNE_48U_24U_else_carry_12_sva <= FpMantRNE_48U_24U_else_carry_12_sva_mx0w0;
      FpMul_8U_23U_FpMul_8U_23U_and_74_itm <= FpMul_8U_23U_FpMul_8U_23U_and_74_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_12_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= 23'b0;
    end
    else if ( core_wen & (~ or_dcpl_176) & (mux_964_nl) ) begin
      mul_loop_mul_12_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= FpMul_8U_23U_p_mant_46_1_12_lpi_1_dfm_3_mx0[45:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_12_sva_1 <= 8'b0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_11_itm <= 1'b0;
      mul_loop_mul_12_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_p_expo_and_11_cse ) begin
      FpMul_8U_23U_p_expo_12_sva_1 <= FpMul_8U_23U_p_expo_12_sva_1_mx0w0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_11_itm <= FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_11_itm_mx0w0;
      mul_loop_mul_12_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
          <= mul_loop_mul_12_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_13_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_181) & (mux_966_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_13_sva_st_2
          <= mul_loop_mul_13_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_13_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= 23'b0;
    end
    else if ( core_wen & (~ or_dcpl_184) & (mux_969_nl) ) begin
      mul_loop_mul_13_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= FpMul_8U_23U_p_mant_46_1_13_lpi_1_dfm_3_mx0[45:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs <= 1'b0;
      FpMantRNE_48U_24U_else_carry_13_sva <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_75_itm <= 1'b0;
    end
    else if ( FpMantRNE_48U_24U_else_and_24_cse ) begin
      mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs <= mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs_mx0w0;
      FpMantRNE_48U_24U_else_carry_13_sva <= FpMantRNE_48U_24U_else_carry_13_sva_mx0w0;
      FpMul_8U_23U_FpMul_8U_23U_and_75_itm <= FpMul_8U_23U_FpMul_8U_23U_and_75_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_13_sva_1 <= 8'b0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_12_itm <= 1'b0;
      mul_loop_mul_13_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_p_expo_and_12_cse ) begin
      FpMul_8U_23U_p_expo_13_sva_1 <= FpMul_8U_23U_p_expo_13_sva_1_mx0w0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_12_itm <= FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_12_itm_mx0w0;
      mul_loop_mul_13_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
          <= mul_loop_mul_13_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_14_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_188) & (mux_971_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_14_sva_st_2
          <= mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs <= 1'b0;
      FpMantRNE_48U_24U_else_carry_14_sva <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_76_itm <= 1'b0;
    end
    else if ( FpMantRNE_48U_24U_else_and_26_cse ) begin
      mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs <= mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs_mx0w0;
      FpMantRNE_48U_24U_else_carry_14_sva <= FpMantRNE_48U_24U_else_carry_14_sva_mx0w0;
      FpMul_8U_23U_FpMul_8U_23U_and_76_itm <= FpMul_8U_23U_FpMul_8U_23U_and_76_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_14_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= 23'b0;
    end
    else if ( core_wen & (~ or_dcpl_191) & (mux_974_nl) ) begin
      mul_loop_mul_14_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= FpMul_8U_23U_p_mant_46_1_14_lpi_1_dfm_3_mx0[45:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_14_sva_1 <= 8'b0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_13_itm <= 1'b0;
      mul_loop_mul_14_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_p_expo_and_13_cse ) begin
      FpMul_8U_23U_p_expo_14_sva_1 <= FpMul_8U_23U_p_expo_14_sva_1_mx0w0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_13_itm <= FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_13_itm_mx0w0;
      mul_loop_mul_14_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
          <= mul_loop_mul_14_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_15_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_195) & (mux_976_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_15_sva_st_2
          <= mul_loop_mul_15_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs <= 1'b0;
      FpMantRNE_48U_24U_else_carry_15_sva <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_77_itm <= 1'b0;
    end
    else if ( FpMantRNE_48U_24U_else_and_28_cse ) begin
      mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs <= mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs_mx0w0;
      FpMantRNE_48U_24U_else_carry_15_sva <= FpMantRNE_48U_24U_else_carry_15_sva_mx0w0;
      FpMul_8U_23U_FpMul_8U_23U_and_77_itm <= FpMul_8U_23U_FpMul_8U_23U_and_77_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_15_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= 23'b0;
    end
    else if ( core_wen & (~ or_dcpl_198) & (mux_979_nl) ) begin
      mul_loop_mul_15_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= FpMul_8U_23U_p_mant_46_1_15_lpi_1_dfm_3_mx0[45:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_15_sva_1 <= 8'b0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_14_itm <= 1'b0;
      mul_loop_mul_15_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_p_expo_and_14_cse ) begin
      FpMul_8U_23U_p_expo_15_sva_1 <= FpMul_8U_23U_p_expo_15_sva_1_mx0w0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_14_itm <= FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_14_itm_mx0w0;
      mul_loop_mul_15_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
          <= mul_loop_mul_15_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_202) & (mux_982_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_2
          <= mul_loop_mul_16_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_48U_24U_else_carry_sva <= 1'b0;
      mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_78_itm <= 1'b0;
    end
    else if ( FpMantRNE_48U_24U_else_carry_and_15_cse ) begin
      FpMantRNE_48U_24U_else_carry_sva <= FpMantRNE_48U_24U_else_carry_sva_mx0w0;
      mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs <= mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs_mx0w0;
      FpMul_8U_23U_FpMul_8U_23U_and_78_itm <= FpMul_8U_23U_FpMul_8U_23U_and_78_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_16_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= 23'b0;
    end
    else if ( core_wen & (~ or_dcpl_205) & (mux_985_nl) ) begin
      mul_loop_mul_16_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_2
          <= FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[45:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_sva_1 <= 8'b0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_15_itm <= 1'b0;
      mul_loop_mul_16_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_p_expo_and_15_cse ) begin
      FpMul_8U_23U_p_expo_sva_1 <= FpMul_8U_23U_p_expo_sva_1_mx0w0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_15_itm <= FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_15_itm_mx0w0;
      mul_loop_mul_16_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm
          <= mul_loop_mul_16_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_8_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_8_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_128_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_8_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_7_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_8_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_7_1_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_8_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_8_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_131_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_8_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_7_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_8_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_7_1_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_8_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_8_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_134_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_8_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_7_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_8_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_7_1_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_8_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_8_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_137_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_8_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_7_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_8_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_7_1_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_8_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_8_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_140_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_8_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_7_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_8_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_7_1_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_8_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_8_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_143_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_8_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_7_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_8_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_7_1_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_8_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_8_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_146_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_8_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_7_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_8_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_7_1_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_8_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_8_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_149_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_8_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_7_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_8_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_7_1_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_8_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_8_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_152_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_8_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_7_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_8_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_7_1_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_8_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_8_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_155_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_8_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_7_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_8_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_7_1_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_8_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_8_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_158_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_8_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_7_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_8_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_7_1_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_8_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_8_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_161_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_8_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_7_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_8_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_7_1_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_8_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_8_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_164_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_8_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_7_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_8_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_7_1_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_8_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_8_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_167_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_8_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_7_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_8_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_7_1_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_8_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_8_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_170_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_8_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_7_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_8_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_7_1_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_8_3_2_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_8_1_0_1 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_173_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_8_3_2_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_7_3_2_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_8_1_0_1 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_7_1_0_1;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_144_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_22_13_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_1_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_65_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_22_13, {and_dcpl_262
          , and_dcpl_266 , and_dcpl_102});
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_7_9_0_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_1_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_64_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_9_0, {and_dcpl_262
          , and_dcpl_266 , and_dcpl_102});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_1_lpi_1_dfm_5 <= 1'b0;
      IsZero_8U_23U_land_2_lpi_1_dfm_5 <= 1'b0;
      IsZero_8U_23U_land_3_lpi_1_dfm_5 <= 1'b0;
      IsZero_8U_23U_land_4_lpi_1_dfm_5 <= 1'b0;
      IsZero_8U_23U_land_5_lpi_1_dfm_5 <= 1'b0;
      IsZero_8U_23U_land_6_lpi_1_dfm_5 <= 1'b0;
      IsZero_8U_23U_land_7_lpi_1_dfm_5 <= 1'b0;
      IsZero_8U_23U_land_8_lpi_1_dfm_5 <= 1'b0;
      IsZero_8U_23U_land_9_lpi_1_dfm_5 <= 1'b0;
      IsZero_8U_23U_land_10_lpi_1_dfm_5 <= 1'b0;
      IsZero_8U_23U_land_11_lpi_1_dfm_5 <= 1'b0;
      IsZero_8U_23U_land_12_lpi_1_dfm_5 <= 1'b0;
      IsZero_8U_23U_land_13_lpi_1_dfm_5 <= 1'b0;
      IsZero_8U_23U_land_14_lpi_1_dfm_5 <= 1'b0;
      IsZero_8U_23U_land_15_lpi_1_dfm_5 <= 1'b0;
      IsZero_8U_23U_land_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_cse ) begin
      IsZero_8U_23U_land_1_lpi_1_dfm_5 <= IsZero_8U_23U_land_1_lpi_1_dfm_7;
      IsZero_8U_23U_land_2_lpi_1_dfm_5 <= IsZero_8U_23U_land_2_lpi_1_dfm_7;
      IsZero_8U_23U_land_3_lpi_1_dfm_5 <= IsZero_8U_23U_land_3_lpi_1_dfm_7;
      IsZero_8U_23U_land_4_lpi_1_dfm_5 <= IsZero_8U_23U_land_4_lpi_1_dfm_7;
      IsZero_8U_23U_land_5_lpi_1_dfm_5 <= IsZero_8U_23U_land_5_lpi_1_dfm_7;
      IsZero_8U_23U_land_6_lpi_1_dfm_5 <= IsZero_8U_23U_land_6_lpi_1_dfm_7;
      IsZero_8U_23U_land_7_lpi_1_dfm_5 <= IsZero_8U_23U_land_7_lpi_1_dfm_7;
      IsZero_8U_23U_land_8_lpi_1_dfm_5 <= IsZero_8U_23U_land_8_lpi_1_dfm_7;
      IsZero_8U_23U_land_9_lpi_1_dfm_5 <= IsZero_8U_23U_land_9_lpi_1_dfm_7;
      IsZero_8U_23U_land_10_lpi_1_dfm_5 <= IsZero_8U_23U_land_10_lpi_1_dfm_7;
      IsZero_8U_23U_land_11_lpi_1_dfm_5 <= IsZero_8U_23U_land_11_lpi_1_dfm_7;
      IsZero_8U_23U_land_12_lpi_1_dfm_5 <= IsZero_8U_23U_land_12_lpi_1_dfm_7;
      IsZero_8U_23U_land_13_lpi_1_dfm_5 <= IsZero_8U_23U_land_13_lpi_1_dfm_7;
      IsZero_8U_23U_land_14_lpi_1_dfm_5 <= IsZero_8U_23U_land_14_lpi_1_dfm_7;
      IsZero_8U_23U_land_15_lpi_1_dfm_5 <= IsZero_8U_23U_land_15_lpi_1_dfm_7;
      IsZero_8U_23U_land_lpi_1_dfm_5 <= IsZero_8U_23U_land_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_1_land_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1140_nl))
        ) begin
      IsZero_8U_23U_1_land_1_lpi_1_dfm_6 <= MUX_s_1_2_2(IsZero_8U_23U_1_land_1_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_1_land_1_lpi_1_dfm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_else_2_if_and_cse & (~ or_dcpl_217) & (~ (mux_1144_nl))
        ) begin
      mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= mul_loop_mul_1_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_18_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_217) ) begin
      FpMul_8U_23U_lor_18_lpi_1_dfm_st <= or_312_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_147_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_22_13_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_2_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_68_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_22_13, {and_dcpl_277
          , and_dcpl_281 , and_dcpl_108});
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_7_9_0_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_2_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_67_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_9_0, {and_dcpl_277
          , and_dcpl_281 , and_dcpl_108});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_1_land_2_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1162_nl))
        ) begin
      IsZero_8U_23U_1_land_2_lpi_1_dfm_6 <= MUX_s_1_2_2(IsZero_8U_23U_1_land_2_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_1_land_2_lpi_1_dfm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_else_2_if_and_cse & (~ or_dcpl_227) & (~ (mux_1167_nl))
        ) begin
      mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= mul_loop_mul_2_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_19_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_227) ) begin
      FpMul_8U_23U_lor_19_lpi_1_dfm_st <= or_2628_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_150_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_22_13_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_3_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_71_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_22_13, {and_dcpl_292
          , and_dcpl_296 , and_dcpl_112});
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_7_9_0_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_3_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_70_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_9_0, {and_dcpl_292
          , and_dcpl_296 , and_dcpl_112});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_1_land_3_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1185_nl))
        ) begin
      IsZero_8U_23U_1_land_3_lpi_1_dfm_6 <= MUX_s_1_2_2(IsZero_8U_23U_1_land_3_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_1_land_3_lpi_1_dfm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_else_2_if_and_cse & (~ or_dcpl_237) & (~ (mux_1189_nl))
        ) begin
      mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= mul_loop_mul_3_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_20_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_237) ) begin
      FpMul_8U_23U_lor_20_lpi_1_dfm_st <= or_363_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_153_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_22_13_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_4_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_74_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_22_13, {and_dcpl_307
          , and_dcpl_311 , and_dcpl_116});
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_7_9_0_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_4_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_73_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_9_0, {and_dcpl_307
          , and_dcpl_311 , and_dcpl_116});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_1_land_4_lpi_1_dfm_4 <= 1'b0;
      IsZero_8U_23U_1_land_6_lpi_1_dfm_4 <= 1'b0;
      IsZero_8U_23U_1_land_7_lpi_1_dfm_4 <= 1'b0;
      IsZero_8U_23U_1_land_10_lpi_1_dfm_4 <= 1'b0;
      IsZero_8U_23U_1_land_11_lpi_1_dfm_4 <= 1'b0;
      IsZero_8U_23U_1_land_12_lpi_1_dfm_4 <= 1'b0;
      IsZero_8U_23U_1_land_14_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( IsZero_8U_23U_1_aelse_and_cse ) begin
      IsZero_8U_23U_1_land_4_lpi_1_dfm_4 <= MUX_s_1_2_2(IsZero_8U_23U_1_land_4_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_1_land_4_lpi_1_dfm, and_dcpl_104);
      IsZero_8U_23U_1_land_6_lpi_1_dfm_4 <= MUX_s_1_2_2(IsZero_8U_23U_1_land_6_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_1_land_6_lpi_1_dfm, and_dcpl_104);
      IsZero_8U_23U_1_land_7_lpi_1_dfm_4 <= MUX_s_1_2_2(IsZero_8U_23U_1_land_7_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_1_land_7_lpi_1_dfm, and_dcpl_104);
      IsZero_8U_23U_1_land_10_lpi_1_dfm_4 <= MUX_s_1_2_2(IsZero_8U_23U_1_land_10_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_1_land_10_lpi_1_dfm, and_dcpl_104);
      IsZero_8U_23U_1_land_11_lpi_1_dfm_4 <= MUX_s_1_2_2(IsZero_8U_23U_1_land_11_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_1_land_11_lpi_1_dfm, and_dcpl_104);
      IsZero_8U_23U_1_land_12_lpi_1_dfm_4 <= MUX_s_1_2_2(IsZero_8U_23U_1_land_12_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_1_land_12_lpi_1_dfm, and_dcpl_104);
      IsZero_8U_23U_1_land_14_lpi_1_dfm_4 <= MUX_s_1_2_2(IsZero_8U_23U_1_land_14_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_1_land_14_lpi_1_dfm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_else_2_if_and_cse & (~ or_dcpl_247) & (~ (mux_1194_nl))
        ) begin
      mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= mul_loop_mul_4_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_21_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_247) ) begin
      FpMul_8U_23U_lor_21_lpi_1_dfm_st <= or_386_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_156_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_22_13_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_5_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_77_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_22_13, {and_dcpl_322
          , and_dcpl_326 , and_dcpl_120});
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_7_9_0_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_5_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_76_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_9_0, {and_dcpl_322
          , and_dcpl_326 , and_dcpl_120});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_1_land_5_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1212_nl))
        ) begin
      IsZero_8U_23U_1_land_5_lpi_1_dfm_6 <= MUX_s_1_2_2(IsZero_8U_23U_1_land_5_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_1_land_5_lpi_1_dfm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_else_2_if_and_cse & (~ or_dcpl_257) & (~ (mux_1218_nl))
        ) begin
      mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= mul_loop_mul_5_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_22_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_257) ) begin
      FpMul_8U_23U_lor_22_lpi_1_dfm_st <= FpMul_8U_23U_lor_22_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_159_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_22_13_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_6_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_80_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_22_13, {and_dcpl_337
          , and_dcpl_341 , and_dcpl_124});
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_7_9_0_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_6_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_79_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_9_0, {and_dcpl_337
          , and_dcpl_341 , and_dcpl_124});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_else_2_if_and_cse & (~ or_dcpl_267) & (~ (mux_1223_nl))
        ) begin
      mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= mul_loop_mul_6_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_23_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_267) ) begin
      FpMul_8U_23U_lor_23_lpi_1_dfm_st <= or_438_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_162_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_22_13_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_7_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_83_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_22_13, {and_dcpl_352
          , and_dcpl_356 , and_dcpl_128});
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_7_9_0_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_7_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_82_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_9_0, {and_dcpl_352
          , and_dcpl_356 , and_dcpl_128});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_else_2_if_and_cse & (~ or_dcpl_277) & (~ (mux_1228_nl))
        ) begin
      mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= mul_loop_mul_7_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_24_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_277) ) begin
      FpMul_8U_23U_lor_24_lpi_1_dfm_st <= or_461_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_165_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_22_13_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_8_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_86_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_22_13, {and_dcpl_367
          , and_dcpl_371 , and_dcpl_132});
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_7_9_0_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_8_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_85_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_9_0, {and_dcpl_367
          , and_dcpl_371 , and_dcpl_132});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_1_land_8_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1246_nl))
        ) begin
      IsZero_8U_23U_1_land_8_lpi_1_dfm_6 <= MUX_s_1_2_2(IsZero_8U_23U_1_land_8_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_1_land_8_lpi_1_dfm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_else_2_if_and_cse & (~ or_dcpl_287) & (~ (mux_1251_nl))
        ) begin
      mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= mul_loop_mul_8_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_25_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_287) ) begin
      FpMul_8U_23U_lor_25_lpi_1_dfm_st <= or_2742_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_168_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_22_13_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_9_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_89_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_22_13, {and_dcpl_382
          , and_dcpl_386 , and_dcpl_136});
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_7_9_0_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_9_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_88_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_9_0, {and_dcpl_382
          , and_dcpl_386 , and_dcpl_136});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_1_land_9_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1269_nl))
        ) begin
      IsZero_8U_23U_1_land_9_lpi_1_dfm_6 <= MUX_s_1_2_2(IsZero_8U_23U_1_land_9_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_1_land_9_lpi_1_dfm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_else_2_if_and_cse & (~ or_dcpl_297) & (~ (mux_1275_nl))
        ) begin
      mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= mul_loop_mul_9_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_26_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_297) ) begin
      FpMul_8U_23U_lor_26_lpi_1_dfm_st <= FpMul_8U_23U_lor_26_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_171_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_22_13_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_10_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_92_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_22_13, {and_dcpl_397
          , and_dcpl_401 , and_dcpl_140});
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_7_9_0_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_10_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_91_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_9_0, {and_dcpl_397
          , and_dcpl_401 , and_dcpl_140});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_else_2_if_and_cse & (~ or_dcpl_307) & (~ (mux_1280_nl))
        ) begin
      mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= mul_loop_mul_10_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_27_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_307) ) begin
      FpMul_8U_23U_lor_27_lpi_1_dfm_st <= FpMul_8U_23U_lor_27_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_174_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_22_13_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_11_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_95_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_22_13, {and_dcpl_412
          , and_dcpl_416 , and_dcpl_144});
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_7_9_0_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_11_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_94_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_9_0, {and_dcpl_412
          , and_dcpl_416 , and_dcpl_144});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_else_2_if_and_cse & (~ or_dcpl_317) & (~ (mux_1285_nl))
        ) begin
      mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= mul_loop_mul_11_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_28_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_317) ) begin
      FpMul_8U_23U_lor_28_lpi_1_dfm_st <= or_570_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_177_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_22_13_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_12_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_98_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_22_13, {and_dcpl_427
          , and_dcpl_431 , and_dcpl_148});
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_7_9_0_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_12_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_97_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_9_0, {and_dcpl_427
          , and_dcpl_431 , and_dcpl_148});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_else_2_if_and_cse & (~ or_dcpl_327) & (~ (mux_1290_nl))
        ) begin
      mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= mul_loop_mul_12_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_29_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_327) ) begin
      FpMul_8U_23U_lor_29_lpi_1_dfm_st <= or_593_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_180_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_22_13_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_13_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_101_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_22_13, {and_dcpl_442
          , and_dcpl_446 , and_dcpl_152});
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_7_9_0_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_13_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_100_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_9_0, {and_dcpl_442
          , and_dcpl_446 , and_dcpl_152});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_1_land_13_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1308_nl))
        ) begin
      IsZero_8U_23U_1_land_13_lpi_1_dfm_6 <= MUX_s_1_2_2(IsZero_8U_23U_1_land_13_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_1_land_13_lpi_1_dfm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_else_2_if_and_cse & (~ or_dcpl_337) & (~ (mux_1313_nl))
        ) begin
      mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= mul_loop_mul_13_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_30_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_337) ) begin
      FpMul_8U_23U_lor_30_lpi_1_dfm_st <= or_616_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_183_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_22_13_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_14_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_104_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_22_13, {and_dcpl_457
          , and_dcpl_461 , and_dcpl_156});
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_7_9_0_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_14_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_103_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_9_0, {and_dcpl_457
          , and_dcpl_461 , and_dcpl_156});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_else_2_if_and_cse & (~ or_dcpl_347) & (~ (mux_1318_nl))
        ) begin
      mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= mul_loop_mul_14_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_31_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_347) ) begin
      FpMul_8U_23U_lor_31_lpi_1_dfm_st <= or_639_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_186_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_22_13_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_15_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_107_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_22_13, {and_dcpl_472
          , and_dcpl_476 , and_dcpl_160});
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_7_9_0_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_15_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_106_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_9_0, {and_dcpl_472
          , and_dcpl_476 , and_dcpl_160});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_1_land_15_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1336_nl))
        ) begin
      IsZero_8U_23U_1_land_15_lpi_1_dfm_6 <= MUX_s_1_2_2(IsZero_8U_23U_1_land_15_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_1_land_15_lpi_1_dfm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_else_2_if_and_cse & (~ or_dcpl_357) & (~ (mux_1340_nl))
        ) begin
      mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= mul_loop_mul_15_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_32_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_357) ) begin
      FpMul_8U_23U_lor_32_lpi_1_dfm_st <= or_662_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_22_13_1 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_9_0_1 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_189_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_22_13_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_110_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_22_13, {and_dcpl_487
          , and_dcpl_491 , and_dcpl_164});
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_7_9_0_1 <= MUX1HOT_v_10_3_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_109_mx0w1,
          FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_9_0, {and_dcpl_487 ,
          and_dcpl_491 , and_dcpl_164});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_1_land_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1358_nl))
        ) begin
      IsZero_8U_23U_1_land_lpi_1_dfm_6 <= MUX_s_1_2_2(IsZero_8U_23U_1_land_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_1_land_lpi_1_dfm, and_dcpl_104);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= 1'b0;
    end
    else if ( FpMul_8U_23U_else_2_if_and_cse & (~ or_dcpl_367) & (~ (mux_1363_nl))
        ) begin
      mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st
          <= mul_loop_mul_16_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_1_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_367) ) begin
      FpMul_8U_23U_lor_1_lpi_1_dfm_st <= or_2885_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_3_2 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_1_0 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3 <= 4'b0;
      FpMul_8U_23U_lor_3_lpi_1_dfm_st <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_12_10 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_3_2 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_3_2_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_1_0 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_1_0_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w0;
      FpMul_8U_23U_lor_3_lpi_1_dfm_st <= FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_tmp;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_12_10_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_3_2 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_1_0 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3 <= 4'b0;
      FpMul_8U_23U_lor_4_lpi_1_dfm_st <= 1'b0;
      IsZero_8U_23U_1_land_2_lpi_1_dfm <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_12_10 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_3_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_3_2 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_3_2_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_1_0 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_1_0_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w0;
      FpMul_8U_23U_lor_4_lpi_1_dfm_st <= FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_2_tmp;
      IsZero_8U_23U_1_land_2_lpi_1_dfm <= IsZero_8U_23U_1_land_2_lpi_1_dfm_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_12_10_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_3_2 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_1_0 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3 <= 4'b0;
      FpMul_8U_23U_lor_5_lpi_1_dfm_st <= 1'b0;
      IsZero_8U_23U_1_land_3_lpi_1_dfm <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_12_10 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_6_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_3_2 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_3_2_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_1_0 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_1_0_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w0;
      FpMul_8U_23U_lor_5_lpi_1_dfm_st <= FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_4_tmp;
      IsZero_8U_23U_1_land_3_lpi_1_dfm <= IsZero_8U_23U_1_land_3_lpi_1_dfm_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_12_10_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_3_2 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_1_0 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3 <= 4'b0;
      FpMul_8U_23U_lor_6_lpi_1_dfm_st <= 1'b0;
      IsZero_8U_23U_1_land_4_lpi_1_dfm <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_12_10 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_9_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_3_2 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_3_2_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_1_0 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_1_0_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3_mx0w0;
      FpMul_8U_23U_lor_6_lpi_1_dfm_st <= FpMul_8U_23U_lor_6_lpi_1_dfm_mx0w0;
      IsZero_8U_23U_1_land_4_lpi_1_dfm <= IsZero_8U_23U_1_land_4_lpi_1_dfm_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_12_10_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_3_2 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_1_0 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3 <= 4'b0;
      FpMul_8U_23U_lor_7_lpi_1_dfm_st <= 1'b0;
      IsZero_8U_23U_1_land_5_lpi_1_dfm <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_12_10 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_12_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_3_2 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_3_2_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_1_0 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_1_0_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3_mx0w0;
      FpMul_8U_23U_lor_7_lpi_1_dfm_st <= FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_8_tmp;
      IsZero_8U_23U_1_land_5_lpi_1_dfm <= IsZero_8U_23U_1_land_5_lpi_1_dfm_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_12_10_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_3_2 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_1_0 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3 <= 4'b0;
      FpMul_8U_23U_lor_8_lpi_1_dfm_st <= 1'b0;
      IsZero_8U_23U_1_land_6_lpi_1_dfm <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_12_10 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_15_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_3_2 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_3_2_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_1_0 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_1_0_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3_mx0w0;
      FpMul_8U_23U_lor_8_lpi_1_dfm_st <= FpMul_8U_23U_lor_8_lpi_1_dfm_mx0w0;
      IsZero_8U_23U_1_land_6_lpi_1_dfm <= IsZero_8U_23U_1_land_6_lpi_1_dfm_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_12_10_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_3_2 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_1_0 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3 <= 4'b0;
      FpMul_8U_23U_lor_9_lpi_1_dfm_st <= 1'b0;
      IsZero_8U_23U_1_land_7_lpi_1_dfm <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_12_10 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_18_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_3_2 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_3_2_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_1_0 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_1_0_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3_mx0w0;
      FpMul_8U_23U_lor_9_lpi_1_dfm_st <= FpMul_8U_23U_lor_9_lpi_1_dfm_mx0w0;
      IsZero_8U_23U_1_land_7_lpi_1_dfm <= IsZero_8U_23U_1_land_7_lpi_1_dfm_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_12_10_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_3_2 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_1_0 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3 <= 4'b0;
      FpMul_8U_23U_lor_10_lpi_1_dfm_st <= 1'b0;
      IsZero_8U_23U_1_land_8_lpi_1_dfm <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_12_10 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_21_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_3_2 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_3_2_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_1_0 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_1_0_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3_mx0w0;
      FpMul_8U_23U_lor_10_lpi_1_dfm_st <= FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_14_tmp;
      IsZero_8U_23U_1_land_8_lpi_1_dfm <= IsZero_8U_23U_1_land_8_lpi_1_dfm_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_12_10_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_3_2 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_1_0 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3 <= 4'b0;
      FpMul_8U_23U_lor_11_lpi_1_dfm_st <= 1'b0;
      IsZero_8U_23U_1_land_9_lpi_1_dfm <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_12_10 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_24_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_3_2 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_3_2_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_1_0 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_1_0_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3_mx0w0;
      FpMul_8U_23U_lor_11_lpi_1_dfm_st <= FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_16_tmp;
      IsZero_8U_23U_1_land_9_lpi_1_dfm <= IsZero_8U_23U_1_land_9_lpi_1_dfm_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_12_10_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_3_2 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_1_0 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3 <= 4'b0;
      FpMul_8U_23U_lor_12_lpi_1_dfm_st <= 1'b0;
      IsZero_8U_23U_1_land_10_lpi_1_dfm <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_12_10 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_27_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_3_2 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_3_2_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_1_0 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_1_0_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3_mx0w0;
      FpMul_8U_23U_lor_12_lpi_1_dfm_st <= FpMul_8U_23U_lor_12_lpi_1_dfm_mx0w0;
      IsZero_8U_23U_1_land_10_lpi_1_dfm <= IsZero_8U_23U_1_land_10_lpi_1_dfm_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_12_10_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_3_2 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_1_0 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3 <= 4'b0;
      FpMul_8U_23U_lor_13_lpi_1_dfm_st <= 1'b0;
      IsZero_8U_23U_1_land_11_lpi_1_dfm <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_12_10 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_30_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_3_2 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_3_2_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_1_0 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_1_0_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3_mx0w0;
      FpMul_8U_23U_lor_13_lpi_1_dfm_st <= FpMul_8U_23U_lor_13_lpi_1_dfm_mx0w0;
      IsZero_8U_23U_1_land_11_lpi_1_dfm <= IsZero_8U_23U_1_land_11_lpi_1_dfm_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_12_10_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_3_2 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_1_0 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3 <= 4'b0;
      FpMul_8U_23U_lor_14_lpi_1_dfm_st <= 1'b0;
      IsZero_8U_23U_1_land_12_lpi_1_dfm <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_12_10 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_33_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_3_2 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_3_2_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_1_0 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_1_0_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3_mx0w0;
      FpMul_8U_23U_lor_14_lpi_1_dfm_st <= FpMul_8U_23U_lor_14_lpi_1_dfm_mx0w0;
      IsZero_8U_23U_1_land_12_lpi_1_dfm <= IsZero_8U_23U_1_land_12_lpi_1_dfm_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_12_10_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_3_2 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_1_0 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3 <= 4'b0;
      FpMul_8U_23U_lor_15_lpi_1_dfm_st <= 1'b0;
      IsZero_8U_23U_1_land_13_lpi_1_dfm <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_12_10 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_36_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_3_2 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_3_2_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_1_0 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_1_0_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3_mx0w0;
      FpMul_8U_23U_lor_15_lpi_1_dfm_st <= FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_24_tmp;
      IsZero_8U_23U_1_land_13_lpi_1_dfm <= IsZero_8U_23U_1_land_13_lpi_1_dfm_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_12_10_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_3_2 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_1_0 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3 <= 4'b0;
      FpMul_8U_23U_lor_16_lpi_1_dfm_st <= 1'b0;
      IsZero_8U_23U_1_land_14_lpi_1_dfm <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_12_10 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_39_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_3_2 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_3_2_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_1_0 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_1_0_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3_mx0w0;
      FpMul_8U_23U_lor_16_lpi_1_dfm_st <= FpMul_8U_23U_lor_16_lpi_1_dfm_mx0w0;
      IsZero_8U_23U_1_land_14_lpi_1_dfm <= IsZero_8U_23U_1_land_14_lpi_1_dfm_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_12_10_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_3_2 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_1_0 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3 <= 4'b0;
      FpMul_8U_23U_lor_17_lpi_1_dfm_st <= 1'b0;
      IsZero_8U_23U_1_land_15_lpi_1_dfm <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_12_10 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_42_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_3_2 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_3_2_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_1_0 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_1_0_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3_mx0w0;
      FpMul_8U_23U_lor_17_lpi_1_dfm_st <= FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_28_tmp;
      IsZero_8U_23U_1_land_15_lpi_1_dfm <= IsZero_8U_23U_1_land_15_lpi_1_dfm_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_12_10_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_3_2 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_1_0 <= 2'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3 <= 4'b0;
      FpMul_8U_23U_lor_lpi_1_dfm_st <= 1'b0;
      IsZero_8U_23U_1_land_lpi_1_dfm <= 1'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_12_10 <= 3'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_and_45_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_3_2 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_3_2_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_1_0 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_1_0_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w0;
      FpMul_8U_23U_lor_lpi_1_dfm_st <= FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_30_tmp;
      IsZero_8U_23U_1_land_lpi_1_dfm <= IsZero_8U_23U_1_land_lpi_1_dfm_mx0w0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_12_10 <= FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_12_10_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_if_land_lpi_1_dfm_st <= 1'b0;
      mul_loop_mul_if_land_15_lpi_1_dfm_st <= 1'b0;
      mul_loop_mul_if_land_14_lpi_1_dfm_st <= 1'b0;
      mul_loop_mul_if_land_13_lpi_1_dfm_st <= 1'b0;
      mul_loop_mul_if_land_12_lpi_1_dfm_st <= 1'b0;
      mul_loop_mul_if_land_11_lpi_1_dfm_st <= 1'b0;
      mul_loop_mul_if_land_10_lpi_1_dfm_st <= 1'b0;
      mul_loop_mul_if_land_9_lpi_1_dfm_st <= 1'b0;
      mul_loop_mul_if_land_8_lpi_1_dfm_st <= 1'b0;
      mul_loop_mul_if_land_7_lpi_1_dfm_st <= 1'b0;
      mul_loop_mul_if_land_6_lpi_1_dfm_st <= 1'b0;
      mul_loop_mul_if_land_5_lpi_1_dfm_st <= 1'b0;
      mul_loop_mul_if_land_4_lpi_1_dfm_st <= 1'b0;
      mul_loop_mul_if_land_3_lpi_1_dfm_st <= 1'b0;
      mul_loop_mul_if_land_2_lpi_1_dfm_st <= 1'b0;
      mul_loop_mul_if_land_1_lpi_1_dfm_st <= 1'b0;
    end
    else if ( mul_loop_mul_if_aelse_and_cse ) begin
      mul_loop_mul_if_land_lpi_1_dfm_st <= nor_44_cse;
      mul_loop_mul_if_land_15_lpi_1_dfm_st <= nor_42_cse;
      mul_loop_mul_if_land_14_lpi_1_dfm_st <= nor_40_cse;
      mul_loop_mul_if_land_13_lpi_1_dfm_st <= nor_39_cse;
      mul_loop_mul_if_land_12_lpi_1_dfm_st <= nor_37_cse;
      mul_loop_mul_if_land_11_lpi_1_dfm_st <= nor_36_cse;
      mul_loop_mul_if_land_10_lpi_1_dfm_st <= nor_35_cse;
      mul_loop_mul_if_land_9_lpi_1_dfm_st <= nor_34_cse;
      mul_loop_mul_if_land_8_lpi_1_dfm_st <= nor_32_cse;
      mul_loop_mul_if_land_7_lpi_1_dfm_st <= nor_30_cse;
      mul_loop_mul_if_land_6_lpi_1_dfm_st <= nor_29_cse;
      mul_loop_mul_if_land_5_lpi_1_dfm_st <= nor_28_cse;
      mul_loop_mul_if_land_4_lpi_1_dfm_st <= nor_26_cse;
      mul_loop_mul_if_land_3_lpi_1_dfm_st <= nor_25_cse;
      mul_loop_mul_if_land_2_lpi_1_dfm_st <= nor_23_cse;
      mul_loop_mul_if_land_1_lpi_1_dfm_st <= nor_21_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_mul_src_1_sva_st <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_53 | and_dcpl_50 | or_dcpl_31 | (fsm_output[0])))
        ) begin
      cfg_mul_src_1_sva_st <= cfg_mul_src_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulIn_data_sva_533 <= 528'b0;
      mul_loop_mul_if_land_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_if_land_15_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_if_land_14_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_if_land_13_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_if_land_12_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_if_land_11_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_if_land_10_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_if_land_9_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_if_land_8_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_if_land_7_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_if_land_6_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_if_land_5_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_if_land_4_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_if_land_3_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_if_land_2_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_if_land_1_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_else_land_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_else_land_15_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_else_land_14_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_else_land_13_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_else_land_12_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_else_land_11_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_else_land_10_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_else_land_9_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_else_land_8_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_else_land_7_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_else_land_6_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_else_land_5_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_else_land_4_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_else_land_3_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_else_land_2_lpi_1_dfm_7 <= 1'b0;
      mul_loop_mul_else_land_1_lpi_1_dfm_7 <= 1'b0;
      io_read_cfg_mul_bypass_rsc_svs_5 <= 1'b0;
    end
    else if ( MulIn_data_and_3_cse ) begin
      MulIn_data_sva_533 <= chn_mul_in_rsci_d_mxwt;
      mul_loop_mul_if_land_lpi_1_dfm_7 <= nor_44_cse;
      mul_loop_mul_if_land_15_lpi_1_dfm_7 <= nor_42_cse;
      mul_loop_mul_if_land_14_lpi_1_dfm_7 <= nor_40_cse;
      mul_loop_mul_if_land_13_lpi_1_dfm_7 <= nor_39_cse;
      mul_loop_mul_if_land_12_lpi_1_dfm_7 <= nor_37_cse;
      mul_loop_mul_if_land_11_lpi_1_dfm_7 <= nor_36_cse;
      mul_loop_mul_if_land_10_lpi_1_dfm_7 <= nor_35_cse;
      mul_loop_mul_if_land_9_lpi_1_dfm_7 <= nor_34_cse;
      mul_loop_mul_if_land_8_lpi_1_dfm_7 <= nor_32_cse;
      mul_loop_mul_if_land_7_lpi_1_dfm_7 <= nor_30_cse;
      mul_loop_mul_if_land_6_lpi_1_dfm_7 <= nor_29_cse;
      mul_loop_mul_if_land_5_lpi_1_dfm_7 <= nor_28_cse;
      mul_loop_mul_if_land_4_lpi_1_dfm_7 <= nor_26_cse;
      mul_loop_mul_if_land_3_lpi_1_dfm_7 <= nor_25_cse;
      mul_loop_mul_if_land_2_lpi_1_dfm_7 <= nor_23_cse;
      mul_loop_mul_if_land_1_lpi_1_dfm_7 <= nor_21_cse;
      mul_loop_mul_else_land_lpi_1_dfm_7 <= ~((chn_mul_in_rsci_d_mxwt[527]) | (~
          cfg_mul_prelu_rsci_d));
      mul_loop_mul_else_land_15_lpi_1_dfm_7 <= ~((chn_mul_in_rsci_d_mxwt[494]) |
          (~ cfg_mul_prelu_rsci_d));
      mul_loop_mul_else_land_14_lpi_1_dfm_7 <= ~((chn_mul_in_rsci_d_mxwt[461]) |
          (~ cfg_mul_prelu_rsci_d));
      mul_loop_mul_else_land_13_lpi_1_dfm_7 <= ~((chn_mul_in_rsci_d_mxwt[428]) |
          (~ cfg_mul_prelu_rsci_d));
      mul_loop_mul_else_land_12_lpi_1_dfm_7 <= ~((chn_mul_in_rsci_d_mxwt[395]) |
          (~ cfg_mul_prelu_rsci_d));
      mul_loop_mul_else_land_11_lpi_1_dfm_7 <= ~((chn_mul_in_rsci_d_mxwt[362]) |
          (~ cfg_mul_prelu_rsci_d));
      mul_loop_mul_else_land_10_lpi_1_dfm_7 <= ~((chn_mul_in_rsci_d_mxwt[329]) |
          (~ cfg_mul_prelu_rsci_d));
      mul_loop_mul_else_land_9_lpi_1_dfm_7 <= ~((chn_mul_in_rsci_d_mxwt[296]) | (~
          cfg_mul_prelu_rsci_d));
      mul_loop_mul_else_land_8_lpi_1_dfm_7 <= ~((chn_mul_in_rsci_d_mxwt[263]) | (~
          cfg_mul_prelu_rsci_d));
      mul_loop_mul_else_land_7_lpi_1_dfm_7 <= ~((chn_mul_in_rsci_d_mxwt[230]) | (~
          cfg_mul_prelu_rsci_d));
      mul_loop_mul_else_land_6_lpi_1_dfm_7 <= ~((chn_mul_in_rsci_d_mxwt[197]) | (~
          cfg_mul_prelu_rsci_d));
      mul_loop_mul_else_land_5_lpi_1_dfm_7 <= ~((chn_mul_in_rsci_d_mxwt[164]) | (~
          cfg_mul_prelu_rsci_d));
      mul_loop_mul_else_land_4_lpi_1_dfm_7 <= ~((chn_mul_in_rsci_d_mxwt[131]) | (~
          cfg_mul_prelu_rsci_d));
      mul_loop_mul_else_land_3_lpi_1_dfm_7 <= ~((chn_mul_in_rsci_d_mxwt[98]) | (~
          cfg_mul_prelu_rsci_d));
      mul_loop_mul_else_land_2_lpi_1_dfm_7 <= ~((chn_mul_in_rsci_d_mxwt[65]) | (~
          cfg_mul_prelu_rsci_d));
      mul_loop_mul_else_land_1_lpi_1_dfm_7 <= ~((chn_mul_in_rsci_d_mxwt[32]) | (~
          cfg_mul_prelu_rsci_d));
      io_read_cfg_mul_bypass_rsc_svs_5 <= cfg_mul_bypass_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_1_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_48_cse ) begin
      IsZero_8U_23U_land_1_lpi_1_dfm_7 <= MUX_s_1_2_2(IsZero_8U_23U_land_1_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_land_1_lpi_1_dfm, and_dcpl_497);
      IsNaN_8U_23U_land_1_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_land_1_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_1_lpi_1_dfm, and_dcpl_497);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_2_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_49_cse ) begin
      IsZero_8U_23U_land_2_lpi_1_dfm_7 <= MUX_s_1_2_2(IsZero_8U_23U_land_2_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_land_2_lpi_1_dfm, and_dcpl_500);
      IsNaN_8U_23U_land_2_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_land_2_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_2_lpi_1_dfm, and_dcpl_500);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_3_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_50_cse ) begin
      IsZero_8U_23U_land_3_lpi_1_dfm_7 <= MUX_s_1_2_2(IsZero_8U_23U_land_3_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_land_3_lpi_1_dfm, and_dcpl_503);
      IsNaN_8U_23U_land_3_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_land_3_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_3_lpi_1_dfm, and_dcpl_503);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_4_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_land_4_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_51_cse ) begin
      IsZero_8U_23U_land_4_lpi_1_dfm_7 <= MUX_s_1_2_2(IsZero_8U_23U_land_4_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_land_4_lpi_1_dfm, and_dcpl_506);
      IsNaN_8U_23U_land_4_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_land_4_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_4_lpi_1_dfm, and_dcpl_506);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_5_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_land_5_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_52_cse ) begin
      IsZero_8U_23U_land_5_lpi_1_dfm_7 <= MUX_s_1_2_2(IsZero_8U_23U_land_5_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_land_5_lpi_1_dfm, and_dcpl_509);
      IsNaN_8U_23U_land_5_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_land_5_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_5_lpi_1_dfm, and_dcpl_509);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_6_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_land_6_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_53_cse ) begin
      IsZero_8U_23U_land_6_lpi_1_dfm_7 <= MUX_s_1_2_2(IsZero_8U_23U_land_6_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_land_6_lpi_1_dfm, and_dcpl_512);
      IsNaN_8U_23U_land_6_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_land_6_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_6_lpi_1_dfm, and_dcpl_512);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_7_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_land_7_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_54_cse ) begin
      IsZero_8U_23U_land_7_lpi_1_dfm_7 <= MUX_s_1_2_2(IsZero_8U_23U_land_7_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_land_7_lpi_1_dfm, and_dcpl_515);
      IsNaN_8U_23U_land_7_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_land_7_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_7_lpi_1_dfm, and_dcpl_515);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_8_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_land_8_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_55_cse ) begin
      IsZero_8U_23U_land_8_lpi_1_dfm_7 <= MUX_s_1_2_2(IsZero_8U_23U_land_8_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_land_8_lpi_1_dfm, and_dcpl_518);
      IsNaN_8U_23U_land_8_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_land_8_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_8_lpi_1_dfm, and_dcpl_518);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_9_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_land_9_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_56_cse ) begin
      IsZero_8U_23U_land_9_lpi_1_dfm_7 <= MUX_s_1_2_2(IsZero_8U_23U_land_9_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_land_9_lpi_1_dfm, and_dcpl_521);
      IsNaN_8U_23U_land_9_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_land_9_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_9_lpi_1_dfm, and_dcpl_521);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_10_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_land_10_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_57_cse ) begin
      IsZero_8U_23U_land_10_lpi_1_dfm_7 <= MUX_s_1_2_2(IsZero_8U_23U_land_10_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_land_10_lpi_1_dfm, and_dcpl_524);
      IsNaN_8U_23U_land_10_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_land_10_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_10_lpi_1_dfm, and_dcpl_524);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_11_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_land_11_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_58_cse ) begin
      IsZero_8U_23U_land_11_lpi_1_dfm_7 <= MUX_s_1_2_2(IsZero_8U_23U_land_11_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_land_11_lpi_1_dfm, and_dcpl_527);
      IsNaN_8U_23U_land_11_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_land_11_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_11_lpi_1_dfm, and_dcpl_527);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_12_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_land_12_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_59_cse ) begin
      IsZero_8U_23U_land_12_lpi_1_dfm_7 <= MUX_s_1_2_2(IsZero_8U_23U_land_12_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_land_12_lpi_1_dfm, and_dcpl_530);
      IsNaN_8U_23U_land_12_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_land_12_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_12_lpi_1_dfm, and_dcpl_530);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_13_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_land_13_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_60_cse ) begin
      IsZero_8U_23U_land_13_lpi_1_dfm_7 <= MUX_s_1_2_2(IsZero_8U_23U_land_13_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_land_13_lpi_1_dfm, and_dcpl_533);
      IsNaN_8U_23U_land_13_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_land_13_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_13_lpi_1_dfm, and_dcpl_533);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_14_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_land_14_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_61_cse ) begin
      IsZero_8U_23U_land_14_lpi_1_dfm_7 <= MUX_s_1_2_2(IsZero_8U_23U_land_14_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_land_14_lpi_1_dfm, and_dcpl_536);
      IsNaN_8U_23U_land_14_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_land_14_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_14_lpi_1_dfm, and_dcpl_536);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_15_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_land_15_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_62_cse ) begin
      IsZero_8U_23U_land_15_lpi_1_dfm_7 <= MUX_s_1_2_2(IsZero_8U_23U_land_15_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_land_15_lpi_1_dfm, and_dcpl_539);
      IsNaN_8U_23U_land_15_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_land_15_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_15_lpi_1_dfm, and_dcpl_539);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_63_cse ) begin
      IsZero_8U_23U_land_lpi_1_dfm_7 <= MUX_s_1_2_2(IsZero_8U_23U_land_lpi_1_dfm_mx0w0,
          IsZero_8U_23U_land_lpi_1_dfm, and_dcpl_542);
      IsNaN_8U_23U_land_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_8U_23U_land_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_lpi_1_dfm, and_dcpl_542);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1446_nl))
        ) begin
      FpMul_8U_23U_lor_1_lpi_1_dfm_6 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_16_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1447_nl)) ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_252_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_1108_rgt | and_1111_rgt | and_1112_rgt) & (~ (mux_1448_nl))
        ) begin
      FpMul_8U_23U_mux_252_itm_3 <= MUX1HOT_s_1_3_2((MulIn_data_sva_534[526]), FpMul_8U_23U_else_5_mux_60_mx0w1,
          FpMul_8U_23U_mux_252_itm, {and_1108_rgt , and_1111_rgt , and_1112_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_32_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1449_nl))
        ) begin
      FpMul_8U_23U_lor_32_lpi_1_dfm_6 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_17_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_15_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1450_nl)) ) begin
      IsNaN_8U_23U_1_land_15_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_15_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_236_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_1117_rgt | and_1120_rgt | and_1121_rgt) & (~ (mux_1452_nl))
        ) begin
      FpMul_8U_23U_mux_236_itm_3 <= MUX1HOT_s_1_3_2((MulIn_data_sva_534[493]), FpMul_8U_23U_else_5_mux_56_mx0w1,
          FpMul_8U_23U_mux_236_itm, {and_1117_rgt , and_1120_rgt , and_1121_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_31_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1453_nl))
        ) begin
      FpMul_8U_23U_lor_31_lpi_1_dfm_6 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_18_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_14_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1454_nl)) ) begin
      IsNaN_8U_23U_1_land_14_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_14_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_220_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_1126_rgt | and_1129_rgt | and_1130_rgt) & (~ (mux_1456_nl))
        ) begin
      FpMul_8U_23U_mux_220_itm_3 <= MUX1HOT_s_1_3_2((MulIn_data_sva_534[460]), FpMul_8U_23U_else_5_mux_52_mx0w1,
          FpMul_8U_23U_mux_220_itm, {and_1126_rgt , and_1129_rgt , and_1130_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_30_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1457_nl))
        ) begin
      FpMul_8U_23U_lor_30_lpi_1_dfm_6 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_19_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_13_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1458_nl)) ) begin
      IsNaN_8U_23U_1_land_13_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_13_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_204_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_1135_rgt | and_1138_rgt | and_1139_rgt) & (~ (mux_1460_nl))
        ) begin
      FpMul_8U_23U_mux_204_itm_3 <= MUX1HOT_s_1_3_2((MulIn_data_sva_534[427]), FpMul_8U_23U_else_5_mux_48_mx0w1,
          FpMul_8U_23U_mux_204_itm, {and_1135_rgt , and_1138_rgt , and_1139_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_29_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1461_nl))
        ) begin
      FpMul_8U_23U_lor_29_lpi_1_dfm_6 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_20_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_12_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1462_nl)) ) begin
      IsNaN_8U_23U_1_land_12_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_12_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_188_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_1144_rgt | and_1147_rgt | and_1148_rgt) & (~ (mux_1464_nl))
        ) begin
      FpMul_8U_23U_mux_188_itm_3 <= MUX1HOT_s_1_3_2((MulIn_data_sva_534[394]), FpMul_8U_23U_else_5_mux_44_mx0w1,
          FpMul_8U_23U_mux_188_itm, {and_1144_rgt , and_1147_rgt , and_1148_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_28_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1465_nl))
        ) begin
      FpMul_8U_23U_lor_28_lpi_1_dfm_6 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_21_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_11_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1466_nl)) ) begin
      IsNaN_8U_23U_1_land_11_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_11_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_172_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_1153_rgt | and_1156_rgt | and_1157_rgt) & (~ (mux_1468_nl))
        ) begin
      FpMul_8U_23U_mux_172_itm_3 <= MUX1HOT_s_1_3_2((MulIn_data_sva_534[361]), FpMul_8U_23U_else_5_mux_40_mx0w1,
          FpMul_8U_23U_mux_172_itm, {and_1153_rgt , and_1156_rgt , and_1157_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_27_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1469_nl))
        ) begin
      FpMul_8U_23U_lor_27_lpi_1_dfm_6 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_22_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_10_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1470_nl)) ) begin
      IsNaN_8U_23U_1_land_10_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_10_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_156_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_1162_rgt | and_1165_rgt | and_1166_rgt) & (~ (mux_1472_nl))
        ) begin
      FpMul_8U_23U_mux_156_itm_3 <= MUX1HOT_s_1_3_2((MulIn_data_sva_534[328]), FpMul_8U_23U_else_5_mux_36_mx0w1,
          FpMul_8U_23U_mux_156_itm, {and_1162_rgt , and_1165_rgt , and_1166_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_26_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1473_nl))
        ) begin
      FpMul_8U_23U_lor_26_lpi_1_dfm_6 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_23_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_9_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1474_nl)) ) begin
      IsNaN_8U_23U_1_land_9_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_9_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_140_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_1171_rgt | and_1174_rgt | and_1175_rgt) & (~ (mux_1476_nl))
        ) begin
      FpMul_8U_23U_mux_140_itm_3 <= MUX1HOT_s_1_3_2((MulIn_data_sva_534[295]), FpMul_8U_23U_else_5_mux_32_mx0w1,
          FpMul_8U_23U_mux_140_itm, {and_1171_rgt , and_1174_rgt , and_1175_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_25_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1477_nl))
        ) begin
      FpMul_8U_23U_lor_25_lpi_1_dfm_6 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_24_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_8_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1478_nl)) ) begin
      IsNaN_8U_23U_1_land_8_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_8_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_124_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_1180_rgt | and_1183_rgt | and_1184_rgt) & (~ (mux_1480_nl))
        ) begin
      FpMul_8U_23U_mux_124_itm_3 <= MUX1HOT_s_1_3_2((MulIn_data_sva_534[262]), FpMul_8U_23U_else_5_mux_28_mx0w1,
          FpMul_8U_23U_mux_124_itm, {and_1180_rgt , and_1183_rgt , and_1184_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_24_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1481_nl))
        ) begin
      FpMul_8U_23U_lor_24_lpi_1_dfm_6 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_25_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_7_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1482_nl)) ) begin
      IsNaN_8U_23U_1_land_7_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_7_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_108_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_1189_rgt | and_1192_rgt | and_1193_rgt) & (~ (mux_1484_nl))
        ) begin
      FpMul_8U_23U_mux_108_itm_3 <= MUX1HOT_s_1_3_2((MulIn_data_sva_534[229]), FpMul_8U_23U_else_5_mux_24_mx0w1,
          FpMul_8U_23U_mux_108_itm, {and_1189_rgt , and_1192_rgt , and_1193_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_23_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1485_nl))
        ) begin
      FpMul_8U_23U_lor_23_lpi_1_dfm_6 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_26_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_6_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1486_nl)) ) begin
      IsNaN_8U_23U_1_land_6_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_6_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_92_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_1198_rgt | and_1201_rgt | and_1202_rgt) & (~ (mux_1488_nl))
        ) begin
      FpMul_8U_23U_mux_92_itm_3 <= MUX1HOT_s_1_3_2((MulIn_data_sva_534[196]), FpMul_8U_23U_else_5_mux_20_mx0w1,
          FpMul_8U_23U_mux_92_itm, {and_1198_rgt , and_1201_rgt , and_1202_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_22_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1489_nl))
        ) begin
      FpMul_8U_23U_lor_22_lpi_1_dfm_6 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_27_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_5_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1490_nl)) ) begin
      IsNaN_8U_23U_1_land_5_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_5_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_76_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_1207_rgt | and_1210_rgt | and_1211_rgt) & (~ (mux_1492_nl))
        ) begin
      FpMul_8U_23U_mux_76_itm_3 <= MUX1HOT_s_1_3_2((MulIn_data_sva_534[163]), FpMul_8U_23U_else_5_mux_16_mx0w1,
          FpMul_8U_23U_mux_76_itm, {and_1207_rgt , and_1210_rgt , and_1211_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_21_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1493_nl))
        ) begin
      FpMul_8U_23U_lor_21_lpi_1_dfm_6 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_28_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_4_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1494_nl)) ) begin
      IsNaN_8U_23U_1_land_4_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_4_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_60_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_1216_rgt | and_1219_rgt | and_1220_rgt) & (~ (mux_1496_nl))
        ) begin
      FpMul_8U_23U_mux_60_itm_3 <= MUX1HOT_s_1_3_2((MulIn_data_sva_534[130]), FpMul_8U_23U_else_5_mux_12_mx0w1,
          FpMul_8U_23U_mux_60_itm, {and_1216_rgt , and_1219_rgt , and_1220_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_20_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1497_nl))
        ) begin
      FpMul_8U_23U_lor_20_lpi_1_dfm_6 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_29_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1498_nl)) ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_44_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_1225_rgt | and_1228_rgt | and_1229_rgt) & (~ (mux_1500_nl))
        ) begin
      FpMul_8U_23U_mux_44_itm_3 <= MUX1HOT_s_1_3_2((MulIn_data_sva_534[97]), FpMul_8U_23U_else_5_mux_8_mx0w1,
          FpMul_8U_23U_mux_44_itm, {and_1225_rgt , and_1228_rgt , and_1229_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_19_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1501_nl))
        ) begin
      FpMul_8U_23U_lor_19_lpi_1_dfm_6 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_30_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1502_nl)) ) begin
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_28_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_1234_rgt | and_1237_rgt | and_1238_rgt) & (~ (mux_1504_nl))
        ) begin
      FpMul_8U_23U_mux_28_itm_3 <= MUX1HOT_s_1_3_2((MulIn_data_sva_534[64]), FpMul_8U_23U_else_5_mux_4_mx0w1,
          FpMul_8U_23U_mux_28_itm, {and_1234_rgt , and_1237_rgt , and_1238_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_18_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_oelse_FpMul_8U_23U_oelse_or_37_cse & (~ (mux_1505_nl))
        ) begin
      FpMul_8U_23U_lor_18_lpi_1_dfm_6 <= FpMul_8U_23U_oelse_1_FpMul_8U_23U_oelse_1_mux_31_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1506_nl)) ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_12_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_1243_rgt | and_1246_rgt | and_1247_rgt) & (~ (mux_1508_nl))
        ) begin
      FpMul_8U_23U_mux_12_itm_3 <= MUX1HOT_s_1_3_2((MulIn_data_sva_534[31]), FpMul_8U_23U_else_5_mux_mx0w1,
          FpMul_8U_23U_mux_12_itm, {and_1243_rgt , and_1246_rgt , and_1247_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_15_sva_9 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1510_nl)) ) begin
      MulOut_data_15_sva_9 <= MulOut_data_15_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_14_sva_9 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1513_nl)) ) begin
      MulOut_data_14_sva_9 <= MulOut_data_14_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_13_sva_9 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1516_nl)) ) begin
      MulOut_data_13_sva_9 <= MulOut_data_13_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_12_sva_9 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1519_nl)) ) begin
      MulOut_data_12_sva_9 <= MulOut_data_12_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_11_sva_9 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1522_nl)) ) begin
      MulOut_data_11_sva_9 <= MulOut_data_11_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_10_sva_9 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1525_nl)) ) begin
      MulOut_data_10_sva_9 <= MulOut_data_10_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_9_sva_9 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1527_nl)) ) begin
      MulOut_data_9_sva_9 <= MulOut_data_9_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_8_sva_9 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1529_nl)) ) begin
      MulOut_data_8_sva_9 <= MulOut_data_8_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_7_sva_9 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1531_nl)) ) begin
      MulOut_data_7_sva_9 <= MulOut_data_7_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_6_sva_9 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1533_nl)) ) begin
      MulOut_data_6_sva_9 <= MulOut_data_6_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_5_sva_9 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1535_nl)) ) begin
      MulOut_data_5_sva_9 <= MulOut_data_5_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_4_sva_9 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1537_nl)) ) begin
      MulOut_data_4_sva_9 <= MulOut_data_4_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_3_sva_9 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1539_nl)) ) begin
      MulOut_data_3_sva_9 <= MulOut_data_3_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_2_sva_9 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1541_nl)) ) begin
      MulOut_data_2_sva_9 <= MulOut_data_2_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_1_sva_9 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1544_nl)) ) begin
      MulOut_data_1_sva_9 <= MulOut_data_1_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_0_sva_9 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ (mux_1547_nl)) ) begin
      MulOut_data_0_sva_9 <= MulOut_data_0_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_187_itm) ) begin
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_7 <= IsNaN_8U_23U_land_1_lpi_1_dfm_st_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_202_itm) ) begin
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_7 <= IsNaN_8U_23U_land_2_lpi_1_dfm_st_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_216_itm) ) begin
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_7 <= IsNaN_8U_23U_land_3_lpi_1_dfm_st_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_4_lpi_1_dfm_st_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_230_itm) ) begin
      IsNaN_8U_23U_land_4_lpi_1_dfm_st_7 <= IsNaN_8U_23U_land_4_lpi_1_dfm_st_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_5_lpi_1_dfm_st_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_245_itm) ) begin
      IsNaN_8U_23U_land_5_lpi_1_dfm_st_7 <= IsNaN_8U_23U_land_5_lpi_1_dfm_st_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_6_lpi_1_dfm_st_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_259_itm) ) begin
      IsNaN_8U_23U_land_6_lpi_1_dfm_st_7 <= IsNaN_8U_23U_land_6_lpi_1_dfm_st_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_7_lpi_1_dfm_st_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_273_itm) ) begin
      IsNaN_8U_23U_land_7_lpi_1_dfm_st_7 <= IsNaN_8U_23U_land_7_lpi_1_dfm_st_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_8_lpi_1_dfm_st_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_288_itm) ) begin
      IsNaN_8U_23U_land_8_lpi_1_dfm_st_7 <= IsNaN_8U_23U_land_8_lpi_1_dfm_st_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_9_lpi_1_dfm_st_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_303_itm) ) begin
      IsNaN_8U_23U_land_9_lpi_1_dfm_st_7 <= IsNaN_8U_23U_land_9_lpi_1_dfm_st_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_10_lpi_1_dfm_st_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_318_itm) ) begin
      IsNaN_8U_23U_land_10_lpi_1_dfm_st_7 <= IsNaN_8U_23U_land_10_lpi_1_dfm_st_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_11_lpi_1_dfm_st_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_332_itm) ) begin
      IsNaN_8U_23U_land_11_lpi_1_dfm_st_7 <= IsNaN_8U_23U_land_11_lpi_1_dfm_st_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_12_lpi_1_dfm_st_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_346_itm) ) begin
      IsNaN_8U_23U_land_12_lpi_1_dfm_st_7 <= IsNaN_8U_23U_land_12_lpi_1_dfm_st_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_13_lpi_1_dfm_st_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_360_itm) ) begin
      IsNaN_8U_23U_land_13_lpi_1_dfm_st_7 <= IsNaN_8U_23U_land_13_lpi_1_dfm_st_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_14_lpi_1_dfm_st_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_374_itm) ) begin
      IsNaN_8U_23U_land_14_lpi_1_dfm_st_7 <= IsNaN_8U_23U_land_14_lpi_1_dfm_st_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_15_lpi_1_dfm_st_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_388_itm) ) begin
      IsNaN_8U_23U_land_15_lpi_1_dfm_st_7 <= IsNaN_8U_23U_land_15_lpi_1_dfm_st_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_st_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_403_itm) ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_st_7 <= IsNaN_8U_23U_land_lpi_1_dfm_st_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_1_sva <= 48'b0;
    end
    else if ( core_wen & (~(or_tmp_608 | mul_loop_mul_if_land_1_lpi_1_dfm_st_7 |
        FpMul_8U_23U_lor_18_lpi_1_dfm_st_3 | or_dcpl_87)) & mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        ) begin
      FpMul_8U_23U_p_mant_p1_1_sva <= mul_loop_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= 1'b0;
    end
    else if ( core_wen & (((~ mul_loop_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1) &
        or_309_cse & (~ reg_FpMul_8U_23U_lor_3_lpi_1_dfm_4_cse) & (cfg_precision==2'b10))
        | and_1252_rgt) & (~ mux_187_itm) ) begin
      mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= MUX_s_1_2_2(mul_loop_mul_1_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_1252_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_2_sva <= 48'b0;
    end
    else if ( core_wen & (~(or_tmp_608 | mul_loop_mul_if_land_2_lpi_1_dfm_st_7 |
        FpMul_8U_23U_lor_19_lpi_1_dfm_st_3 | or_dcpl_87)) & mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        ) begin
      FpMul_8U_23U_p_mant_p1_2_sva <= mul_loop_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= 1'b0;
    end
    else if ( core_wen & (((~ mul_loop_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1) &
        or_309_cse & (~ reg_FpMul_8U_23U_lor_4_lpi_1_dfm_4_cse) & (cfg_precision==2'b10))
        | and_1257_rgt) & (~ mux_202_itm) ) begin
      mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= MUX_s_1_2_2(mul_loop_mul_2_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_1257_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_3_sva <= 48'b0;
    end
    else if ( core_wen & (~(or_tmp_608 | mul_loop_mul_if_land_3_lpi_1_dfm_st_7 |
        FpMul_8U_23U_lor_20_lpi_1_dfm_st_3 | or_dcpl_87)) & mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        ) begin
      FpMul_8U_23U_p_mant_p1_3_sva <= mul_loop_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= 1'b0;
    end
    else if ( core_wen & (((~ mul_loop_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1) &
        or_309_cse & (~ reg_FpMul_8U_23U_lor_5_lpi_1_dfm_4_cse) & (cfg_precision==2'b10))
        | and_1262_rgt) & (~ mux_216_itm) ) begin
      mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= MUX_s_1_2_2(mul_loop_mul_3_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_1262_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_4_sva <= 48'b0;
    end
    else if ( core_wen & (~(or_dcpl_95 | mul_loop_mul_if_land_4_lpi_1_dfm_st_7 |
        FpMul_8U_23U_lor_21_lpi_1_dfm_st_3 | or_90_cse)) & mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        ) begin
      FpMul_8U_23U_p_mant_p1_4_sva <= mul_loop_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= 1'b0;
    end
    else if ( core_wen & (((~ mul_loop_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1) &
        or_309_cse & (~ reg_FpMul_8U_23U_lor_6_lpi_1_dfm_4_cse) & (cfg_precision==2'b10))
        | and_1267_rgt) & (~ mux_230_itm) ) begin
      mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= MUX_s_1_2_2(mul_loop_mul_4_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_1267_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_5_sva <= 48'b0;
    end
    else if ( core_wen & (~(or_tmp_608 | mul_loop_mul_if_land_5_lpi_1_dfm_st_7 |
        FpMul_8U_23U_lor_22_lpi_1_dfm_st_3 | or_dcpl_87)) & mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        ) begin
      FpMul_8U_23U_p_mant_p1_5_sva <= mul_loop_mul_5_FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= 1'b0;
    end
    else if ( core_wen & (((~ mul_loop_mul_5_FpMul_8U_23U_oelse_1_acc_itm_9_1) &
        or_309_cse & (~ reg_FpMul_8U_23U_lor_7_lpi_1_dfm_4_cse) & (cfg_precision==2'b10))
        | and_1272_rgt) & (~ mux_245_itm) ) begin
      mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= MUX_s_1_2_2(mul_loop_mul_5_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_1272_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_6_sva <= 48'b0;
    end
    else if ( core_wen & (~(or_tmp_608 | mul_loop_mul_if_land_6_lpi_1_dfm_st_7 |
        FpMul_8U_23U_lor_23_lpi_1_dfm_st_3 | or_dcpl_87)) & mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        ) begin
      FpMul_8U_23U_p_mant_p1_6_sva <= mul_loop_mul_6_FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= 1'b0;
    end
    else if ( core_wen & (((~ mul_loop_mul_6_FpMul_8U_23U_oelse_1_acc_itm_9_1) &
        or_309_cse & (~ reg_FpMul_8U_23U_lor_8_lpi_1_dfm_4_cse) & (cfg_precision==2'b10))
        | and_1277_rgt) & (~ mux_259_itm) ) begin
      mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= MUX_s_1_2_2(mul_loop_mul_6_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_1277_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_7_sva <= 48'b0;
    end
    else if ( core_wen & (~(or_tmp_608 | mul_loop_mul_if_land_7_lpi_1_dfm_st_7 |
        FpMul_8U_23U_lor_24_lpi_1_dfm_st_3 | or_dcpl_87)) & mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        ) begin
      FpMul_8U_23U_p_mant_p1_7_sva <= mul_loop_mul_7_FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= 1'b0;
    end
    else if ( core_wen & (((~ mul_loop_mul_7_FpMul_8U_23U_oelse_1_acc_itm_9_1) &
        or_309_cse & (~ reg_FpMul_8U_23U_lor_9_lpi_1_dfm_4_cse) & (cfg_precision==2'b10))
        | and_1282_rgt) & (~ mux_273_itm) ) begin
      mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= MUX_s_1_2_2(mul_loop_mul_7_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_1282_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_8_sva <= 48'b0;
    end
    else if ( core_wen & (~(or_tmp_608 | mul_loop_mul_if_land_8_lpi_1_dfm_st_7 |
        FpMul_8U_23U_lor_25_lpi_1_dfm_st_3 | or_dcpl_87)) & mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        ) begin
      FpMul_8U_23U_p_mant_p1_8_sva <= mul_loop_mul_8_FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= 1'b0;
    end
    else if ( core_wen & (((~ mul_loop_mul_8_FpMul_8U_23U_oelse_1_acc_itm_9_1) &
        or_309_cse & (~ reg_FpMul_8U_23U_lor_10_lpi_1_dfm_4_cse) & (cfg_precision==2'b10))
        | and_1287_rgt) & (~ mux_288_itm) ) begin
      mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= MUX_s_1_2_2(mul_loop_mul_8_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_1287_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_9_sva <= 48'b0;
    end
    else if ( core_wen & (~(or_tmp_608 | mul_loop_mul_if_land_9_lpi_1_dfm_st_7 |
        FpMul_8U_23U_lor_26_lpi_1_dfm_st_3 | or_dcpl_87)) & mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        ) begin
      FpMul_8U_23U_p_mant_p1_9_sva <= mul_loop_mul_9_FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= 1'b0;
    end
    else if ( core_wen & (((~ mul_loop_mul_9_FpMul_8U_23U_oelse_1_acc_itm_9_1) &
        or_309_cse & (~ reg_FpMul_8U_23U_lor_11_lpi_1_dfm_4_cse) & (cfg_precision==2'b10))
        | and_1292_rgt) & (~ mux_303_itm) ) begin
      mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= MUX_s_1_2_2(mul_loop_mul_9_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_1292_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_10_sva <= 48'b0;
    end
    else if ( core_wen & (~(or_tmp_608 | mul_loop_mul_if_land_10_lpi_1_dfm_st_7 |
        FpMul_8U_23U_lor_27_lpi_1_dfm_st_3 | or_dcpl_87)) & mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        ) begin
      FpMul_8U_23U_p_mant_p1_10_sva <= mul_loop_mul_10_FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= 1'b0;
    end
    else if ( core_wen & (((~ mul_loop_mul_10_FpMul_8U_23U_oelse_1_acc_itm_9_1) &
        or_309_cse & (~ reg_FpMul_8U_23U_lor_12_lpi_1_dfm_4_cse) & (cfg_precision==2'b10))
        | and_1297_rgt) & (~ mux_318_itm) ) begin
      mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= MUX_s_1_2_2(mul_loop_mul_10_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_1297_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_11_sva <= 48'b0;
    end
    else if ( core_wen & (~(or_dcpl_95 | mul_loop_mul_if_land_11_lpi_1_dfm_st_7 |
        FpMul_8U_23U_lor_28_lpi_1_dfm_st_3 | or_90_cse)) & mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        ) begin
      FpMul_8U_23U_p_mant_p1_11_sva <= mul_loop_mul_11_FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= 1'b0;
    end
    else if ( core_wen & (((~ mul_loop_mul_11_FpMul_8U_23U_oelse_1_acc_itm_9_1) &
        or_309_cse & (~ reg_FpMul_8U_23U_lor_13_lpi_1_dfm_4_cse) & (cfg_precision==2'b10))
        | and_1302_rgt) & (~ mux_332_itm) ) begin
      mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= MUX_s_1_2_2(mul_loop_mul_11_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_1302_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_12_sva <= 48'b0;
    end
    else if ( core_wen & (~(or_dcpl_95 | mul_loop_mul_if_land_12_lpi_1_dfm_st_7 |
        FpMul_8U_23U_lor_29_lpi_1_dfm_st_3 | or_90_cse)) & mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        ) begin
      FpMul_8U_23U_p_mant_p1_12_sva <= mul_loop_mul_12_FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= 1'b0;
    end
    else if ( core_wen & (((~ mul_loop_mul_12_FpMul_8U_23U_oelse_1_acc_itm_9_1) &
        or_309_cse & (~ reg_FpMul_8U_23U_lor_14_lpi_1_dfm_4_cse) & (cfg_precision==2'b10))
        | and_1307_rgt) & (~ mux_346_itm) ) begin
      mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= MUX_s_1_2_2(mul_loop_mul_12_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_1307_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_13_sva <= 48'b0;
    end
    else if ( core_wen & (~(or_dcpl_95 | mul_loop_mul_if_land_13_lpi_1_dfm_st_7 |
        FpMul_8U_23U_lor_30_lpi_1_dfm_st_3 | or_90_cse)) & mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        ) begin
      FpMul_8U_23U_p_mant_p1_13_sva <= mul_loop_mul_13_FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= 1'b0;
    end
    else if ( core_wen & (((~ mul_loop_mul_13_FpMul_8U_23U_oelse_1_acc_itm_9_1) &
        or_309_cse & (~ reg_FpMul_8U_23U_lor_15_lpi_1_dfm_4_cse) & (cfg_precision==2'b10))
        | and_1312_rgt) & (~ mux_360_itm) ) begin
      mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= MUX_s_1_2_2(mul_loop_mul_13_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_1312_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_14_sva <= 48'b0;
    end
    else if ( core_wen & (~(or_tmp_608 | mul_loop_mul_if_land_14_lpi_1_dfm_st_7 |
        FpMul_8U_23U_lor_31_lpi_1_dfm_st_3 | or_dcpl_87)) & mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        ) begin
      FpMul_8U_23U_p_mant_p1_14_sva <= mul_loop_mul_14_FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= 1'b0;
    end
    else if ( core_wen & (((~ mul_loop_mul_14_FpMul_8U_23U_oelse_1_acc_itm_9_1) &
        or_309_cse & (~ reg_FpMul_8U_23U_lor_16_lpi_1_dfm_4_cse) & (cfg_precision==2'b10))
        | and_1317_rgt) & (~ mux_374_itm) ) begin
      mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= MUX_s_1_2_2(mul_loop_mul_14_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_1317_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_15_sva <= 48'b0;
    end
    else if ( core_wen & (~(or_tmp_608 | mul_loop_mul_if_land_15_lpi_1_dfm_st_7 |
        FpMul_8U_23U_lor_32_lpi_1_dfm_st_3 | or_dcpl_87)) & mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        ) begin
      FpMul_8U_23U_p_mant_p1_15_sva <= mul_loop_mul_15_FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= 1'b0;
    end
    else if ( core_wen & (((~ mul_loop_mul_15_FpMul_8U_23U_oelse_1_acc_itm_9_1) &
        or_309_cse & (~ reg_FpMul_8U_23U_lor_17_lpi_1_dfm_4_cse) & (cfg_precision==2'b10))
        | and_1322_rgt) & (~ mux_388_itm) ) begin
      mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= MUX_s_1_2_2(mul_loop_mul_15_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_1322_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_sva <= 48'b0;
    end
    else if ( core_wen & (~(or_tmp_608 | mul_loop_mul_if_land_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3
        | or_dcpl_87)) & mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        ) begin
      FpMul_8U_23U_p_mant_p1_sva <= mul_loop_mul_16_FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= 1'b0;
    end
    else if ( core_wen & (((~ mul_loop_mul_16_FpMul_8U_23U_oelse_1_acc_itm_9_1) &
        or_309_cse & (~ reg_FpMul_8U_23U_lor_lpi_1_dfm_4_cse) & (cfg_precision==2'b10))
        | and_1327_rgt) & (~ mux_403_itm) ) begin
      mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
          <= MUX_s_1_2_2(mul_loop_mul_16_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_1327_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_1_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( FpMul_8U_23U_else_2_if_and_cse & (~ or_dcpl_373) & (~ (mux_1445_nl))
        ) begin
      IsZero_8U_23U_1_land_1_lpi_1_dfm <= IsZero_8U_23U_1_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_tmp_204 | mul_loop_mul_if_land_1_lpi_1_dfm_st_6 |
        mul_loop_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1 | and_dcpl_50 | reg_FpMul_8U_23U_lor_3_lpi_1_dfm_4_cse
        | or_90_cse)) ) begin
      mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= mul_loop_mul_1_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_12_itm <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_770 & (~ mul_loop_mul_if_land_1_lpi_1_dfm_st_6)
        & IsNaN_8U_23U_land_1_lpi_1_dfm_9 & and_dcpl_85) | FpMul_8U_23U_mux_12_itm_mx0c1)
        ) begin
      FpMul_8U_23U_mux_12_itm <= MUX_s_1_2_2((MulIn_data_sva_534[31]), FpMul_8U_23U_else_5_mux_mx0w1,
          FpMul_8U_23U_mux_12_itm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_tmp_204 | mul_loop_mul_if_land_2_lpi_1_dfm_st_6 |
        mul_loop_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1 | and_dcpl_50 | reg_FpMul_8U_23U_lor_4_lpi_1_dfm_4_cse
        | or_90_cse)) ) begin
      mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= mul_loop_mul_2_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_28_itm <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_770 & (~ mul_loop_mul_if_land_2_lpi_1_dfm_st_6)
        & IsNaN_8U_23U_land_2_lpi_1_dfm_9 & and_dcpl_85) | FpMul_8U_23U_mux_28_itm_mx0c1)
        ) begin
      FpMul_8U_23U_mux_28_itm <= MUX_s_1_2_2((MulIn_data_sva_534[64]), FpMul_8U_23U_else_5_mux_4_mx0w1,
          FpMul_8U_23U_mux_28_itm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_tmp_204 | mul_loop_mul_if_land_3_lpi_1_dfm_st_6 |
        mul_loop_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1 | and_dcpl_50 | reg_FpMul_8U_23U_lor_5_lpi_1_dfm_4_cse
        | or_90_cse)) ) begin
      mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= mul_loop_mul_3_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_44_itm <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_770 & (~ mul_loop_mul_if_land_3_lpi_1_dfm_st_6)
        & IsNaN_8U_23U_land_3_lpi_1_dfm_9 & and_dcpl_85) | FpMul_8U_23U_mux_44_itm_mx0c1)
        ) begin
      FpMul_8U_23U_mux_44_itm <= MUX_s_1_2_2((MulIn_data_sva_534[97]), FpMul_8U_23U_else_5_mux_8_mx0w1,
          FpMul_8U_23U_mux_44_itm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_tmp_204 | mul_loop_mul_if_land_4_lpi_1_dfm_st_6 |
        mul_loop_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1 | and_dcpl_50 | reg_FpMul_8U_23U_lor_6_lpi_1_dfm_4_cse
        | or_90_cse)) ) begin
      mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= mul_loop_mul_4_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_60_itm <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_770 & (~ mul_loop_mul_if_land_4_lpi_1_dfm_st_6)
        & IsNaN_8U_23U_land_4_lpi_1_dfm_9 & and_dcpl_85) | FpMul_8U_23U_mux_60_itm_mx0c1)
        ) begin
      FpMul_8U_23U_mux_60_itm <= MUX_s_1_2_2((MulIn_data_sva_534[130]), FpMul_8U_23U_else_5_mux_12_mx0w1,
          FpMul_8U_23U_mux_60_itm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_tmp_204 | mul_loop_mul_if_land_5_lpi_1_dfm_st_6 |
        mul_loop_mul_5_FpMul_8U_23U_oelse_1_acc_itm_9_1 | and_dcpl_50 | reg_FpMul_8U_23U_lor_7_lpi_1_dfm_4_cse
        | or_90_cse)) ) begin
      mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= mul_loop_mul_5_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_76_itm <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_770 & (~ mul_loop_mul_if_land_5_lpi_1_dfm_st_6)
        & IsNaN_8U_23U_land_5_lpi_1_dfm_9 & and_dcpl_85) | FpMul_8U_23U_mux_76_itm_mx0c1)
        ) begin
      FpMul_8U_23U_mux_76_itm <= MUX_s_1_2_2((MulIn_data_sva_534[163]), FpMul_8U_23U_else_5_mux_16_mx0w1,
          FpMul_8U_23U_mux_76_itm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_tmp_204 | mul_loop_mul_if_land_6_lpi_1_dfm_st_6 |
        mul_loop_mul_6_FpMul_8U_23U_oelse_1_acc_itm_9_1 | and_dcpl_50 | reg_FpMul_8U_23U_lor_8_lpi_1_dfm_4_cse
        | or_90_cse)) ) begin
      mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= mul_loop_mul_6_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_92_itm <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_770 & (~ mul_loop_mul_if_land_6_lpi_1_dfm_st_6)
        & IsNaN_8U_23U_land_6_lpi_1_dfm_9 & and_dcpl_85) | FpMul_8U_23U_mux_92_itm_mx0c1)
        ) begin
      FpMul_8U_23U_mux_92_itm <= MUX_s_1_2_2((MulIn_data_sva_534[196]), FpMul_8U_23U_else_5_mux_20_mx0w1,
          FpMul_8U_23U_mux_92_itm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_tmp_204 | mul_loop_mul_if_land_7_lpi_1_dfm_st_6 |
        mul_loop_mul_7_FpMul_8U_23U_oelse_1_acc_itm_9_1 | and_dcpl_50 | reg_FpMul_8U_23U_lor_9_lpi_1_dfm_4_cse
        | or_90_cse)) ) begin
      mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= mul_loop_mul_7_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_108_itm <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_770 & (~ mul_loop_mul_if_land_7_lpi_1_dfm_st_6)
        & IsNaN_8U_23U_land_7_lpi_1_dfm_9 & and_dcpl_85) | FpMul_8U_23U_mux_108_itm_mx0c1)
        ) begin
      FpMul_8U_23U_mux_108_itm <= MUX_s_1_2_2((MulIn_data_sva_534[229]), FpMul_8U_23U_else_5_mux_24_mx0w1,
          FpMul_8U_23U_mux_108_itm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_tmp_204 | mul_loop_mul_if_land_8_lpi_1_dfm_st_6 |
        mul_loop_mul_8_FpMul_8U_23U_oelse_1_acc_itm_9_1 | and_dcpl_50 | reg_FpMul_8U_23U_lor_10_lpi_1_dfm_4_cse
        | or_90_cse)) ) begin
      mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= mul_loop_mul_8_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_124_itm <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_770 & (~ mul_loop_mul_if_land_8_lpi_1_dfm_st_6)
        & IsNaN_8U_23U_land_8_lpi_1_dfm_9 & and_dcpl_85) | FpMul_8U_23U_mux_124_itm_mx0c1)
        ) begin
      FpMul_8U_23U_mux_124_itm <= MUX_s_1_2_2((MulIn_data_sva_534[262]), FpMul_8U_23U_else_5_mux_28_mx0w1,
          FpMul_8U_23U_mux_124_itm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_tmp_204 | mul_loop_mul_if_land_9_lpi_1_dfm_st_6 |
        mul_loop_mul_9_FpMul_8U_23U_oelse_1_acc_itm_9_1 | and_dcpl_50 | reg_FpMul_8U_23U_lor_11_lpi_1_dfm_4_cse
        | or_90_cse)) ) begin
      mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= mul_loop_mul_9_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_140_itm <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_770 & (~ mul_loop_mul_if_land_9_lpi_1_dfm_st_6)
        & IsNaN_8U_23U_land_9_lpi_1_dfm_9 & and_dcpl_85) | FpMul_8U_23U_mux_140_itm_mx0c1)
        ) begin
      FpMul_8U_23U_mux_140_itm <= MUX_s_1_2_2((MulIn_data_sva_534[295]), FpMul_8U_23U_else_5_mux_32_mx0w1,
          FpMul_8U_23U_mux_140_itm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_tmp_204 | mul_loop_mul_if_land_10_lpi_1_dfm_st_6 |
        mul_loop_mul_10_FpMul_8U_23U_oelse_1_acc_itm_9_1 | and_dcpl_50 | reg_FpMul_8U_23U_lor_12_lpi_1_dfm_4_cse
        | or_90_cse)) ) begin
      mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= mul_loop_mul_10_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_156_itm <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_770 & (~ mul_loop_mul_if_land_10_lpi_1_dfm_st_6)
        & IsNaN_8U_23U_land_10_lpi_1_dfm_9 & and_dcpl_85) | FpMul_8U_23U_mux_156_itm_mx0c1)
        ) begin
      FpMul_8U_23U_mux_156_itm <= MUX_s_1_2_2((MulIn_data_sva_534[328]), FpMul_8U_23U_else_5_mux_36_mx0w1,
          FpMul_8U_23U_mux_156_itm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_tmp_204 | mul_loop_mul_if_land_11_lpi_1_dfm_st_6 |
        mul_loop_mul_11_FpMul_8U_23U_oelse_1_acc_itm_9_1 | and_dcpl_50 | reg_FpMul_8U_23U_lor_13_lpi_1_dfm_4_cse
        | or_90_cse)) ) begin
      mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= mul_loop_mul_11_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_172_itm <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_770 & (~ mul_loop_mul_if_land_11_lpi_1_dfm_st_6)
        & IsNaN_8U_23U_land_11_lpi_1_dfm_9 & and_dcpl_85) | FpMul_8U_23U_mux_172_itm_mx0c1)
        ) begin
      FpMul_8U_23U_mux_172_itm <= MUX_s_1_2_2((MulIn_data_sva_534[361]), FpMul_8U_23U_else_5_mux_40_mx0w1,
          FpMul_8U_23U_mux_172_itm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_tmp_204 | mul_loop_mul_if_land_12_lpi_1_dfm_st_6 |
        mul_loop_mul_12_FpMul_8U_23U_oelse_1_acc_itm_9_1 | and_dcpl_50 | reg_FpMul_8U_23U_lor_14_lpi_1_dfm_4_cse
        | or_90_cse)) ) begin
      mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= mul_loop_mul_12_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_188_itm <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_770 & (~ mul_loop_mul_if_land_12_lpi_1_dfm_st_6)
        & IsNaN_8U_23U_land_12_lpi_1_dfm_9 & and_dcpl_85) | FpMul_8U_23U_mux_188_itm_mx0c1)
        ) begin
      FpMul_8U_23U_mux_188_itm <= MUX_s_1_2_2((MulIn_data_sva_534[394]), FpMul_8U_23U_else_5_mux_44_mx0w1,
          FpMul_8U_23U_mux_188_itm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_tmp_204 | mul_loop_mul_if_land_13_lpi_1_dfm_st_6 |
        mul_loop_mul_13_FpMul_8U_23U_oelse_1_acc_itm_9_1 | and_dcpl_50 | reg_FpMul_8U_23U_lor_15_lpi_1_dfm_4_cse
        | or_90_cse)) ) begin
      mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= mul_loop_mul_13_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_204_itm <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_770 & (~ mul_loop_mul_if_land_13_lpi_1_dfm_st_6)
        & IsNaN_8U_23U_land_13_lpi_1_dfm_9 & and_dcpl_85) | FpMul_8U_23U_mux_204_itm_mx0c1)
        ) begin
      FpMul_8U_23U_mux_204_itm <= MUX_s_1_2_2((MulIn_data_sva_534[427]), FpMul_8U_23U_else_5_mux_48_mx0w1,
          FpMul_8U_23U_mux_204_itm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_tmp_204 | mul_loop_mul_if_land_14_lpi_1_dfm_st_6 |
        mul_loop_mul_14_FpMul_8U_23U_oelse_1_acc_itm_9_1 | and_dcpl_50 | reg_FpMul_8U_23U_lor_16_lpi_1_dfm_4_cse
        | or_90_cse)) ) begin
      mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= mul_loop_mul_14_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_220_itm <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_770 & (~ mul_loop_mul_if_land_14_lpi_1_dfm_st_6)
        & IsNaN_8U_23U_land_14_lpi_1_dfm_9 & and_dcpl_85) | FpMul_8U_23U_mux_220_itm_mx0c1)
        ) begin
      FpMul_8U_23U_mux_220_itm <= MUX_s_1_2_2((MulIn_data_sva_534[460]), FpMul_8U_23U_else_5_mux_52_mx0w1,
          FpMul_8U_23U_mux_220_itm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_tmp_204 | mul_loop_mul_if_land_15_lpi_1_dfm_st_6 |
        mul_loop_mul_15_FpMul_8U_23U_oelse_1_acc_itm_9_1 | and_dcpl_50 | reg_FpMul_8U_23U_lor_17_lpi_1_dfm_4_cse
        | or_90_cse)) ) begin
      mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= mul_loop_mul_15_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_236_itm <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_770 & (~ mul_loop_mul_if_land_15_lpi_1_dfm_st_6)
        & IsNaN_8U_23U_land_15_lpi_1_dfm_9 & and_dcpl_85) | FpMul_8U_23U_mux_236_itm_mx0c1)
        ) begin
      FpMul_8U_23U_mux_236_itm <= MUX_s_1_2_2((MulIn_data_sva_534[493]), FpMul_8U_23U_else_5_mux_56_mx0w1,
          FpMul_8U_23U_mux_236_itm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_tmp_204 | mul_loop_mul_if_land_lpi_1_dfm_st_6 | mul_loop_mul_16_FpMul_8U_23U_oelse_1_acc_itm_9_1
        | and_dcpl_50 | reg_FpMul_8U_23U_lor_lpi_1_dfm_4_cse | or_90_cse)) ) begin
      mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs
          <= mul_loop_mul_16_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_252_itm <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_770 & (~ mul_loop_mul_if_land_lpi_1_dfm_st_6)
        & IsNaN_8U_23U_land_lpi_1_dfm_9 & and_dcpl_85) | FpMul_8U_23U_mux_252_itm_mx0c1)
        ) begin
      FpMul_8U_23U_mux_252_itm <= MUX_s_1_2_2((MulIn_data_sva_534[526]), FpMul_8U_23U_else_5_mux_60_mx0w1,
          FpMul_8U_23U_mux_252_itm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1548_nl) ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 <= ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_9_0_mx1!=10'b0000000000))
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_3_2_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_1_lpi_1_dfm_3_1_0_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w0==4'b1111);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1549_nl) ) begin
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 <= ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_9_0_mx1!=10'b0000000000))
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_3_2_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_2_lpi_1_dfm_3_1_0_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w0==4'b1111);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1550_nl) ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 <= ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_9_0_mx1!=10'b0000000000))
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_3_2_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_3_lpi_1_dfm_3_1_0_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w0==4'b1111);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_4_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1551_nl) ) begin
      IsNaN_8U_23U_1_land_4_lpi_1_dfm_7 <= ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_9_0_mx1!=10'b0000000000))
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_3_2_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_4_lpi_1_dfm_3_1_0_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_4_lpi_1_dfm_3_mx0w0==4'b1111);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_5_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1552_nl) ) begin
      IsNaN_8U_23U_1_land_5_lpi_1_dfm_7 <= ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_9_0_mx1!=10'b0000000000))
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_3_2_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_5_lpi_1_dfm_3_1_0_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_5_lpi_1_dfm_3_mx0w0==4'b1111);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_6_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1553_nl) ) begin
      IsNaN_8U_23U_1_land_6_lpi_1_dfm_7 <= ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_9_0_mx1!=10'b0000000000))
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_3_2_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_6_lpi_1_dfm_3_1_0_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_6_lpi_1_dfm_3_mx0w0==4'b1111);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_7_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1554_nl) ) begin
      IsNaN_8U_23U_1_land_7_lpi_1_dfm_7 <= ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_9_0_mx1!=10'b0000000000))
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_3_2_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_7_lpi_1_dfm_3_1_0_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_7_lpi_1_dfm_3_mx0w0==4'b1111);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_8_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1555_nl) ) begin
      IsNaN_8U_23U_1_land_8_lpi_1_dfm_7 <= ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_9_0_mx1!=10'b0000000000))
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_3_2_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_8_lpi_1_dfm_3_1_0_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_8_lpi_1_dfm_3_mx0w0==4'b1111);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_9_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1556_nl) ) begin
      IsNaN_8U_23U_1_land_9_lpi_1_dfm_7 <= ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_9_0_mx1!=10'b0000000000))
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_3_2_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_9_lpi_1_dfm_3_1_0_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_9_lpi_1_dfm_3_mx0w0==4'b1111);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_10_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1557_nl) ) begin
      IsNaN_8U_23U_1_land_10_lpi_1_dfm_7 <= ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_9_0_mx1!=10'b0000000000))
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_3_2_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_10_lpi_1_dfm_3_1_0_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_10_lpi_1_dfm_3_mx0w0==4'b1111);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_11_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1558_nl) ) begin
      IsNaN_8U_23U_1_land_11_lpi_1_dfm_7 <= ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_9_0_mx1!=10'b0000000000))
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_3_2_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_11_lpi_1_dfm_3_1_0_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_11_lpi_1_dfm_3_mx0w0==4'b1111);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_12_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1559_nl) ) begin
      IsNaN_8U_23U_1_land_12_lpi_1_dfm_7 <= ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_9_0_mx1!=10'b0000000000))
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_3_2_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_12_lpi_1_dfm_3_1_0_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_12_lpi_1_dfm_3_mx0w0==4'b1111);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_13_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1560_nl) ) begin
      IsNaN_8U_23U_1_land_13_lpi_1_dfm_7 <= ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_9_0_mx1!=10'b0000000000))
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_3_2_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_13_lpi_1_dfm_3_1_0_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_13_lpi_1_dfm_3_mx0w0==4'b1111);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_14_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1561_nl) ) begin
      IsNaN_8U_23U_1_land_14_lpi_1_dfm_7 <= ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_9_0_mx1!=10'b0000000000))
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_3_2_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_14_lpi_1_dfm_3_1_0_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_14_lpi_1_dfm_3_mx0w0==4'b1111);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_15_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1562_nl) ) begin
      IsNaN_8U_23U_1_land_15_lpi_1_dfm_7 <= ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_9_0_mx1!=10'b0000000000))
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_3_2_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_15_lpi_1_dfm_3_1_0_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_15_lpi_1_dfm_3_mx0w0==4'b1111);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1563_nl) ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_7 <= ((FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_22_13_mx1!=10'b0000000000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_12_10_mx0w0!=3'b000)
          | (FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_9_0_mx1!=10'b0000000000))
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_3_2_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_7_4_lpi_1_dfm_3_1_0_mx0w0==2'b11)
          & (FpExpoWidthInc_5U_8U_23U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w0==4'b1111);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_1_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_65_mx0w1,
          and_dcpl_879);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_1_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_1_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_64_mx0w1,
          and_dcpl_879);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_3_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_2_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_68_mx0w1,
          and_dcpl_891);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_2_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_2_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_67_mx0w1,
          and_dcpl_891);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_6_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_3_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_71_mx0w1,
          and_dcpl_903);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_3_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_3_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_70_mx0w1,
          and_dcpl_903);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_9_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_4_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_74_mx0w1,
          and_dcpl_915);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_4_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_4_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_73_mx0w1,
          and_dcpl_915);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_12_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_5_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_77_mx0w1,
          and_dcpl_927);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_5_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_5_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_76_mx0w1,
          and_dcpl_927);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_15_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_6_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_80_mx0w1,
          and_dcpl_939);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_6_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_6_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_79_mx0w1,
          and_dcpl_939);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_18_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_7_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_83_mx0w1,
          and_dcpl_951);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_7_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_7_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_82_mx0w1,
          and_dcpl_951);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_21_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_8_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_86_mx0w1,
          and_dcpl_963);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_8_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_8_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_85_mx0w1,
          and_dcpl_963);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_24_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_9_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_89_mx0w1,
          and_dcpl_975);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_9_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_9_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_88_mx0w1,
          and_dcpl_975);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_27_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_10_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_92_mx0w1,
          and_dcpl_987);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_10_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_10_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_91_mx0w1,
          and_dcpl_987);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_30_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_11_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_95_mx0w1,
          and_dcpl_999);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_11_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_11_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_94_mx0w1,
          and_dcpl_999);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_33_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_12_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_98_mx0w1,
          and_dcpl_1011);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_12_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_12_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_97_mx0w1,
          and_dcpl_1011);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_36_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_13_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_101_mx0w1,
          and_dcpl_1023);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_13_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_13_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_100_mx0w1,
          and_dcpl_1023);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_39_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_14_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_104_mx0w1,
          and_dcpl_1035);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_14_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_14_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_103_mx0w1,
          and_dcpl_1035);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_42_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_15_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_107_mx0w1,
          and_dcpl_1047);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_15_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_15_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_106_mx0w1,
          and_dcpl_1047);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_22_13 <= 10'b0;
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_9_0 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_and_45_cse ) begin
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_22_13 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_22_13_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_110_mx0w1,
          and_dcpl_1059);
      FpExpoWidthInc_5U_8U_23U_1U_1U_o_mant_lpi_1_dfm_3_9_0 <= MUX_v_10_2_2(FpMantWidthInc_5U_10U_23U_1U_1U_o_mant_9_0_lpi_1_dfm,
          FpExpoWidthInc_5U_8U_23U_1U_1U_FpExpoWidthInc_5U_8U_23U_1U_1U_or_109_mx0w1,
          and_dcpl_1059);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_1_lpi_1_dfm <= 1'b0;
      IsNaN_8U_23U_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_16_cse ) begin
      IsZero_8U_23U_land_1_lpi_1_dfm <= IsZero_8U_23U_land_1_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_land_1_lpi_1_dfm <= IsNaN_8U_23U_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_2_lpi_1_dfm <= 1'b0;
      IsNaN_8U_23U_land_2_lpi_1_dfm <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_17_cse ) begin
      IsZero_8U_23U_land_2_lpi_1_dfm <= IsZero_8U_23U_land_2_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_land_2_lpi_1_dfm <= IsNaN_8U_23U_land_2_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_3_lpi_1_dfm <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_18_cse ) begin
      IsZero_8U_23U_land_3_lpi_1_dfm <= IsZero_8U_23U_land_3_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_land_3_lpi_1_dfm <= IsNaN_8U_23U_land_3_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_4_lpi_1_dfm <= 1'b0;
      IsNaN_8U_23U_land_4_lpi_1_dfm <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_19_cse ) begin
      IsZero_8U_23U_land_4_lpi_1_dfm <= IsZero_8U_23U_land_4_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_land_4_lpi_1_dfm <= IsNaN_8U_23U_land_4_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_5_lpi_1_dfm <= 1'b0;
      IsNaN_8U_23U_land_5_lpi_1_dfm <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_20_cse ) begin
      IsZero_8U_23U_land_5_lpi_1_dfm <= IsZero_8U_23U_land_5_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_land_5_lpi_1_dfm <= IsNaN_8U_23U_land_5_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_6_lpi_1_dfm <= 1'b0;
      IsNaN_8U_23U_land_6_lpi_1_dfm <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_21_cse ) begin
      IsZero_8U_23U_land_6_lpi_1_dfm <= IsZero_8U_23U_land_6_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_land_6_lpi_1_dfm <= IsNaN_8U_23U_land_6_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_7_lpi_1_dfm <= 1'b0;
      IsNaN_8U_23U_land_7_lpi_1_dfm <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_22_cse ) begin
      IsZero_8U_23U_land_7_lpi_1_dfm <= IsZero_8U_23U_land_7_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_land_7_lpi_1_dfm <= IsNaN_8U_23U_land_7_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_8_lpi_1_dfm <= 1'b0;
      IsNaN_8U_23U_land_8_lpi_1_dfm <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_23_cse ) begin
      IsZero_8U_23U_land_8_lpi_1_dfm <= IsZero_8U_23U_land_8_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_land_8_lpi_1_dfm <= IsNaN_8U_23U_land_8_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_9_lpi_1_dfm <= 1'b0;
      IsNaN_8U_23U_land_9_lpi_1_dfm <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_24_cse ) begin
      IsZero_8U_23U_land_9_lpi_1_dfm <= IsZero_8U_23U_land_9_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_land_9_lpi_1_dfm <= IsNaN_8U_23U_land_9_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_10_lpi_1_dfm <= 1'b0;
      IsNaN_8U_23U_land_10_lpi_1_dfm <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_25_cse ) begin
      IsZero_8U_23U_land_10_lpi_1_dfm <= IsZero_8U_23U_land_10_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_land_10_lpi_1_dfm <= IsNaN_8U_23U_land_10_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_11_lpi_1_dfm <= 1'b0;
      IsNaN_8U_23U_land_11_lpi_1_dfm <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_26_cse ) begin
      IsZero_8U_23U_land_11_lpi_1_dfm <= IsZero_8U_23U_land_11_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_land_11_lpi_1_dfm <= IsNaN_8U_23U_land_11_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_12_lpi_1_dfm <= 1'b0;
      IsNaN_8U_23U_land_12_lpi_1_dfm <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_27_cse ) begin
      IsZero_8U_23U_land_12_lpi_1_dfm <= IsZero_8U_23U_land_12_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_land_12_lpi_1_dfm <= IsNaN_8U_23U_land_12_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_13_lpi_1_dfm <= 1'b0;
      IsNaN_8U_23U_land_13_lpi_1_dfm <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_28_cse ) begin
      IsZero_8U_23U_land_13_lpi_1_dfm <= IsZero_8U_23U_land_13_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_land_13_lpi_1_dfm <= IsNaN_8U_23U_land_13_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_14_lpi_1_dfm <= 1'b0;
      IsNaN_8U_23U_land_14_lpi_1_dfm <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_29_cse ) begin
      IsZero_8U_23U_land_14_lpi_1_dfm <= IsZero_8U_23U_land_14_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_land_14_lpi_1_dfm <= IsNaN_8U_23U_land_14_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_15_lpi_1_dfm <= 1'b0;
      IsNaN_8U_23U_land_15_lpi_1_dfm <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_30_cse ) begin
      IsZero_8U_23U_land_15_lpi_1_dfm <= IsZero_8U_23U_land_15_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_land_15_lpi_1_dfm <= IsNaN_8U_23U_land_15_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_lpi_1_dfm <= 1'b0;
      IsNaN_8U_23U_land_lpi_1_dfm <= 1'b0;
    end
    else if ( IsZero_8U_23U_aelse_and_31_cse ) begin
      IsZero_8U_23U_land_lpi_1_dfm <= IsZero_8U_23U_land_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_land_lpi_1_dfm <= IsNaN_8U_23U_land_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_15_sva_8 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1565_nl) ) begin
      MulOut_data_15_sva_8 <= conv_s2u_49_49($signed((MulIn_data_sva_533[527:495]))
          * $signed(({else_MulOp_data_15_15_lpi_1_dfm_mx0 , else_MulOp_data_15_14_10_lpi_1_dfm_mx0
          , else_MulOp_data_15_9_0_lpi_1_dfm_mx0})));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_14_sva_8 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1567_nl) ) begin
      MulOut_data_14_sva_8 <= conv_s2u_49_49($signed((MulIn_data_sva_533[494:462]))
          * $signed(({else_MulOp_data_14_15_lpi_1_dfm_mx0 , else_MulOp_data_14_14_10_lpi_1_dfm_mx0
          , else_MulOp_data_14_9_0_lpi_1_dfm_mx0})));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_13_sva_8 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1569_nl) ) begin
      MulOut_data_13_sva_8 <= conv_s2u_49_49($signed((MulIn_data_sva_533[461:429]))
          * $signed(({else_MulOp_data_13_15_lpi_1_dfm_mx0 , else_MulOp_data_13_14_10_lpi_1_dfm_mx0
          , else_MulOp_data_13_9_0_lpi_1_dfm_mx0})));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_12_sva_8 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1571_nl) ) begin
      MulOut_data_12_sva_8 <= conv_s2u_49_49($signed((MulIn_data_sva_533[428:396]))
          * $signed(({else_MulOp_data_12_15_lpi_1_dfm_mx0 , else_MulOp_data_12_14_10_lpi_1_dfm_mx0
          , else_MulOp_data_12_9_0_lpi_1_dfm_mx0})));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_11_sva_8 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1573_nl) ) begin
      MulOut_data_11_sva_8 <= conv_s2u_49_49($signed((MulIn_data_sva_533[395:363]))
          * $signed(({else_MulOp_data_11_15_lpi_1_dfm_mx0 , else_MulOp_data_11_14_10_lpi_1_dfm_mx0
          , else_MulOp_data_11_9_0_lpi_1_dfm_mx0})));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_10_sva_8 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1575_nl) ) begin
      MulOut_data_10_sva_8 <= conv_s2u_49_49($signed((MulIn_data_sva_533[362:330]))
          * $signed(({else_MulOp_data_10_15_lpi_1_dfm_mx0 , else_MulOp_data_10_14_10_lpi_1_dfm_mx0
          , else_MulOp_data_10_9_0_lpi_1_dfm_mx0})));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_9_sva_8 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1577_nl) ) begin
      MulOut_data_9_sva_8 <= conv_s2u_49_49($signed((MulIn_data_sva_533[329:297]))
          * $signed(({else_MulOp_data_9_15_lpi_1_dfm_mx0 , else_MulOp_data_9_14_10_lpi_1_dfm_mx0
          , else_MulOp_data_9_9_0_lpi_1_dfm_mx0})));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_8_sva_8 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1579_nl) ) begin
      MulOut_data_8_sva_8 <= conv_s2u_49_49($signed((MulIn_data_sva_533[296:264]))
          * $signed(({else_MulOp_data_8_15_lpi_1_dfm_mx0 , else_MulOp_data_8_14_10_lpi_1_dfm_mx0
          , else_MulOp_data_8_9_0_lpi_1_dfm_mx0})));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_7_sva_8 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1581_nl) ) begin
      MulOut_data_7_sva_8 <= conv_s2u_49_49($signed((MulIn_data_sva_533[263:231]))
          * $signed(({else_MulOp_data_7_15_lpi_1_dfm_mx0 , else_MulOp_data_7_14_10_lpi_1_dfm_mx0
          , else_MulOp_data_7_9_0_lpi_1_dfm_mx0})));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_6_sva_8 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1583_nl) ) begin
      MulOut_data_6_sva_8 <= conv_s2u_49_49($signed((MulIn_data_sva_533[230:198]))
          * $signed(({else_MulOp_data_6_15_lpi_1_dfm_mx0 , else_MulOp_data_6_14_10_lpi_1_dfm_mx0
          , else_MulOp_data_6_9_0_lpi_1_dfm_mx0})));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_5_sva_8 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1585_nl) ) begin
      MulOut_data_5_sva_8 <= conv_s2u_49_49($signed((MulIn_data_sva_533[197:165]))
          * $signed(({else_MulOp_data_5_15_lpi_1_dfm_mx0 , else_MulOp_data_5_14_10_lpi_1_dfm_mx0
          , else_MulOp_data_5_9_0_lpi_1_dfm_mx0})));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_4_sva_8 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1587_nl) ) begin
      MulOut_data_4_sva_8 <= conv_s2u_49_49($signed((MulIn_data_sva_533[164:132]))
          * $signed(({else_MulOp_data_4_15_lpi_1_dfm_mx0 , else_MulOp_data_4_14_10_lpi_1_dfm_mx0
          , else_MulOp_data_4_9_0_lpi_1_dfm_mx0})));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_3_sva_8 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1589_nl) ) begin
      MulOut_data_3_sva_8 <= conv_s2u_49_49($signed((MulIn_data_sva_533[131:99]))
          * $signed(({else_MulOp_data_3_15_lpi_1_dfm_mx0 , else_MulOp_data_3_14_10_lpi_1_dfm_mx0
          , else_MulOp_data_3_9_0_lpi_1_dfm_mx0})));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_2_sva_8 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1591_nl) ) begin
      MulOut_data_2_sva_8 <= conv_s2u_49_49($signed((MulIn_data_sva_533[98:66]))
          * $signed(({else_MulOp_data_2_15_lpi_1_dfm_mx0 , else_MulOp_data_2_14_10_lpi_1_dfm_mx0
          , else_MulOp_data_2_9_0_lpi_1_dfm_mx0})));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_1_sva_8 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1593_nl) ) begin
      MulOut_data_1_sva_8 <= conv_s2u_49_49($signed((MulIn_data_sva_533[65:33]))
          * $signed(({else_MulOp_data_1_15_lpi_1_dfm_mx0 , else_MulOp_data_1_14_10_lpi_1_dfm_mx0
          , else_MulOp_data_1_9_0_lpi_1_dfm_mx0})));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulOut_data_0_sva_8 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1595_nl) ) begin
      MulOut_data_0_sva_8 <= conv_s2u_49_49($signed((MulIn_data_sva_533[32:0])) *
          $signed(({else_MulOp_data_0_15_lpi_1_dfm_mx0 , else_MulOp_data_0_14_10_lpi_1_dfm_mx0
          , else_MulOp_data_0_9_0_lpi_1_dfm_mx0})));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_156_itm) ) begin
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_6 <= IsNaN_8U_23U_land_1_lpi_1_dfm_st_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_157_itm) ) begin
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_6 <= IsNaN_8U_23U_land_2_lpi_1_dfm_st_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_158_itm) ) begin
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_6 <= IsNaN_8U_23U_land_3_lpi_1_dfm_st_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_4_lpi_1_dfm_st_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_159_itm) ) begin
      IsNaN_8U_23U_land_4_lpi_1_dfm_st_6 <= IsNaN_8U_23U_land_4_lpi_1_dfm_st_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_5_lpi_1_dfm_st_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_160_itm) ) begin
      IsNaN_8U_23U_land_5_lpi_1_dfm_st_6 <= IsNaN_8U_23U_land_5_lpi_1_dfm_st_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_6_lpi_1_dfm_st_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_161_itm) ) begin
      IsNaN_8U_23U_land_6_lpi_1_dfm_st_6 <= IsNaN_8U_23U_land_6_lpi_1_dfm_st_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_7_lpi_1_dfm_st_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_162_itm) ) begin
      IsNaN_8U_23U_land_7_lpi_1_dfm_st_6 <= IsNaN_8U_23U_land_7_lpi_1_dfm_st_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_8_lpi_1_dfm_st_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_163_itm) ) begin
      IsNaN_8U_23U_land_8_lpi_1_dfm_st_6 <= IsNaN_8U_23U_land_8_lpi_1_dfm_st_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_9_lpi_1_dfm_st_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_164_itm) ) begin
      IsNaN_8U_23U_land_9_lpi_1_dfm_st_6 <= IsNaN_8U_23U_land_9_lpi_1_dfm_st_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_10_lpi_1_dfm_st_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_165_itm) ) begin
      IsNaN_8U_23U_land_10_lpi_1_dfm_st_6 <= IsNaN_8U_23U_land_10_lpi_1_dfm_st_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_11_lpi_1_dfm_st_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_166_itm) ) begin
      IsNaN_8U_23U_land_11_lpi_1_dfm_st_6 <= IsNaN_8U_23U_land_11_lpi_1_dfm_st_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_12_lpi_1_dfm_st_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_167_itm) ) begin
      IsNaN_8U_23U_land_12_lpi_1_dfm_st_6 <= IsNaN_8U_23U_land_12_lpi_1_dfm_st_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_13_lpi_1_dfm_st_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_168_itm) ) begin
      IsNaN_8U_23U_land_13_lpi_1_dfm_st_6 <= IsNaN_8U_23U_land_13_lpi_1_dfm_st_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_14_lpi_1_dfm_st_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_169_itm) ) begin
      IsNaN_8U_23U_land_14_lpi_1_dfm_st_6 <= IsNaN_8U_23U_land_14_lpi_1_dfm_st_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_15_lpi_1_dfm_st_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_170_itm) ) begin
      IsNaN_8U_23U_land_15_lpi_1_dfm_st_6 <= IsNaN_8U_23U_land_15_lpi_1_dfm_st_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_st_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (~ mux_171_itm) ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_st_6 <= IsNaN_8U_23U_land_lpi_1_dfm_st_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_nan_to_zero_op_sign_1_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1596_nl) ) begin
      mul_nan_to_zero_op_sign_1_lpi_1_dfm_4 <= else_MulOp_data_0_15_lpi_1_dfm_mx0
          & (~ mul_nan_to_zero_land_1_lpi_1_dfm);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_nan_to_zero_op_sign_2_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1597_nl) ) begin
      mul_nan_to_zero_op_sign_2_lpi_1_dfm_4 <= else_MulOp_data_1_15_lpi_1_dfm_mx0
          & (~ mul_nan_to_zero_land_2_lpi_1_dfm);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_nan_to_zero_op_sign_3_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1598_nl) ) begin
      mul_nan_to_zero_op_sign_3_lpi_1_dfm_4 <= else_MulOp_data_2_15_lpi_1_dfm_mx0
          & (~ mul_nan_to_zero_land_3_lpi_1_dfm);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_nan_to_zero_op_sign_4_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1599_nl) ) begin
      mul_nan_to_zero_op_sign_4_lpi_1_dfm_4 <= else_MulOp_data_3_15_lpi_1_dfm_mx0
          & (~ mul_nan_to_zero_land_4_lpi_1_dfm);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_nan_to_zero_op_sign_5_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1600_nl) ) begin
      mul_nan_to_zero_op_sign_5_lpi_1_dfm_4 <= else_MulOp_data_4_15_lpi_1_dfm_mx0
          & (~ mul_nan_to_zero_land_5_lpi_1_dfm);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_nan_to_zero_op_sign_6_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1601_nl) ) begin
      mul_nan_to_zero_op_sign_6_lpi_1_dfm_4 <= else_MulOp_data_5_15_lpi_1_dfm_mx0
          & (~ mul_nan_to_zero_land_6_lpi_1_dfm);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_nan_to_zero_op_sign_7_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1602_nl) ) begin
      mul_nan_to_zero_op_sign_7_lpi_1_dfm_4 <= else_MulOp_data_6_15_lpi_1_dfm_mx0
          & (~ mul_nan_to_zero_land_7_lpi_1_dfm);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_nan_to_zero_op_sign_8_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1603_nl) ) begin
      mul_nan_to_zero_op_sign_8_lpi_1_dfm_4 <= else_MulOp_data_7_15_lpi_1_dfm_mx0
          & (~ mul_nan_to_zero_land_8_lpi_1_dfm);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_nan_to_zero_op_sign_9_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1604_nl) ) begin
      mul_nan_to_zero_op_sign_9_lpi_1_dfm_4 <= else_MulOp_data_8_15_lpi_1_dfm_mx0
          & (~ mul_nan_to_zero_land_9_lpi_1_dfm);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_nan_to_zero_op_sign_10_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1605_nl) ) begin
      mul_nan_to_zero_op_sign_10_lpi_1_dfm_4 <= else_MulOp_data_9_15_lpi_1_dfm_mx0
          & (~ mul_nan_to_zero_land_10_lpi_1_dfm);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_nan_to_zero_op_sign_11_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1606_nl) ) begin
      mul_nan_to_zero_op_sign_11_lpi_1_dfm_4 <= else_MulOp_data_10_15_lpi_1_dfm_mx0
          & (~ mul_nan_to_zero_land_11_lpi_1_dfm);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_nan_to_zero_op_sign_12_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1607_nl) ) begin
      mul_nan_to_zero_op_sign_12_lpi_1_dfm_4 <= else_MulOp_data_11_15_lpi_1_dfm_mx0
          & (~ mul_nan_to_zero_land_12_lpi_1_dfm);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_nan_to_zero_op_sign_13_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1608_nl) ) begin
      mul_nan_to_zero_op_sign_13_lpi_1_dfm_4 <= else_MulOp_data_12_15_lpi_1_dfm_mx0
          & (~ mul_nan_to_zero_land_13_lpi_1_dfm);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_nan_to_zero_op_sign_14_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1609_nl) ) begin
      mul_nan_to_zero_op_sign_14_lpi_1_dfm_4 <= else_MulOp_data_13_15_lpi_1_dfm_mx0
          & (~ mul_nan_to_zero_land_14_lpi_1_dfm);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_nan_to_zero_op_sign_15_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1610_nl) ) begin
      mul_nan_to_zero_op_sign_15_lpi_1_dfm_4 <= else_MulOp_data_14_15_lpi_1_dfm_mx0
          & (~ mul_nan_to_zero_land_15_lpi_1_dfm);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_nan_to_zero_op_sign_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_50) & (mux_1611_nl) ) begin
      mul_nan_to_zero_op_sign_lpi_1_dfm_4 <= else_MulOp_data_15_15_lpi_1_dfm_mx0
          & (~ mul_nan_to_zero_land_lpi_1_dfm);
    end
  end
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_33_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_1_sva[9:0]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_1_lpi_1_dfm[9:0]), mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_32_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_33_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_1_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_33_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_32_nl),
      10'b1111111111, FpMul_8U_23U_lor_33_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_32_nl = MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_1_sva[12:10]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_1_lpi_1_dfm[12:10]), mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_31_nl = ~(MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_32_nl),
      3'b111, FpMul_8U_23U_is_inf_1_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_32_nl = ~(MUX_v_3_2_2((FpMul_8U_23U_nor_31_nl),
      3'b111, FpMul_8U_23U_lor_33_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_34_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_1_sva[22:13]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_1_lpi_1_dfm[22:13]), mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_34_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_1_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_16_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_nl),
      10'b1111111111, FpMul_8U_23U_lor_33_lpi_1_dfm));
  assign SetToInf_8U_23U_mux_nl = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_lpi_1_dfm_1[3:0]),
      FpMul_8U_23U_FpMul_8U_23U_and_itm_2);
  assign FpMul_8U_23U_oelse_2_not_64_nl = ~ FpMul_8U_23U_lor_33_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_95_nl = MUX_v_4_2_2(4'b0000, (SetToInf_8U_23U_mux_nl),
      (FpMul_8U_23U_oelse_2_not_64_nl));
  assign FpMul_8U_23U_oelse_2_not_96_nl = ~ FpMul_8U_23U_lor_33_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_97_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_1_lpi_1_dfm[1:0]),
      (FpMul_8U_23U_oelse_2_not_96_nl));
  assign FpMul_8U_23U_oelse_2_not_112_nl = ~ FpMul_8U_23U_lor_33_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_96_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_1_lpi_1_dfm[3:2]),
      (FpMul_8U_23U_oelse_2_not_112_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_35_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_2_sva[9:0]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_2_lpi_1_dfm[9:0]), mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_34_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_35_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_2_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_35_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_34_nl),
      10'b1111111111, FpMul_8U_23U_lor_34_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_36_nl = MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_2_sva[12:10]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_2_lpi_1_dfm[12:10]), mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_33_nl = ~(MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_36_nl),
      3'b111, FpMul_8U_23U_is_inf_2_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_34_nl = ~(MUX_v_3_2_2((FpMul_8U_23U_nor_33_nl),
      3'b111, FpMul_8U_23U_lor_34_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_37_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_2_sva[22:13]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_2_lpi_1_dfm[22:13]), mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_16_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_37_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_2_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_17_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_16_nl),
      10'b1111111111, FpMul_8U_23U_lor_34_lpi_1_dfm));
  assign SetToInf_8U_23U_mux_2_nl = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_lpi_1_dfm_1[3:0]),
      FpMul_8U_23U_FpMul_8U_23U_and_64_itm_2);
  assign FpMul_8U_23U_oelse_2_not_66_nl = ~ FpMul_8U_23U_lor_34_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_98_nl = MUX_v_4_2_2(4'b0000, (SetToInf_8U_23U_mux_2_nl),
      (FpMul_8U_23U_oelse_2_not_66_nl));
  assign FpMul_8U_23U_oelse_2_not_97_nl = ~ FpMul_8U_23U_lor_34_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_100_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_2_lpi_1_dfm[1:0]),
      (FpMul_8U_23U_oelse_2_not_97_nl));
  assign FpMul_8U_23U_oelse_2_not_113_nl = ~ FpMul_8U_23U_lor_34_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_99_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_2_lpi_1_dfm[3:2]),
      (FpMul_8U_23U_oelse_2_not_113_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_38_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_3_sva[9:0]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_3_lpi_1_dfm[9:0]), mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_36_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_38_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_3_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_37_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_36_nl),
      10'b1111111111, FpMul_8U_23U_lor_35_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_39_nl = MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_3_sva[12:10]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_3_lpi_1_dfm[12:10]), mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_35_nl = ~(MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_39_nl),
      3'b111, FpMul_8U_23U_is_inf_3_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_36_nl = ~(MUX_v_3_2_2((FpMul_8U_23U_nor_35_nl),
      3'b111, FpMul_8U_23U_lor_35_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_40_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_3_sva[22:13]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_3_lpi_1_dfm[22:13]), mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_17_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_40_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_3_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_18_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_17_nl),
      10'b1111111111, FpMul_8U_23U_lor_35_lpi_1_dfm));
  assign SetToInf_8U_23U_mux_4_nl = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_lpi_1_dfm_1[3:0]),
      FpMul_8U_23U_FpMul_8U_23U_and_65_itm_2);
  assign FpMul_8U_23U_oelse_2_not_68_nl = ~ FpMul_8U_23U_lor_35_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_101_nl = MUX_v_4_2_2(4'b0000, (SetToInf_8U_23U_mux_4_nl),
      (FpMul_8U_23U_oelse_2_not_68_nl));
  assign FpMul_8U_23U_oelse_2_not_98_nl = ~ FpMul_8U_23U_lor_35_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_103_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_3_lpi_1_dfm[1:0]),
      (FpMul_8U_23U_oelse_2_not_98_nl));
  assign FpMul_8U_23U_oelse_2_not_114_nl = ~ FpMul_8U_23U_lor_35_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_102_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_3_lpi_1_dfm[3:2]),
      (FpMul_8U_23U_oelse_2_not_114_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_41_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_4_sva[9:0]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_4_lpi_1_dfm[9:0]), mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_38_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_41_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_4_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_39_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_38_nl),
      10'b1111111111, FpMul_8U_23U_lor_36_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_42_nl = MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_4_sva[12:10]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_4_lpi_1_dfm[12:10]), mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_37_nl = ~(MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_42_nl),
      3'b111, FpMul_8U_23U_is_inf_4_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_38_nl = ~(MUX_v_3_2_2((FpMul_8U_23U_nor_37_nl),
      3'b111, FpMul_8U_23U_lor_36_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_43_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_4_sva[22:13]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_4_lpi_1_dfm[22:13]), mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_18_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_43_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_4_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_19_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_18_nl),
      10'b1111111111, FpMul_8U_23U_lor_36_lpi_1_dfm));
  assign SetToInf_8U_23U_mux_6_nl = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_4_lpi_1_dfm_1[3:0]),
      FpMul_8U_23U_FpMul_8U_23U_and_66_itm_2);
  assign FpMul_8U_23U_oelse_2_not_70_nl = ~ FpMul_8U_23U_lor_36_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_104_nl = MUX_v_4_2_2(4'b0000, (SetToInf_8U_23U_mux_6_nl),
      (FpMul_8U_23U_oelse_2_not_70_nl));
  assign FpMul_8U_23U_oelse_2_not_99_nl = ~ FpMul_8U_23U_lor_36_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_106_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_4_lpi_1_dfm[1:0]),
      (FpMul_8U_23U_oelse_2_not_99_nl));
  assign FpMul_8U_23U_oelse_2_not_115_nl = ~ FpMul_8U_23U_lor_36_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_105_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_4_lpi_1_dfm[3:2]),
      (FpMul_8U_23U_oelse_2_not_115_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_44_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_5_sva[9:0]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_5_lpi_1_dfm[9:0]), mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_40_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_44_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_5_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_41_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_40_nl),
      10'b1111111111, FpMul_8U_23U_lor_37_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_45_nl = MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_5_sva[12:10]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_5_lpi_1_dfm[12:10]), mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_39_nl = ~(MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_45_nl),
      3'b111, FpMul_8U_23U_is_inf_5_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_40_nl = ~(MUX_v_3_2_2((FpMul_8U_23U_nor_39_nl),
      3'b111, FpMul_8U_23U_lor_37_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_46_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_5_sva[22:13]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_5_lpi_1_dfm[22:13]), mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_19_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_46_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_5_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_20_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_19_nl),
      10'b1111111111, FpMul_8U_23U_lor_37_lpi_1_dfm));
  assign SetToInf_8U_23U_mux_8_nl = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_5_lpi_1_dfm_1[3:0]),
      FpMul_8U_23U_FpMul_8U_23U_and_67_itm_2);
  assign FpMul_8U_23U_oelse_2_not_72_nl = ~ FpMul_8U_23U_lor_37_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_107_nl = MUX_v_4_2_2(4'b0000, (SetToInf_8U_23U_mux_8_nl),
      (FpMul_8U_23U_oelse_2_not_72_nl));
  assign FpMul_8U_23U_oelse_2_not_100_nl = ~ FpMul_8U_23U_lor_37_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_109_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_5_lpi_1_dfm[1:0]),
      (FpMul_8U_23U_oelse_2_not_100_nl));
  assign FpMul_8U_23U_oelse_2_not_116_nl = ~ FpMul_8U_23U_lor_37_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_108_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_5_lpi_1_dfm[3:2]),
      (FpMul_8U_23U_oelse_2_not_116_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_47_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_6_sva[9:0]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_6_lpi_1_dfm[9:0]), mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_42_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_47_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_6_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_43_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_42_nl),
      10'b1111111111, FpMul_8U_23U_lor_38_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_48_nl = MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_6_sva[12:10]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_6_lpi_1_dfm[12:10]), mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_41_nl = ~(MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_48_nl),
      3'b111, FpMul_8U_23U_is_inf_6_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_42_nl = ~(MUX_v_3_2_2((FpMul_8U_23U_nor_41_nl),
      3'b111, FpMul_8U_23U_lor_38_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_49_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_6_sva[22:13]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_6_lpi_1_dfm[22:13]), mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_20_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_49_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_6_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_21_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_20_nl),
      10'b1111111111, FpMul_8U_23U_lor_38_lpi_1_dfm));
  assign SetToInf_8U_23U_mux_10_nl = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_6_lpi_1_dfm_1[3:0]),
      FpMul_8U_23U_FpMul_8U_23U_and_68_itm_2);
  assign FpMul_8U_23U_oelse_2_not_74_nl = ~ FpMul_8U_23U_lor_38_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_110_nl = MUX_v_4_2_2(4'b0000, (SetToInf_8U_23U_mux_10_nl),
      (FpMul_8U_23U_oelse_2_not_74_nl));
  assign FpMul_8U_23U_oelse_2_not_101_nl = ~ FpMul_8U_23U_lor_38_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_112_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_6_lpi_1_dfm[1:0]),
      (FpMul_8U_23U_oelse_2_not_101_nl));
  assign FpMul_8U_23U_oelse_2_not_117_nl = ~ FpMul_8U_23U_lor_38_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_111_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_6_lpi_1_dfm[3:2]),
      (FpMul_8U_23U_oelse_2_not_117_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_50_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_7_sva[9:0]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_7_lpi_1_dfm[9:0]), mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_44_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_50_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_7_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_45_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_44_nl),
      10'b1111111111, FpMul_8U_23U_lor_39_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_51_nl = MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_7_sva[12:10]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_7_lpi_1_dfm[12:10]), mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_43_nl = ~(MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_51_nl),
      3'b111, FpMul_8U_23U_is_inf_7_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_44_nl = ~(MUX_v_3_2_2((FpMul_8U_23U_nor_43_nl),
      3'b111, FpMul_8U_23U_lor_39_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_52_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_7_sva[22:13]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_7_lpi_1_dfm[22:13]), mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_21_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_52_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_7_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_22_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_21_nl),
      10'b1111111111, FpMul_8U_23U_lor_39_lpi_1_dfm));
  assign SetToInf_8U_23U_mux_12_nl = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_7_lpi_1_dfm_1[3:0]),
      FpMul_8U_23U_FpMul_8U_23U_and_69_itm_2);
  assign FpMul_8U_23U_oelse_2_not_76_nl = ~ FpMul_8U_23U_lor_39_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_113_nl = MUX_v_4_2_2(4'b0000, (SetToInf_8U_23U_mux_12_nl),
      (FpMul_8U_23U_oelse_2_not_76_nl));
  assign FpMul_8U_23U_oelse_2_not_102_nl = ~ FpMul_8U_23U_lor_39_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_115_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_7_lpi_1_dfm[1:0]),
      (FpMul_8U_23U_oelse_2_not_102_nl));
  assign FpMul_8U_23U_oelse_2_not_118_nl = ~ FpMul_8U_23U_lor_39_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_114_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_7_lpi_1_dfm[3:2]),
      (FpMul_8U_23U_oelse_2_not_118_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_53_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_8_sva[9:0]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_8_lpi_1_dfm[9:0]), mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_46_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_53_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_8_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_47_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_46_nl),
      10'b1111111111, FpMul_8U_23U_lor_40_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_54_nl = MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_8_sva[12:10]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_8_lpi_1_dfm[12:10]), mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_45_nl = ~(MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_54_nl),
      3'b111, FpMul_8U_23U_is_inf_8_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_46_nl = ~(MUX_v_3_2_2((FpMul_8U_23U_nor_45_nl),
      3'b111, FpMul_8U_23U_lor_40_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_55_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_8_sva[22:13]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_8_lpi_1_dfm[22:13]), mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_22_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_55_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_8_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_23_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_22_nl),
      10'b1111111111, FpMul_8U_23U_lor_40_lpi_1_dfm));
  assign SetToInf_8U_23U_mux_14_nl = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_8_lpi_1_dfm_1[3:0]),
      FpMul_8U_23U_FpMul_8U_23U_and_70_itm_2);
  assign FpMul_8U_23U_oelse_2_not_78_nl = ~ FpMul_8U_23U_lor_40_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_116_nl = MUX_v_4_2_2(4'b0000, (SetToInf_8U_23U_mux_14_nl),
      (FpMul_8U_23U_oelse_2_not_78_nl));
  assign FpMul_8U_23U_oelse_2_not_103_nl = ~ FpMul_8U_23U_lor_40_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_118_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_8_lpi_1_dfm[1:0]),
      (FpMul_8U_23U_oelse_2_not_103_nl));
  assign FpMul_8U_23U_oelse_2_not_119_nl = ~ FpMul_8U_23U_lor_40_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_117_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_8_lpi_1_dfm[3:2]),
      (FpMul_8U_23U_oelse_2_not_119_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_56_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_9_sva[9:0]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_9_lpi_1_dfm[9:0]), mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_48_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_56_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_9_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_49_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_48_nl),
      10'b1111111111, FpMul_8U_23U_lor_41_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_57_nl = MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_9_sva[12:10]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_9_lpi_1_dfm[12:10]), mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_47_nl = ~(MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_57_nl),
      3'b111, FpMul_8U_23U_is_inf_9_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_48_nl = ~(MUX_v_3_2_2((FpMul_8U_23U_nor_47_nl),
      3'b111, FpMul_8U_23U_lor_41_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_16_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_9_sva[22:13]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_9_lpi_1_dfm[22:13]), mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_23_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_16_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_9_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_24_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_23_nl),
      10'b1111111111, FpMul_8U_23U_lor_41_lpi_1_dfm));
  assign SetToInf_8U_23U_mux_16_nl = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_9_lpi_1_dfm_1[3:0]),
      FpMul_8U_23U_FpMul_8U_23U_and_71_itm_2);
  assign FpMul_8U_23U_oelse_2_not_80_nl = ~ FpMul_8U_23U_lor_41_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_119_nl = MUX_v_4_2_2(4'b0000, (SetToInf_8U_23U_mux_16_nl),
      (FpMul_8U_23U_oelse_2_not_80_nl));
  assign FpMul_8U_23U_oelse_2_not_104_nl = ~ FpMul_8U_23U_lor_41_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_121_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_9_lpi_1_dfm[1:0]),
      (FpMul_8U_23U_oelse_2_not_104_nl));
  assign FpMul_8U_23U_oelse_2_not_120_nl = ~ FpMul_8U_23U_lor_41_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_120_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_9_lpi_1_dfm[3:2]),
      (FpMul_8U_23U_oelse_2_not_120_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_58_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_10_sva[9:0]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_10_lpi_1_dfm[9:0]), mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_50_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_58_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_10_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_51_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_50_nl),
      10'b1111111111, FpMul_8U_23U_lor_42_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_59_nl = MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_10_sva[12:10]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_10_lpi_1_dfm[12:10]), mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_49_nl = ~(MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_59_nl),
      3'b111, FpMul_8U_23U_is_inf_10_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_50_nl = ~(MUX_v_3_2_2((FpMul_8U_23U_nor_49_nl),
      3'b111, FpMul_8U_23U_lor_42_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_18_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_10_sva[22:13]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_10_lpi_1_dfm[22:13]), mul_loop_mul_10_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_24_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_18_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_10_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_25_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_24_nl),
      10'b1111111111, FpMul_8U_23U_lor_42_lpi_1_dfm));
  assign SetToInf_8U_23U_mux_18_nl = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_10_lpi_1_dfm_1[3:0]),
      FpMul_8U_23U_FpMul_8U_23U_and_72_itm_2);
  assign FpMul_8U_23U_oelse_2_not_82_nl = ~ FpMul_8U_23U_lor_42_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_122_nl = MUX_v_4_2_2(4'b0000, (SetToInf_8U_23U_mux_18_nl),
      (FpMul_8U_23U_oelse_2_not_82_nl));
  assign FpMul_8U_23U_oelse_2_not_105_nl = ~ FpMul_8U_23U_lor_42_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_124_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_10_lpi_1_dfm[1:0]),
      (FpMul_8U_23U_oelse_2_not_105_nl));
  assign FpMul_8U_23U_oelse_2_not_121_nl = ~ FpMul_8U_23U_lor_42_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_123_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_10_lpi_1_dfm[3:2]),
      (FpMul_8U_23U_oelse_2_not_121_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_60_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_11_sva[9:0]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_11_lpi_1_dfm[9:0]), mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_52_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_60_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_11_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_53_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_52_nl),
      10'b1111111111, FpMul_8U_23U_lor_43_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_61_nl = MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_11_sva[12:10]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_11_lpi_1_dfm[12:10]), mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_51_nl = ~(MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_61_nl),
      3'b111, FpMul_8U_23U_is_inf_11_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_52_nl = ~(MUX_v_3_2_2((FpMul_8U_23U_nor_51_nl),
      3'b111, FpMul_8U_23U_lor_43_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_20_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_11_sva[22:13]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_11_lpi_1_dfm[22:13]), mul_loop_mul_11_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_25_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_20_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_11_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_26_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_25_nl),
      10'b1111111111, FpMul_8U_23U_lor_43_lpi_1_dfm));
  assign SetToInf_8U_23U_mux_20_nl = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_11_lpi_1_dfm_1[3:0]),
      FpMul_8U_23U_FpMul_8U_23U_and_73_itm_2);
  assign FpMul_8U_23U_oelse_2_not_84_nl = ~ FpMul_8U_23U_lor_43_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_125_nl = MUX_v_4_2_2(4'b0000, (SetToInf_8U_23U_mux_20_nl),
      (FpMul_8U_23U_oelse_2_not_84_nl));
  assign FpMul_8U_23U_oelse_2_not_106_nl = ~ FpMul_8U_23U_lor_43_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_127_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_11_lpi_1_dfm[1:0]),
      (FpMul_8U_23U_oelse_2_not_106_nl));
  assign FpMul_8U_23U_oelse_2_not_122_nl = ~ FpMul_8U_23U_lor_43_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_126_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_11_lpi_1_dfm[3:2]),
      (FpMul_8U_23U_oelse_2_not_122_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_62_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_12_sva[9:0]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_12_lpi_1_dfm[9:0]), mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_54_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_62_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_12_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_55_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_54_nl),
      10'b1111111111, FpMul_8U_23U_lor_44_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_63_nl = MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_12_sva[12:10]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_12_lpi_1_dfm[12:10]), mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_53_nl = ~(MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_63_nl),
      3'b111, FpMul_8U_23U_is_inf_12_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_54_nl = ~(MUX_v_3_2_2((FpMul_8U_23U_nor_53_nl),
      3'b111, FpMul_8U_23U_lor_44_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_22_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_12_sva[22:13]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_12_lpi_1_dfm[22:13]), mul_loop_mul_12_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_26_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_22_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_12_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_27_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_26_nl),
      10'b1111111111, FpMul_8U_23U_lor_44_lpi_1_dfm));
  assign SetToInf_8U_23U_mux_22_nl = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_12_lpi_1_dfm_1[3:0]),
      FpMul_8U_23U_FpMul_8U_23U_and_74_itm_2);
  assign FpMul_8U_23U_oelse_2_not_86_nl = ~ FpMul_8U_23U_lor_44_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_128_nl = MUX_v_4_2_2(4'b0000, (SetToInf_8U_23U_mux_22_nl),
      (FpMul_8U_23U_oelse_2_not_86_nl));
  assign FpMul_8U_23U_oelse_2_not_107_nl = ~ FpMul_8U_23U_lor_44_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_130_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_12_lpi_1_dfm[1:0]),
      (FpMul_8U_23U_oelse_2_not_107_nl));
  assign FpMul_8U_23U_oelse_2_not_123_nl = ~ FpMul_8U_23U_lor_44_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_129_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_12_lpi_1_dfm[3:2]),
      (FpMul_8U_23U_oelse_2_not_123_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_64_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_13_sva[9:0]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_13_lpi_1_dfm[9:0]), mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_56_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_64_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_13_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_57_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_56_nl),
      10'b1111111111, FpMul_8U_23U_lor_45_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_65_nl = MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_13_sva[12:10]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_13_lpi_1_dfm[12:10]), mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_55_nl = ~(MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_65_nl),
      3'b111, FpMul_8U_23U_is_inf_13_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_56_nl = ~(MUX_v_3_2_2((FpMul_8U_23U_nor_55_nl),
      3'b111, FpMul_8U_23U_lor_45_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_24_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_13_sva[22:13]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_13_lpi_1_dfm[22:13]), mul_loop_mul_13_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_27_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_24_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_13_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_28_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_27_nl),
      10'b1111111111, FpMul_8U_23U_lor_45_lpi_1_dfm));
  assign SetToInf_8U_23U_mux_24_nl = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_13_lpi_1_dfm_1[3:0]),
      FpMul_8U_23U_FpMul_8U_23U_and_75_itm_2);
  assign FpMul_8U_23U_oelse_2_not_88_nl = ~ FpMul_8U_23U_lor_45_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_131_nl = MUX_v_4_2_2(4'b0000, (SetToInf_8U_23U_mux_24_nl),
      (FpMul_8U_23U_oelse_2_not_88_nl));
  assign FpMul_8U_23U_oelse_2_not_108_nl = ~ FpMul_8U_23U_lor_45_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_133_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_13_lpi_1_dfm[1:0]),
      (FpMul_8U_23U_oelse_2_not_108_nl));
  assign FpMul_8U_23U_oelse_2_not_124_nl = ~ FpMul_8U_23U_lor_45_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_132_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_13_lpi_1_dfm[3:2]),
      (FpMul_8U_23U_oelse_2_not_124_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_66_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_14_sva[9:0]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_14_lpi_1_dfm[9:0]), mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_58_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_66_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_14_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_59_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_58_nl),
      10'b1111111111, FpMul_8U_23U_lor_46_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_67_nl = MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_14_sva[12:10]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_14_lpi_1_dfm[12:10]), mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_57_nl = ~(MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_67_nl),
      3'b111, FpMul_8U_23U_is_inf_14_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_58_nl = ~(MUX_v_3_2_2((FpMul_8U_23U_nor_57_nl),
      3'b111, FpMul_8U_23U_lor_46_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_26_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_14_sva[22:13]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_14_lpi_1_dfm[22:13]), mul_loop_mul_14_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_28_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_26_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_14_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_29_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_28_nl),
      10'b1111111111, FpMul_8U_23U_lor_46_lpi_1_dfm));
  assign SetToInf_8U_23U_mux_26_nl = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_14_lpi_1_dfm_1[3:0]),
      FpMul_8U_23U_FpMul_8U_23U_and_76_itm_2);
  assign FpMul_8U_23U_oelse_2_not_90_nl = ~ FpMul_8U_23U_lor_46_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_134_nl = MUX_v_4_2_2(4'b0000, (SetToInf_8U_23U_mux_26_nl),
      (FpMul_8U_23U_oelse_2_not_90_nl));
  assign FpMul_8U_23U_oelse_2_not_109_nl = ~ FpMul_8U_23U_lor_46_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_136_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_14_lpi_1_dfm[1:0]),
      (FpMul_8U_23U_oelse_2_not_109_nl));
  assign FpMul_8U_23U_oelse_2_not_125_nl = ~ FpMul_8U_23U_lor_46_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_135_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_14_lpi_1_dfm[3:2]),
      (FpMul_8U_23U_oelse_2_not_125_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_68_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_15_sva[9:0]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_15_lpi_1_dfm[9:0]), mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_60_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_68_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_15_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_61_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_60_nl),
      10'b1111111111, FpMul_8U_23U_lor_47_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_69_nl = MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_15_sva[12:10]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_15_lpi_1_dfm[12:10]), mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_59_nl = ~(MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_69_nl),
      3'b111, FpMul_8U_23U_is_inf_15_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_60_nl = ~(MUX_v_3_2_2((FpMul_8U_23U_nor_59_nl),
      3'b111, FpMul_8U_23U_lor_47_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_28_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_15_sva[22:13]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_15_lpi_1_dfm[22:13]), mul_loop_mul_15_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_29_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_28_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_15_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_30_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_29_nl),
      10'b1111111111, FpMul_8U_23U_lor_47_lpi_1_dfm));
  assign SetToInf_8U_23U_mux_28_nl = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_15_lpi_1_dfm_1[3:0]),
      FpMul_8U_23U_FpMul_8U_23U_and_77_itm_2);
  assign FpMul_8U_23U_oelse_2_not_92_nl = ~ FpMul_8U_23U_lor_47_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_137_nl = MUX_v_4_2_2(4'b0000, (SetToInf_8U_23U_mux_28_nl),
      (FpMul_8U_23U_oelse_2_not_92_nl));
  assign FpMul_8U_23U_oelse_2_not_110_nl = ~ FpMul_8U_23U_lor_47_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_139_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_15_lpi_1_dfm[1:0]),
      (FpMul_8U_23U_oelse_2_not_110_nl));
  assign FpMul_8U_23U_oelse_2_not_126_nl = ~ FpMul_8U_23U_lor_47_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_138_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_15_lpi_1_dfm[3:2]),
      (FpMul_8U_23U_oelse_2_not_126_nl));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_70_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_sva[9:0]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_lpi_1_dfm[9:0]), mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_62_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_70_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_63_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_62_nl),
      10'b1111111111, FpMul_8U_23U_lor_2_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_71_nl = MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_sva[12:10]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_lpi_1_dfm[12:10]), mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_61_nl = ~(MUX_v_3_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_71_nl),
      3'b111, FpMul_8U_23U_is_inf_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_62_nl = ~(MUX_v_3_2_2((FpMul_8U_23U_nor_61_nl),
      3'b111, FpMul_8U_23U_lor_2_lpi_1_dfm));
  assign FpMantWidthDec_8U_47U_23U_0U_0U_mux_30_nl = MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_sva[22:13]),
      (FpMantWidthDec_8U_47U_23U_0U_0U_o_mant_lpi_1_dfm[22:13]), mul_loop_mul_16_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_nor_30_nl = ~(MUX_v_10_2_2((FpMantWidthDec_8U_47U_23U_0U_0U_mux_30_nl),
      10'b1111111111, FpMul_8U_23U_is_inf_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_31_nl = ~(MUX_v_10_2_2((FpMul_8U_23U_nor_30_nl),
      10'b1111111111, FpMul_8U_23U_lor_2_lpi_1_dfm));
  assign SetToInf_8U_23U_mux_30_nl = MUX_v_4_2_2(4'b1110, (FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_lpi_1_dfm_1[3:0]),
      FpMul_8U_23U_FpMul_8U_23U_and_78_itm_2);
  assign FpMul_8U_23U_oelse_2_not_94_nl = ~ FpMul_8U_23U_lor_2_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_140_nl = MUX_v_4_2_2(4'b0000, (SetToInf_8U_23U_mux_30_nl),
      (FpMul_8U_23U_oelse_2_not_94_nl));
  assign FpMul_8U_23U_oelse_2_not_111_nl = ~ FpMul_8U_23U_lor_2_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_142_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_lpi_1_dfm[1:0]),
      (FpMul_8U_23U_oelse_2_not_111_nl));
  assign FpMul_8U_23U_oelse_2_not_127_nl = ~ FpMul_8U_23U_lor_2_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_141_nl = MUX_v_2_2_2(2'b00, (FpMul_8U_23U_o_expo_7_4_lpi_1_dfm[3:2]),
      (FpMul_8U_23U_oelse_2_not_127_nl));
  assign mux_16_nl = MUX_s_1_2_2(mux_tmp_8, mux_tmp_1, mul_loop_mul_if_land_1_lpi_1_dfm_st);
  assign mux_17_nl = MUX_s_1_2_2(mux_tmp_8, mux_tmp_1, nor_21_cse);
  assign mux_18_nl = MUX_s_1_2_2((mux_17_nl), (mux_16_nl), or_90_cse);
  assign mux_19_nl = MUX_s_1_2_2(mux_tmp_1, (mux_18_nl), chn_mul_in_rsci_bawt);
  assign mux_26_nl = MUX_s_1_2_2(mux_tmp_18, mux_tmp_14, mul_loop_mul_if_land_2_lpi_1_dfm_st);
  assign mux_27_nl = MUX_s_1_2_2(mux_tmp_18, mux_tmp_14, nor_23_cse);
  assign mux_28_nl = MUX_s_1_2_2((mux_27_nl), (mux_26_nl), or_90_cse);
  assign mux_29_nl = MUX_s_1_2_2(mux_tmp_14, (mux_28_nl), chn_mul_in_rsci_bawt);
  assign mux_36_nl = MUX_s_1_2_2(mux_tmp_28, mux_tmp_24, mul_loop_mul_if_land_3_lpi_1_dfm_st);
  assign mux_37_nl = MUX_s_1_2_2(mux_tmp_28, mux_tmp_24, nor_25_cse);
  assign mux_38_nl = MUX_s_1_2_2((mux_37_nl), (mux_36_nl), or_90_cse);
  assign mux_39_nl = MUX_s_1_2_2(mux_tmp_24, (mux_38_nl), chn_mul_in_rsci_bawt);
  assign mux_46_nl = MUX_s_1_2_2(mux_tmp_38, mux_tmp_34, mul_loop_mul_if_land_4_lpi_1_dfm_st);
  assign mux_47_nl = MUX_s_1_2_2(mux_tmp_38, mux_tmp_34, nor_26_cse);
  assign mux_48_nl = MUX_s_1_2_2((mux_47_nl), (mux_46_nl), or_90_cse);
  assign mux_49_nl = MUX_s_1_2_2(mux_tmp_34, (mux_48_nl), chn_mul_in_rsci_bawt);
  assign mux_56_nl = MUX_s_1_2_2(mux_tmp_48, mux_tmp_44, mul_loop_mul_if_land_5_lpi_1_dfm_st);
  assign mux_57_nl = MUX_s_1_2_2(mux_tmp_48, mux_tmp_44, nor_28_cse);
  assign mux_58_nl = MUX_s_1_2_2((mux_57_nl), (mux_56_nl), or_90_cse);
  assign mux_59_nl = MUX_s_1_2_2(mux_tmp_44, (mux_58_nl), chn_mul_in_rsci_bawt);
  assign mux_63_nl = MUX_s_1_2_2(mux_tmp_55, mux_tmp_53, mul_loop_mul_if_land_6_lpi_1_dfm_st);
  assign mux_64_nl = MUX_s_1_2_2(mux_tmp_55, mux_tmp_53, nor_29_cse);
  assign mux_65_nl = MUX_s_1_2_2((mux_64_nl), (mux_63_nl), or_90_cse);
  assign mux_66_nl = MUX_s_1_2_2(mux_tmp_53, (mux_65_nl), chn_mul_in_rsci_bawt);
  assign mux_70_nl = MUX_s_1_2_2(mux_tmp_62, mux_tmp_60, mul_loop_mul_if_land_7_lpi_1_dfm_st);
  assign mux_71_nl = MUX_s_1_2_2(mux_tmp_62, mux_tmp_60, nor_30_cse);
  assign mux_72_nl = MUX_s_1_2_2((mux_71_nl), (mux_70_nl), or_90_cse);
  assign mux_73_nl = MUX_s_1_2_2(mux_tmp_60, (mux_72_nl), chn_mul_in_rsci_bawt);
  assign mux_80_nl = MUX_s_1_2_2(mux_tmp_72, mux_tmp_68, mul_loop_mul_if_land_8_lpi_1_dfm_st);
  assign mux_81_nl = MUX_s_1_2_2(mux_tmp_72, mux_tmp_68, nor_32_cse);
  assign mux_82_nl = MUX_s_1_2_2((mux_81_nl), (mux_80_nl), or_90_cse);
  assign mux_83_nl = MUX_s_1_2_2(mux_tmp_68, (mux_82_nl), chn_mul_in_rsci_bawt);
  assign mux_90_nl = MUX_s_1_2_2(mux_tmp_82, mux_tmp_78, mul_loop_mul_if_land_9_lpi_1_dfm_st);
  assign mux_91_nl = MUX_s_1_2_2(mux_tmp_82, mux_tmp_78, nor_34_cse);
  assign mux_92_nl = MUX_s_1_2_2((mux_91_nl), (mux_90_nl), or_90_cse);
  assign mux_93_nl = MUX_s_1_2_2(mux_tmp_78, (mux_92_nl), chn_mul_in_rsci_bawt);
  assign mux_97_nl = MUX_s_1_2_2(mux_tmp_89, mux_tmp_87, mul_loop_mul_if_land_10_lpi_1_dfm_st);
  assign mux_98_nl = MUX_s_1_2_2(mux_tmp_89, mux_tmp_87, nor_35_cse);
  assign mux_99_nl = MUX_s_1_2_2((mux_98_nl), (mux_97_nl), or_90_cse);
  assign mux_100_nl = MUX_s_1_2_2(mux_tmp_87, (mux_99_nl), chn_mul_in_rsci_bawt);
  assign mux_104_nl = MUX_s_1_2_2(mux_tmp_96, mux_tmp_94, mul_loop_mul_if_land_11_lpi_1_dfm_st);
  assign mux_105_nl = MUX_s_1_2_2(mux_tmp_96, mux_tmp_94, nor_36_cse);
  assign mux_106_nl = MUX_s_1_2_2((mux_105_nl), (mux_104_nl), or_90_cse);
  assign mux_107_nl = MUX_s_1_2_2(mux_tmp_94, (mux_106_nl), chn_mul_in_rsci_bawt);
  assign mux_111_nl = MUX_s_1_2_2(mux_tmp_103, mux_tmp_101, mul_loop_mul_if_land_12_lpi_1_dfm_st);
  assign mux_112_nl = MUX_s_1_2_2(mux_tmp_103, mux_tmp_101, nor_37_cse);
  assign mux_113_nl = MUX_s_1_2_2((mux_112_nl), (mux_111_nl), or_90_cse);
  assign mux_114_nl = MUX_s_1_2_2(mux_tmp_101, (mux_113_nl), chn_mul_in_rsci_bawt);
  assign mux_121_nl = MUX_s_1_2_2(mux_tmp_113, mux_tmp_109, mul_loop_mul_if_land_13_lpi_1_dfm_st);
  assign mux_122_nl = MUX_s_1_2_2(mux_tmp_113, mux_tmp_109, nor_39_cse);
  assign mux_123_nl = MUX_s_1_2_2((mux_122_nl), (mux_121_nl), or_90_cse);
  assign mux_124_nl = MUX_s_1_2_2(mux_tmp_109, (mux_123_nl), chn_mul_in_rsci_bawt);
  assign mux_128_nl = MUX_s_1_2_2(mux_tmp_120, mux_tmp_118, mul_loop_mul_if_land_14_lpi_1_dfm_st);
  assign mux_129_nl = MUX_s_1_2_2(mux_tmp_120, mux_tmp_118, nor_40_cse);
  assign mux_130_nl = MUX_s_1_2_2((mux_129_nl), (mux_128_nl), or_90_cse);
  assign mux_131_nl = MUX_s_1_2_2(mux_tmp_118, (mux_130_nl), chn_mul_in_rsci_bawt);
  assign mux_138_nl = MUX_s_1_2_2(mux_tmp_130, mux_tmp_126, mul_loop_mul_if_land_15_lpi_1_dfm_st);
  assign mux_139_nl = MUX_s_1_2_2(mux_tmp_130, mux_tmp_126, nor_42_cse);
  assign mux_140_nl = MUX_s_1_2_2((mux_139_nl), (mux_138_nl), or_90_cse);
  assign mux_141_nl = MUX_s_1_2_2(mux_tmp_126, (mux_140_nl), chn_mul_in_rsci_bawt);
  assign mux_148_nl = MUX_s_1_2_2(mux_tmp_140, mux_tmp_136, mul_loop_mul_if_land_lpi_1_dfm_st);
  assign mux_149_nl = MUX_s_1_2_2(mux_tmp_140, mux_tmp_136, nor_44_cse);
  assign mux_150_nl = MUX_s_1_2_2((mux_149_nl), (mux_148_nl), or_90_cse);
  assign mux_151_nl = MUX_s_1_2_2(mux_tmp_136, (mux_150_nl), chn_mul_in_rsci_bawt);
  assign mux_185_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_18_lpi_1_dfm_st, or_312_cse, nor_53_cse);
  assign nor_1489_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_1_lpi_1_dfm_st_6 | (mux_185_nl));
  assign mux_186_nl = MUX_s_1_2_2(nor_1490_cse, (nor_1489_nl), or_309_cse);
  assign or_335_nl = FpMul_8U_23U_lor_19_lpi_1_dfm_st | mul_loop_mul_if_land_2_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign mux_198_nl = MUX_s_1_2_2(or_tmp_248, (or_335_nl), or_309_cse);
  assign or_342_nl = mul_loop_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1 | mul_loop_mul_if_land_2_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2) | reg_FpMul_8U_23U_lor_4_lpi_1_dfm_4_cse;
  assign mux_200_nl = MUX_s_1_2_2(or_tmp_248, (or_342_nl), or_309_cse);
  assign mux_201_nl = MUX_s_1_2_2((mux_200_nl), (mux_198_nl), or_90_cse);
  assign mux_214_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_20_lpi_1_dfm_st, or_363_cse, nor_53_cse);
  assign nor_1475_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_3_lpi_1_dfm_st_6 | (mux_214_nl));
  assign nor_1476_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_3_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_20_lpi_1_dfm_st_3);
  assign mux_215_nl = MUX_s_1_2_2((nor_1476_nl), (nor_1475_nl), or_309_cse);
  assign mux_228_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_21_lpi_1_dfm_st, or_386_cse, nor_53_cse);
  assign nor_1469_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_4_lpi_1_dfm_st_6 | (mux_228_nl));
  assign nor_1470_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_4_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_21_lpi_1_dfm_st_3);
  assign mux_229_nl = MUX_s_1_2_2((nor_1470_nl), (nor_1469_nl), or_309_cse);
  assign or_409_nl = FpMul_8U_23U_lor_22_lpi_1_dfm_st | mul_loop_mul_if_land_5_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign mux_241_nl = MUX_s_1_2_2(or_tmp_322, (or_409_nl), or_309_cse);
  assign or_417_nl = reg_FpMul_8U_23U_lor_7_lpi_1_dfm_4_cse | mul_loop_mul_5_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | mul_loop_mul_if_land_5_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign mux_243_nl = MUX_s_1_2_2(or_tmp_322, (or_417_nl), or_309_cse);
  assign mux_244_nl = MUX_s_1_2_2((mux_243_nl), (mux_241_nl), or_90_cse);
  assign mux_257_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_23_lpi_1_dfm_st, or_438_cse, nor_53_cse);
  assign nor_1459_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_6_lpi_1_dfm_st_6 | (mux_257_nl));
  assign nor_1460_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_6_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_23_lpi_1_dfm_st_3);
  assign mux_258_nl = MUX_s_1_2_2((nor_1460_nl), (nor_1459_nl), or_309_cse);
  assign mux_271_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_24_lpi_1_dfm_st, or_461_cse, nor_53_cse);
  assign nor_1453_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_7_lpi_1_dfm_st_6 | (mux_271_nl));
  assign nor_1454_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_7_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_24_lpi_1_dfm_st_3);
  assign mux_272_nl = MUX_s_1_2_2((nor_1454_nl), (nor_1453_nl), or_309_cse);
  assign or_484_nl = FpMul_8U_23U_lor_25_lpi_1_dfm_st | mul_loop_mul_if_land_8_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign mux_284_nl = MUX_s_1_2_2(or_tmp_397, (or_484_nl), or_309_cse);
  assign or_491_nl = mul_loop_mul_8_FpMul_8U_23U_oelse_1_acc_itm_9_1 | mul_loop_mul_if_land_8_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2) | reg_FpMul_8U_23U_lor_10_lpi_1_dfm_4_cse;
  assign mux_286_nl = MUX_s_1_2_2(or_tmp_397, (or_491_nl), or_309_cse);
  assign mux_287_nl = MUX_s_1_2_2((mux_286_nl), (mux_284_nl), or_90_cse);
  assign or_512_nl = FpMul_8U_23U_lor_26_lpi_1_dfm_st | mul_loop_mul_if_land_9_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign mux_299_nl = MUX_s_1_2_2(or_tmp_425, (or_512_nl), or_309_cse);
  assign or_520_nl = reg_FpMul_8U_23U_lor_11_lpi_1_dfm_4_cse | mul_loop_mul_9_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | mul_loop_mul_if_land_9_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign mux_301_nl = MUX_s_1_2_2(or_tmp_425, (or_520_nl), or_309_cse);
  assign mux_302_nl = MUX_s_1_2_2((mux_301_nl), (mux_299_nl), or_90_cse);
  assign or_541_nl = FpMul_8U_23U_lor_27_lpi_1_dfm_st | mul_loop_mul_if_land_10_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign mux_314_nl = MUX_s_1_2_2(or_tmp_454, (or_541_nl), or_309_cse);
  assign mux_316_nl = MUX_s_1_2_2(or_tmp_454, or_tmp_460, or_309_cse);
  assign mux_317_nl = MUX_s_1_2_2((mux_316_nl), (mux_314_nl), or_90_cse);
  assign mux_330_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_28_lpi_1_dfm_st, or_570_cse, nor_53_cse);
  assign nor_1435_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_11_lpi_1_dfm_st_6 | (mux_330_nl));
  assign nor_1436_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_11_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_28_lpi_1_dfm_st_3);
  assign mux_331_nl = MUX_s_1_2_2((nor_1436_nl), (nor_1435_nl), or_309_cse);
  assign mux_344_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_29_lpi_1_dfm_st, or_593_cse, nor_53_cse);
  assign nor_1429_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_12_lpi_1_dfm_st_6 | (mux_344_nl));
  assign nor_1430_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_12_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_29_lpi_1_dfm_st_3);
  assign mux_345_nl = MUX_s_1_2_2((nor_1430_nl), (nor_1429_nl), or_309_cse);
  assign mux_358_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_30_lpi_1_dfm_st, or_616_cse, nor_53_cse);
  assign nor_1423_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_13_lpi_1_dfm_st_6 | (mux_358_nl));
  assign nor_1424_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_13_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_30_lpi_1_dfm_st_3);
  assign mux_359_nl = MUX_s_1_2_2((nor_1424_nl), (nor_1423_nl), or_309_cse);
  assign mux_372_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_31_lpi_1_dfm_st, or_639_cse, nor_53_cse);
  assign nor_1417_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_14_lpi_1_dfm_st_6 | (mux_372_nl));
  assign nor_1418_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_14_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_31_lpi_1_dfm_st_3);
  assign mux_373_nl = MUX_s_1_2_2((nor_1418_nl), (nor_1417_nl), or_309_cse);
  assign mux_386_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_32_lpi_1_dfm_st, or_662_cse, nor_53_cse);
  assign nor_1411_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_15_lpi_1_dfm_st_6 | (mux_386_nl));
  assign nor_1412_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_15_lpi_1_dfm_st_7 | FpMul_8U_23U_lor_32_lpi_1_dfm_st_3);
  assign mux_387_nl = MUX_s_1_2_2((nor_1412_nl), (nor_1411_nl), or_309_cse);
  assign or_685_nl = FpMul_8U_23U_lor_1_lpi_1_dfm_st | mul_loop_mul_if_land_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign mux_399_nl = MUX_s_1_2_2(or_tmp_598, (or_685_nl), or_309_cse);
  assign or_692_nl = mul_loop_mul_16_FpMul_8U_23U_oelse_1_acc_itm_9_1 | mul_loop_mul_if_land_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2) | reg_FpMul_8U_23U_lor_lpi_1_dfm_4_cse;
  assign mux_401_nl = MUX_s_1_2_2(or_tmp_598, (or_692_nl), or_309_cse);
  assign mux_402_nl = MUX_s_1_2_2((mux_401_nl), (mux_399_nl), or_90_cse);
  assign or_707_nl = mul_loop_mul_if_land_1_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | (~ main_stage_v_4);
  assign mux_408_nl = MUX_s_1_2_2((or_707_nl), mux_tmp_399, or_309_cse);
  assign or_713_nl = (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt
      | mux_tmp_402;
  assign mux_411_nl = MUX_s_1_2_2(mux_tmp_402, mux_tmp_403, or_309_cse);
  assign mux_412_nl = MUX_s_1_2_2((mux_411_nl), (or_713_nl), mul_loop_mul_else_land_1_lpi_1_dfm_9);
  assign or_726_nl = mul_loop_mul_if_land_2_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | (~ main_stage_v_4);
  assign mux_415_nl = MUX_s_1_2_2((or_726_nl), mux_tmp_406, or_309_cse);
  assign or_732_nl = (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt
      | mux_tmp_409;
  assign mux_417_nl = MUX_s_1_2_2(mux_tmp_409, mux_tmp_403, or_309_cse);
  assign mux_418_nl = MUX_s_1_2_2((mux_417_nl), (or_732_nl), mul_loop_mul_else_land_2_lpi_1_dfm_9);
  assign or_742_nl = mul_loop_mul_if_land_3_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | (~ main_stage_v_4);
  assign mux_421_nl = MUX_s_1_2_2((or_742_nl), mux_tmp_412, or_309_cse);
  assign or_751_nl = mul_loop_mul_else_land_3_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_424_nl = MUX_s_1_2_2((or_751_nl), mux_tmp_415, or_309_cse);
  assign or_760_nl = mul_loop_mul_if_land_4_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | (~ main_stage_v_4);
  assign mux_427_nl = MUX_s_1_2_2((or_760_nl), mux_tmp_418, or_309_cse);
  assign or_769_nl = mul_loop_mul_else_land_4_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_430_nl = MUX_s_1_2_2((or_769_nl), mux_tmp_421, or_309_cse);
  assign or_778_nl = mul_loop_mul_if_land_5_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | (~ main_stage_v_4);
  assign mux_433_nl = MUX_s_1_2_2((or_778_nl), mux_tmp_424, or_309_cse);
  assign or_787_nl = mul_loop_mul_else_land_5_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_436_nl = MUX_s_1_2_2((or_787_nl), mux_tmp_427, or_309_cse);
  assign or_796_nl = mul_loop_mul_if_land_6_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | (~ main_stage_v_4);
  assign mux_439_nl = MUX_s_1_2_2((or_796_nl), mux_tmp_430, or_309_cse);
  assign or_805_nl = mul_loop_mul_else_land_6_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_442_nl = MUX_s_1_2_2((or_805_nl), mux_tmp_433, or_309_cse);
  assign or_814_nl = mul_loop_mul_if_land_7_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | (~ main_stage_v_4);
  assign mux_445_nl = MUX_s_1_2_2((or_814_nl), mux_tmp_436, or_309_cse);
  assign or_823_nl = mul_loop_mul_else_land_7_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_448_nl = MUX_s_1_2_2((or_823_nl), mux_tmp_439, or_309_cse);
  assign or_832_nl = mul_loop_mul_if_land_8_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | (~ main_stage_v_4);
  assign mux_451_nl = MUX_s_1_2_2((or_832_nl), mux_tmp_442, or_309_cse);
  assign or_841_nl = mul_loop_mul_else_land_8_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_454_nl = MUX_s_1_2_2((or_841_nl), mux_tmp_445, or_309_cse);
  assign or_850_nl = mul_loop_mul_if_land_9_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | (~ main_stage_v_4);
  assign mux_457_nl = MUX_s_1_2_2((or_850_nl), mux_tmp_448, or_309_cse);
  assign or_859_nl = mul_loop_mul_else_land_9_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_460_nl = MUX_s_1_2_2((or_859_nl), mux_tmp_451, or_309_cse);
  assign or_868_nl = mul_loop_mul_if_land_10_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | (~ main_stage_v_4);
  assign mux_463_nl = MUX_s_1_2_2((or_868_nl), mux_tmp_454, or_309_cse);
  assign or_877_nl = mul_loop_mul_else_land_10_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_466_nl = MUX_s_1_2_2((or_877_nl), mux_tmp_457, or_309_cse);
  assign or_886_nl = mul_loop_mul_if_land_11_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | (~ main_stage_v_4);
  assign mux_469_nl = MUX_s_1_2_2((or_886_nl), mux_tmp_460, or_309_cse);
  assign or_892_nl = (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt
      | mux_tmp_463;
  assign mux_471_nl = MUX_s_1_2_2(mux_tmp_463, mux_tmp_403, or_309_cse);
  assign mux_472_nl = MUX_s_1_2_2((mux_471_nl), (or_892_nl), mul_loop_mul_else_land_11_lpi_1_dfm_9);
  assign or_902_nl = mul_loop_mul_if_land_12_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | (~ main_stage_v_4);
  assign mux_475_nl = MUX_s_1_2_2((or_902_nl), mux_tmp_466, or_309_cse);
  assign or_908_nl = (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt
      | mux_tmp_469;
  assign mux_477_nl = MUX_s_1_2_2(mux_tmp_469, mux_tmp_403, or_309_cse);
  assign mux_478_nl = MUX_s_1_2_2((mux_477_nl), (or_908_nl), mul_loop_mul_else_land_12_lpi_1_dfm_9);
  assign or_918_nl = mul_loop_mul_if_land_13_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | (~ main_stage_v_4);
  assign mux_481_nl = MUX_s_1_2_2((or_918_nl), mux_tmp_472, or_309_cse);
  assign or_924_nl = (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt
      | mux_tmp_475;
  assign mux_483_nl = MUX_s_1_2_2(mux_tmp_475, mux_tmp_403, or_309_cse);
  assign mux_484_nl = MUX_s_1_2_2((mux_483_nl), (or_924_nl), mul_loop_mul_else_land_13_lpi_1_dfm_9);
  assign or_934_nl = mul_loop_mul_if_land_14_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | (~ main_stage_v_4);
  assign mux_487_nl = MUX_s_1_2_2((or_934_nl), mux_tmp_478, or_309_cse);
  assign or_940_nl = (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt
      | mux_tmp_481;
  assign mux_489_nl = MUX_s_1_2_2(mux_tmp_481, mux_tmp_403, or_309_cse);
  assign mux_490_nl = MUX_s_1_2_2((mux_489_nl), (or_940_nl), mul_loop_mul_else_land_14_lpi_1_dfm_9);
  assign or_950_nl = mul_loop_mul_if_land_15_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | (~ main_stage_v_4);
  assign mux_493_nl = MUX_s_1_2_2((or_950_nl), mux_tmp_484, or_309_cse);
  assign or_956_nl = (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt
      | mux_tmp_487;
  assign mux_495_nl = MUX_s_1_2_2(mux_tmp_487, mux_tmp_403, or_309_cse);
  assign mux_496_nl = MUX_s_1_2_2((mux_495_nl), (or_956_nl), mul_loop_mul_else_land_15_lpi_1_dfm_9);
  assign or_966_nl = mul_loop_mul_if_land_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | (~ main_stage_v_4);
  assign mux_499_nl = MUX_s_1_2_2((or_966_nl), mux_tmp_490, or_309_cse);
  assign or_975_nl = mul_loop_mul_else_land_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_502_nl = MUX_s_1_2_2((or_975_nl), mux_tmp_493, or_309_cse);
  assign nor_1676_nl = ~(IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 | FpMul_8U_23U_lor_18_lpi_1_dfm_st_3
      | not_tmp_1326);
  assign or_4963_nl = IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 | (~(FpMul_8U_23U_lor_18_lpi_1_dfm_st_3
      | not_tmp_1326));
  assign mux_1693_nl = MUX_s_1_2_2((or_4963_nl), (nor_1676_nl), IsNaN_8U_23U_land_1_lpi_1_dfm_st_7);
  assign nor_1393_nl = ~((~((~ (mul_loop_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 | FpMul_8U_23U_lor_18_lpi_1_dfm_6))
      | IsNaN_8U_23U_land_1_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8
      | mul_loop_mul_if_land_1_lpi_1_dfm_9);
  assign nor_1395_nl = ~((~ FpMul_8U_23U_lor_18_lpi_1_dfm_6) | IsNaN_8U_23U_land_1_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 | mul_loop_mul_if_land_1_lpi_1_dfm_9);
  assign mux_510_nl = MUX_s_1_2_2((nor_1395_nl), (nor_1393_nl), mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign nor_1396_nl = ~((~ or_tmp_893) | IsNaN_8U_23U_land_1_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 | mul_loop_mul_if_land_1_lpi_1_dfm_9);
  assign mux_511_nl = MUX_s_1_2_2((nor_1396_nl), (mux_510_nl), nor_53_cse);
  assign and_2230_nl = nor_129_cse & (mux_511_nl);
  assign nor_1397_nl = ~((~ main_stage_v_4) | IsNaN_8U_23U_land_1_lpi_1_dfm_11 |
      mul_loop_mul_if_land_1_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | mul_loop_mul_if_land_1_lpi_1_dfm_st_8 | IsNaN_8U_23U_1_land_1_lpi_1_dfm_9
      | FpMul_8U_23U_lor_18_lpi_1_dfm_st_4 | (~(mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
      & or_tmp_898 & ((~ mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs_2) | mul_loop_mul_1_FpMantRNE_48U_24U_else_and_svs_st_2))));
  assign mux_512_nl = MUX_s_1_2_2((nor_1397_nl), (and_2230_nl), or_309_cse);
  assign nor_1390_nl = ~(FpMul_8U_23U_lor_18_lpi_1_dfm_st_4 | mul_loop_mul_if_land_1_lpi_1_dfm_st_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4));
  assign mux_514_nl = MUX_s_1_2_2((nor_1390_nl), nor_1490_cse, or_309_cse);
  assign or_1023_nl = mul_loop_mul_if_land_1_lpi_1_dfm_st_8 | mul_loop_mul_if_land_1_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_515_nl = MUX_s_1_2_2((or_1023_nl), or_tmp_932, or_309_cse);
  assign nor_1381_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_1_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_1_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 | mul_loop_mul_if_land_1_lpi_1_dfm_9);
  assign nor_1382_nl = ~(nor_1383_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_1_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_1_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 | mul_loop_mul_if_land_1_lpi_1_dfm_9);
  assign nor_1384_nl = ~((FpMul_8U_23U_p_mant_p1_1_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_1_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_1_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8
      | mul_loop_mul_if_land_1_lpi_1_dfm_9);
  assign mux_517_nl = MUX_s_1_2_2((nor_1384_nl), (nor_1382_nl), nor_133_cse);
  assign and_2229_nl = mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_517_nl);
  assign nor_1385_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_1_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_1_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8
      | mul_loop_mul_if_land_1_lpi_1_dfm_9);
  assign mux_518_nl = MUX_s_1_2_2((nor_1385_nl), (and_2229_nl), nor_53_cse);
  assign mux_519_nl = MUX_s_1_2_2((mux_518_nl), (nor_1381_nl), FpMul_8U_23U_lor_18_lpi_1_dfm_6);
  assign nor_1386_nl = ~((~ or_tmp_898) | (~ main_stage_v_4) | IsNaN_8U_23U_land_1_lpi_1_dfm_11
      | mul_loop_mul_if_land_1_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_8 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_1_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_1_lpi_1_dfm_9);
  assign mux_520_nl = MUX_s_1_2_2((nor_1386_nl), (mux_519_nl), or_309_cse);
  assign nor_1671_nl = ~(IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 | FpMul_8U_23U_lor_19_lpi_1_dfm_st_3
      | not_tmp_1344);
  assign or_4960_nl = IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 | (~(FpMul_8U_23U_lor_19_lpi_1_dfm_st_3
      | not_tmp_1344));
  assign mux_1698_nl = MUX_s_1_2_2((or_4960_nl), (nor_1671_nl), IsNaN_8U_23U_land_2_lpi_1_dfm_st_7);
  assign nor_1359_nl = ~((~((~ (mul_loop_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 | FpMul_8U_23U_lor_19_lpi_1_dfm_6))
      | IsNaN_8U_23U_land_2_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_2_lpi_1_dfm_8
      | mul_loop_mul_if_land_2_lpi_1_dfm_9);
  assign nor_1361_nl = ~((~ FpMul_8U_23U_lor_19_lpi_1_dfm_6) | IsNaN_8U_23U_land_2_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 | mul_loop_mul_if_land_2_lpi_1_dfm_9);
  assign mux_534_nl = MUX_s_1_2_2((nor_1361_nl), (nor_1359_nl), mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign nor_1362_nl = ~((~ or_tmp_975) | IsNaN_8U_23U_land_2_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 | mul_loop_mul_if_land_2_lpi_1_dfm_9);
  assign mux_535_nl = MUX_s_1_2_2((nor_1362_nl), (mux_534_nl), nor_53_cse);
  assign and_2224_nl = nor_145_cse & (mux_535_nl);
  assign nor_1363_nl = ~((~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8 |
      IsNaN_8U_23U_land_2_lpi_1_dfm_11 | mul_loop_mul_if_land_2_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | mul_loop_mul_if_land_2_lpi_1_dfm_st_8 | IsNaN_8U_23U_1_land_2_lpi_1_dfm_9
      | FpMul_8U_23U_lor_19_lpi_1_dfm_st_4 | (~(mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
      & or_tmp_980 & ((~ mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs_2) | mul_loop_mul_2_FpMantRNE_48U_24U_else_and_svs_st_2))));
  assign mux_536_nl = MUX_s_1_2_2((nor_1363_nl), (and_2224_nl), or_309_cse);
  assign or_1098_nl = FpMul_8U_23U_lor_19_lpi_1_dfm_st_4 | mul_loop_mul_if_land_2_lpi_1_dfm_st_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_538_nl = MUX_s_1_2_2((or_1098_nl), or_tmp_248, or_309_cse);
  assign or_1103_nl = mul_loop_mul_if_land_2_lpi_1_dfm_st_8 | mul_loop_mul_if_land_2_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_539_nl = MUX_s_1_2_2((or_1103_nl), or_tmp_1012, or_309_cse);
  assign nor_1349_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_2_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_2_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 | mul_loop_mul_if_land_2_lpi_1_dfm_9);
  assign nor_1350_nl = ~(nor_1351_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_2_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_2_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 | mul_loop_mul_if_land_2_lpi_1_dfm_9);
  assign nor_1352_nl = ~((FpMul_8U_23U_p_mant_p1_2_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_2_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_2_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_2_lpi_1_dfm_8
      | mul_loop_mul_if_land_2_lpi_1_dfm_9);
  assign mux_541_nl = MUX_s_1_2_2((nor_1352_nl), (nor_1350_nl), nor_149_cse);
  assign and_2223_nl = mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_541_nl);
  assign nor_1353_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_64_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_2_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_2_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_2_lpi_1_dfm_8
      | mul_loop_mul_if_land_2_lpi_1_dfm_9);
  assign mux_542_nl = MUX_s_1_2_2((nor_1353_nl), (and_2223_nl), nor_53_cse);
  assign mux_543_nl = MUX_s_1_2_2((mux_542_nl), (nor_1349_nl), FpMul_8U_23U_lor_19_lpi_1_dfm_6);
  assign nor_1354_nl = ~((~ or_tmp_980) | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_2_lpi_1_dfm_11 | mul_loop_mul_if_land_2_lpi_1_dfm_10 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_2_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_2_lpi_1_dfm_9);
  assign mux_544_nl = MUX_s_1_2_2((nor_1354_nl), (mux_543_nl), or_309_cse);
  assign nor_1666_nl = ~(IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 | FpMul_8U_23U_lor_20_lpi_1_dfm_st_3
      | not_tmp_1362);
  assign or_4957_nl = IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 | (~(FpMul_8U_23U_lor_20_lpi_1_dfm_st_3
      | not_tmp_1362));
  assign mux_1703_nl = MUX_s_1_2_2((or_4957_nl), (nor_1666_nl), IsNaN_8U_23U_land_3_lpi_1_dfm_st_7);
  assign nor_1327_nl = ~((~((~ (mul_loop_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 | FpMul_8U_23U_lor_20_lpi_1_dfm_6))
      | IsNaN_8U_23U_land_3_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_3_lpi_1_dfm_8
      | mul_loop_mul_if_land_3_lpi_1_dfm_9);
  assign nor_1329_nl = ~((~ FpMul_8U_23U_lor_20_lpi_1_dfm_6) | IsNaN_8U_23U_land_3_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 | mul_loop_mul_if_land_3_lpi_1_dfm_9);
  assign mux_558_nl = MUX_s_1_2_2((nor_1329_nl), (nor_1327_nl), mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign nor_1330_nl = ~((~ or_tmp_1055) | IsNaN_8U_23U_land_3_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 | mul_loop_mul_if_land_3_lpi_1_dfm_9);
  assign mux_559_nl = MUX_s_1_2_2((nor_1330_nl), (mux_558_nl), nor_53_cse);
  assign and_2218_nl = nor_161_cse & (mux_559_nl);
  assign nor_1331_nl = ~((~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8 |
      IsNaN_8U_23U_land_3_lpi_1_dfm_11 | mul_loop_mul_if_land_3_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | mul_loop_mul_if_land_3_lpi_1_dfm_st_8 | IsNaN_8U_23U_1_land_3_lpi_1_dfm_9
      | FpMul_8U_23U_lor_20_lpi_1_dfm_st_4 | (~(mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
      & or_tmp_1060 & ((~ mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs_2) | mul_loop_mul_3_FpMantRNE_48U_24U_else_and_svs_st_2))));
  assign mux_560_nl = MUX_s_1_2_2((nor_1331_nl), (and_2218_nl), or_309_cse);
  assign nor_1323_nl = ~(or_tmp_1088 | (~ main_stage_v_3));
  assign nor_1324_nl = ~(FpMul_8U_23U_lor_20_lpi_1_dfm_st_4 | mul_loop_mul_if_land_3_lpi_1_dfm_st_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4));
  assign mux_562_nl = MUX_s_1_2_2((nor_1324_nl), (nor_1323_nl), or_309_cse);
  assign or_1185_nl = mul_loop_mul_if_land_3_lpi_1_dfm_st_8 | mul_loop_mul_if_land_3_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_563_nl = MUX_s_1_2_2((or_1185_nl), or_tmp_1094, or_309_cse);
  assign nor_1315_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_3_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_3_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 | mul_loop_mul_if_land_3_lpi_1_dfm_9);
  assign nor_1316_nl = ~(nor_1317_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_3_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_3_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 | mul_loop_mul_if_land_3_lpi_1_dfm_9);
  assign nor_1318_nl = ~((FpMul_8U_23U_p_mant_p1_3_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_3_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_3_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_3_lpi_1_dfm_8
      | mul_loop_mul_if_land_3_lpi_1_dfm_9);
  assign mux_565_nl = MUX_s_1_2_2((nor_1318_nl), (nor_1316_nl), nor_165_cse);
  assign and_2217_nl = mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_565_nl);
  assign nor_1319_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_65_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_3_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_3_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_3_lpi_1_dfm_8
      | mul_loop_mul_if_land_3_lpi_1_dfm_9);
  assign mux_566_nl = MUX_s_1_2_2((nor_1319_nl), (and_2217_nl), nor_53_cse);
  assign mux_567_nl = MUX_s_1_2_2((mux_566_nl), (nor_1315_nl), FpMul_8U_23U_lor_20_lpi_1_dfm_6);
  assign nor_1320_nl = ~((~ or_tmp_1060) | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_3_lpi_1_dfm_11 | mul_loop_mul_if_land_3_lpi_1_dfm_10 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_3_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_3_lpi_1_dfm_9);
  assign mux_568_nl = MUX_s_1_2_2((nor_1320_nl), (mux_567_nl), or_309_cse);
  assign nor_1661_nl = ~(IsNaN_8U_23U_1_land_4_lpi_1_dfm_8 | FpMul_8U_23U_lor_21_lpi_1_dfm_st_3
      | not_tmp_1380);
  assign or_4954_nl = IsNaN_8U_23U_1_land_4_lpi_1_dfm_8 | (~(FpMul_8U_23U_lor_21_lpi_1_dfm_st_3
      | not_tmp_1380));
  assign mux_1708_nl = MUX_s_1_2_2((or_4954_nl), (nor_1661_nl), IsNaN_8U_23U_land_4_lpi_1_dfm_st_7);
  assign nor_1293_nl = ~((~((~ (mul_loop_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 | FpMul_8U_23U_lor_21_lpi_1_dfm_6))
      | IsNaN_8U_23U_land_4_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_4_lpi_1_dfm_8
      | mul_loop_mul_if_land_4_lpi_1_dfm_9);
  assign nor_1295_nl = ~((~ FpMul_8U_23U_lor_21_lpi_1_dfm_6) | IsNaN_8U_23U_land_4_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_4_lpi_1_dfm_8 | mul_loop_mul_if_land_4_lpi_1_dfm_9);
  assign mux_582_nl = MUX_s_1_2_2((nor_1295_nl), (nor_1293_nl), mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign nor_1296_nl = ~((~ or_tmp_1137) | IsNaN_8U_23U_land_4_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_4_lpi_1_dfm_8 | mul_loop_mul_if_land_4_lpi_1_dfm_9);
  assign mux_583_nl = MUX_s_1_2_2((nor_1296_nl), (mux_582_nl), nor_53_cse);
  assign and_2212_nl = nor_177_cse & (mux_583_nl);
  assign nor_1297_nl = ~((~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8 |
      IsNaN_8U_23U_land_4_lpi_1_dfm_11 | mul_loop_mul_if_land_4_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | mul_loop_mul_if_land_4_lpi_1_dfm_st_8 | IsNaN_8U_23U_1_land_4_lpi_1_dfm_9
      | FpMul_8U_23U_lor_21_lpi_1_dfm_st_4 | (~(mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
      & or_tmp_1142 & ((~ mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs_2) | mul_loop_mul_4_FpMantRNE_48U_24U_else_and_svs_st_2))));
  assign mux_584_nl = MUX_s_1_2_2((nor_1297_nl), (and_2212_nl), or_309_cse);
  assign or_1260_nl = (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt
      | FpMul_8U_23U_lor_21_lpi_1_dfm_st_4 | mul_loop_mul_if_land_4_lpi_1_dfm_st_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign or_1263_nl = FpMul_8U_23U_lor_21_lpi_1_dfm_st_4 | mul_loop_mul_if_land_4_lpi_1_dfm_st_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_587_nl = MUX_s_1_2_2((or_1263_nl), or_tmp_302, or_309_cse);
  assign mux_588_nl = MUX_s_1_2_2((mux_587_nl), (or_1260_nl), FpMul_8U_23U_lor_21_lpi_1_dfm_st_3);
  assign or_1268_nl = mul_loop_mul_if_land_4_lpi_1_dfm_st_8 | mul_loop_mul_if_land_4_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_589_nl = MUX_s_1_2_2((or_1268_nl), or_tmp_1177, or_309_cse);
  assign nor_1285_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_4_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_4_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_4_lpi_1_dfm_8 | mul_loop_mul_if_land_4_lpi_1_dfm_9);
  assign nor_1286_nl = ~(nor_1287_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_4_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_4_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_4_lpi_1_dfm_8 | mul_loop_mul_if_land_4_lpi_1_dfm_9);
  assign nor_1288_nl = ~((FpMul_8U_23U_p_mant_p1_4_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_4_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_4_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_4_lpi_1_dfm_8
      | mul_loop_mul_if_land_4_lpi_1_dfm_9);
  assign mux_591_nl = MUX_s_1_2_2((nor_1288_nl), (nor_1286_nl), nor_181_cse);
  assign and_2211_nl = mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_591_nl);
  assign nor_1289_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_66_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_4_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_4_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_4_lpi_1_dfm_8
      | mul_loop_mul_if_land_4_lpi_1_dfm_9);
  assign mux_592_nl = MUX_s_1_2_2((nor_1289_nl), (and_2211_nl), nor_53_cse);
  assign mux_593_nl = MUX_s_1_2_2((mux_592_nl), (nor_1285_nl), FpMul_8U_23U_lor_21_lpi_1_dfm_6);
  assign nor_1290_nl = ~((~ or_tmp_1142) | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_4_lpi_1_dfm_11 | mul_loop_mul_if_land_4_lpi_1_dfm_10 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_4_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_4_lpi_1_dfm_9);
  assign mux_594_nl = MUX_s_1_2_2((nor_1290_nl), (mux_593_nl), or_309_cse);
  assign nor_1656_nl = ~(IsNaN_8U_23U_1_land_5_lpi_1_dfm_8 | FpMul_8U_23U_lor_22_lpi_1_dfm_st_3
      | not_tmp_1398);
  assign or_4951_nl = IsNaN_8U_23U_1_land_5_lpi_1_dfm_8 | (~(FpMul_8U_23U_lor_22_lpi_1_dfm_st_3
      | not_tmp_1398));
  assign mux_1713_nl = MUX_s_1_2_2((or_4951_nl), (nor_1656_nl), IsNaN_8U_23U_land_5_lpi_1_dfm_st_7);
  assign nor_1263_nl = ~((~((~ (mul_loop_mul_5_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_5_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 | FpMul_8U_23U_lor_22_lpi_1_dfm_6))
      | IsNaN_8U_23U_land_5_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_5_lpi_1_dfm_8
      | mul_loop_mul_if_land_5_lpi_1_dfm_9);
  assign nor_1265_nl = ~((~ FpMul_8U_23U_lor_22_lpi_1_dfm_6) | IsNaN_8U_23U_land_5_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_5_lpi_1_dfm_8 | mul_loop_mul_if_land_5_lpi_1_dfm_9);
  assign mux_608_nl = MUX_s_1_2_2((nor_1265_nl), (nor_1263_nl), mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign nor_1266_nl = ~((~ or_tmp_1220) | IsNaN_8U_23U_land_5_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_5_lpi_1_dfm_8 | mul_loop_mul_if_land_5_lpi_1_dfm_9);
  assign mux_609_nl = MUX_s_1_2_2((nor_1266_nl), (mux_608_nl), nor_53_cse);
  assign and_2206_nl = nor_193_cse & (mux_609_nl);
  assign nor_1267_nl = ~((~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8 |
      IsNaN_8U_23U_land_5_lpi_1_dfm_11 | mul_loop_mul_if_land_5_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | mul_loop_mul_if_land_5_lpi_1_dfm_st_8 | IsNaN_8U_23U_1_land_5_lpi_1_dfm_9
      | FpMul_8U_23U_lor_22_lpi_1_dfm_st_4 | (~(mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
      & or_tmp_1225 & ((~ mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs_2) | mul_loop_mul_5_FpMantRNE_48U_24U_else_and_svs_st_2))));
  assign mux_610_nl = MUX_s_1_2_2((nor_1267_nl), (and_2206_nl), or_309_cse);
  assign or_1343_nl = FpMul_8U_23U_lor_22_lpi_1_dfm_st_4 | mul_loop_mul_if_land_5_lpi_1_dfm_st_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_612_nl = MUX_s_1_2_2((or_1343_nl), or_tmp_322, or_309_cse);
  assign or_1348_nl = mul_loop_mul_if_land_5_lpi_1_dfm_st_8 | mul_loop_mul_if_land_5_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_613_nl = MUX_s_1_2_2((or_1348_nl), or_tmp_1257, or_309_cse);
  assign nor_1253_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_5_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_5_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_5_lpi_1_dfm_8 | mul_loop_mul_if_land_5_lpi_1_dfm_9);
  assign nor_1254_nl = ~(nor_1255_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_5_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_5_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_5_lpi_1_dfm_8 | mul_loop_mul_if_land_5_lpi_1_dfm_9);
  assign nor_1256_nl = ~((FpMul_8U_23U_p_mant_p1_5_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_5_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_5_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_5_lpi_1_dfm_8
      | mul_loop_mul_if_land_5_lpi_1_dfm_9);
  assign mux_615_nl = MUX_s_1_2_2((nor_1256_nl), (nor_1254_nl), nor_197_cse);
  assign and_2205_nl = mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_615_nl);
  assign nor_1257_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_67_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_5_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_5_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_5_lpi_1_dfm_8
      | mul_loop_mul_if_land_5_lpi_1_dfm_9);
  assign mux_616_nl = MUX_s_1_2_2((nor_1257_nl), (and_2205_nl), nor_53_cse);
  assign mux_617_nl = MUX_s_1_2_2((mux_616_nl), (nor_1253_nl), FpMul_8U_23U_lor_22_lpi_1_dfm_6);
  assign nor_1258_nl = ~((~ or_tmp_1225) | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_5_lpi_1_dfm_11 | mul_loop_mul_if_land_5_lpi_1_dfm_10 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_5_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_5_lpi_1_dfm_9);
  assign mux_618_nl = MUX_s_1_2_2((nor_1258_nl), (mux_617_nl), or_309_cse);
  assign nor_1651_nl = ~(IsNaN_8U_23U_1_land_6_lpi_1_dfm_8 | FpMul_8U_23U_lor_23_lpi_1_dfm_st_3
      | not_tmp_1416);
  assign or_4948_nl = IsNaN_8U_23U_1_land_6_lpi_1_dfm_8 | (~(FpMul_8U_23U_lor_23_lpi_1_dfm_st_3
      | not_tmp_1416));
  assign mux_1718_nl = MUX_s_1_2_2((or_4948_nl), (nor_1651_nl), IsNaN_8U_23U_land_6_lpi_1_dfm_st_7);
  assign nor_1231_nl = ~((~((~ (mul_loop_mul_6_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_6_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 | FpMul_8U_23U_lor_23_lpi_1_dfm_6))
      | IsNaN_8U_23U_land_6_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_6_lpi_1_dfm_8
      | mul_loop_mul_if_land_6_lpi_1_dfm_9);
  assign nor_1233_nl = ~((~ FpMul_8U_23U_lor_23_lpi_1_dfm_6) | IsNaN_8U_23U_land_6_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_6_lpi_1_dfm_8 | mul_loop_mul_if_land_6_lpi_1_dfm_9);
  assign mux_632_nl = MUX_s_1_2_2((nor_1233_nl), (nor_1231_nl), mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign nor_1234_nl = ~((~ or_tmp_1300) | IsNaN_8U_23U_land_6_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_6_lpi_1_dfm_8 | mul_loop_mul_if_land_6_lpi_1_dfm_9);
  assign mux_633_nl = MUX_s_1_2_2((nor_1234_nl), (mux_632_nl), nor_53_cse);
  assign and_2200_nl = nor_209_cse & (mux_633_nl);
  assign nor_1235_nl = ~((~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8 |
      IsNaN_8U_23U_land_6_lpi_1_dfm_11 | mul_loop_mul_if_land_6_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | mul_loop_mul_if_land_6_lpi_1_dfm_st_8 | IsNaN_8U_23U_1_land_6_lpi_1_dfm_9
      | FpMul_8U_23U_lor_23_lpi_1_dfm_st_4 | (~(mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
      & or_tmp_1305 & ((~ mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs_2) | mul_loop_mul_6_FpMantRNE_48U_24U_else_and_svs_st_2))));
  assign mux_634_nl = MUX_s_1_2_2((nor_1235_nl), (and_2200_nl), or_309_cse);
  assign nor_1227_nl = ~(or_tmp_1333 | (~ main_stage_v_3));
  assign nor_1228_nl = ~(FpMul_8U_23U_lor_23_lpi_1_dfm_st_4 | mul_loop_mul_if_land_6_lpi_1_dfm_st_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4));
  assign mux_636_nl = MUX_s_1_2_2((nor_1228_nl), (nor_1227_nl), or_309_cse);
  assign or_1430_nl = mul_loop_mul_if_land_6_lpi_1_dfm_st_8 | mul_loop_mul_if_land_6_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_637_nl = MUX_s_1_2_2((or_1430_nl), or_tmp_1339, or_309_cse);
  assign nor_1219_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_6_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_6_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_6_lpi_1_dfm_8 | mul_loop_mul_if_land_6_lpi_1_dfm_9);
  assign nor_1220_nl = ~(nor_1221_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_6_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_6_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_6_lpi_1_dfm_8 | mul_loop_mul_if_land_6_lpi_1_dfm_9);
  assign nor_1222_nl = ~((FpMul_8U_23U_p_mant_p1_6_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_6_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_6_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_6_lpi_1_dfm_8
      | mul_loop_mul_if_land_6_lpi_1_dfm_9);
  assign mux_639_nl = MUX_s_1_2_2((nor_1222_nl), (nor_1220_nl), nor_213_cse);
  assign and_2199_nl = mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_639_nl);
  assign nor_1223_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_68_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_6_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_6_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_6_lpi_1_dfm_8
      | mul_loop_mul_if_land_6_lpi_1_dfm_9);
  assign mux_640_nl = MUX_s_1_2_2((nor_1223_nl), (and_2199_nl), nor_53_cse);
  assign mux_641_nl = MUX_s_1_2_2((mux_640_nl), (nor_1219_nl), FpMul_8U_23U_lor_23_lpi_1_dfm_6);
  assign nor_1224_nl = ~((~ or_tmp_1305) | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_6_lpi_1_dfm_11 | mul_loop_mul_if_land_6_lpi_1_dfm_10 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_6_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_6_lpi_1_dfm_9);
  assign mux_642_nl = MUX_s_1_2_2((nor_1224_nl), (mux_641_nl), or_309_cse);
  assign nor_1646_nl = ~(IsNaN_8U_23U_1_land_7_lpi_1_dfm_8 | FpMul_8U_23U_lor_24_lpi_1_dfm_st_3
      | not_tmp_1434);
  assign or_4945_nl = IsNaN_8U_23U_1_land_7_lpi_1_dfm_8 | (~(FpMul_8U_23U_lor_24_lpi_1_dfm_st_3
      | not_tmp_1434));
  assign mux_1723_nl = MUX_s_1_2_2((or_4945_nl), (nor_1646_nl), IsNaN_8U_23U_land_7_lpi_1_dfm_st_7);
  assign nor_1197_nl = ~((~((~ (mul_loop_mul_7_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_7_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 | FpMul_8U_23U_lor_24_lpi_1_dfm_6))
      | IsNaN_8U_23U_land_7_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_7_lpi_1_dfm_8
      | mul_loop_mul_if_land_7_lpi_1_dfm_9);
  assign nor_1199_nl = ~((~ FpMul_8U_23U_lor_24_lpi_1_dfm_6) | IsNaN_8U_23U_land_7_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_7_lpi_1_dfm_8 | mul_loop_mul_if_land_7_lpi_1_dfm_9);
  assign mux_656_nl = MUX_s_1_2_2((nor_1199_nl), (nor_1197_nl), mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign nor_1200_nl = ~((~ or_tmp_1382) | IsNaN_8U_23U_land_7_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_7_lpi_1_dfm_8 | mul_loop_mul_if_land_7_lpi_1_dfm_9);
  assign mux_657_nl = MUX_s_1_2_2((nor_1200_nl), (mux_656_nl), nor_53_cse);
  assign and_2194_nl = nor_225_cse & (mux_657_nl);
  assign nor_1201_nl = ~((~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8 |
      IsNaN_8U_23U_land_7_lpi_1_dfm_11 | mul_loop_mul_if_land_7_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | mul_loop_mul_if_land_7_lpi_1_dfm_st_8 | IsNaN_8U_23U_1_land_7_lpi_1_dfm_9
      | FpMul_8U_23U_lor_24_lpi_1_dfm_st_4 | (~(mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
      & or_tmp_1387 & ((~ mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs_2) | mul_loop_mul_7_FpMantRNE_48U_24U_else_and_svs_st_2))));
  assign mux_658_nl = MUX_s_1_2_2((nor_1201_nl), (and_2194_nl), or_309_cse);
  assign nor_1193_nl = ~(or_tmp_1415 | (~ main_stage_v_3));
  assign nor_1194_nl = ~(FpMul_8U_23U_lor_24_lpi_1_dfm_st_4 | mul_loop_mul_if_land_7_lpi_1_dfm_st_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4));
  assign mux_660_nl = MUX_s_1_2_2((nor_1194_nl), (nor_1193_nl), or_309_cse);
  assign or_1512_nl = mul_loop_mul_if_land_7_lpi_1_dfm_st_8 | mul_loop_mul_if_land_7_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_661_nl = MUX_s_1_2_2((or_1512_nl), or_tmp_1421, or_309_cse);
  assign nor_1185_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_7_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_7_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_7_lpi_1_dfm_8 | mul_loop_mul_if_land_7_lpi_1_dfm_9);
  assign nor_1186_nl = ~(nor_1187_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_7_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_7_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_7_lpi_1_dfm_8 | mul_loop_mul_if_land_7_lpi_1_dfm_9);
  assign nor_1188_nl = ~((FpMul_8U_23U_p_mant_p1_7_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_7_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_7_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_7_lpi_1_dfm_8
      | mul_loop_mul_if_land_7_lpi_1_dfm_9);
  assign mux_663_nl = MUX_s_1_2_2((nor_1188_nl), (nor_1186_nl), nor_229_cse);
  assign and_2193_nl = mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_663_nl);
  assign nor_1189_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_69_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_7_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_7_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_7_lpi_1_dfm_8
      | mul_loop_mul_if_land_7_lpi_1_dfm_9);
  assign mux_664_nl = MUX_s_1_2_2((nor_1189_nl), (and_2193_nl), nor_53_cse);
  assign mux_665_nl = MUX_s_1_2_2((mux_664_nl), (nor_1185_nl), FpMul_8U_23U_lor_24_lpi_1_dfm_6);
  assign nor_1190_nl = ~((~ or_tmp_1387) | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_7_lpi_1_dfm_11 | mul_loop_mul_if_land_7_lpi_1_dfm_10 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_7_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_7_lpi_1_dfm_9);
  assign mux_666_nl = MUX_s_1_2_2((nor_1190_nl), (mux_665_nl), or_309_cse);
  assign nor_1641_nl = ~(IsNaN_8U_23U_1_land_8_lpi_1_dfm_8 | FpMul_8U_23U_lor_25_lpi_1_dfm_st_3
      | not_tmp_1452);
  assign or_4942_nl = IsNaN_8U_23U_1_land_8_lpi_1_dfm_8 | (~(FpMul_8U_23U_lor_25_lpi_1_dfm_st_3
      | not_tmp_1452));
  assign mux_1728_nl = MUX_s_1_2_2((or_4942_nl), (nor_1641_nl), IsNaN_8U_23U_land_8_lpi_1_dfm_st_7);
  assign nor_1163_nl = ~((~((~ (mul_loop_mul_8_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_8_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 | FpMul_8U_23U_lor_25_lpi_1_dfm_6))
      | IsNaN_8U_23U_land_8_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_8_lpi_1_dfm_8
      | mul_loop_mul_if_land_8_lpi_1_dfm_9);
  assign nor_1165_nl = ~((~ FpMul_8U_23U_lor_25_lpi_1_dfm_6) | IsNaN_8U_23U_land_8_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_8_lpi_1_dfm_8 | mul_loop_mul_if_land_8_lpi_1_dfm_9);
  assign mux_680_nl = MUX_s_1_2_2((nor_1165_nl), (nor_1163_nl), mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign nor_1166_nl = ~((~ or_tmp_1464) | IsNaN_8U_23U_land_8_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_8_lpi_1_dfm_8 | mul_loop_mul_if_land_8_lpi_1_dfm_9);
  assign mux_681_nl = MUX_s_1_2_2((nor_1166_nl), (mux_680_nl), nor_53_cse);
  assign and_2188_nl = nor_241_cse & (mux_681_nl);
  assign nor_1167_nl = ~((~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8 |
      IsNaN_8U_23U_land_8_lpi_1_dfm_11 | mul_loop_mul_if_land_8_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | mul_loop_mul_if_land_8_lpi_1_dfm_st_8 | IsNaN_8U_23U_1_land_8_lpi_1_dfm_9
      | FpMul_8U_23U_lor_25_lpi_1_dfm_st_4 | (~(mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
      & or_tmp_1469 & ((~ mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs_2) | mul_loop_mul_8_FpMantRNE_48U_24U_else_and_svs_st_2))));
  assign mux_682_nl = MUX_s_1_2_2((nor_1167_nl), (and_2188_nl), or_309_cse);
  assign or_1587_nl = FpMul_8U_23U_lor_25_lpi_1_dfm_st_4 | mul_loop_mul_if_land_8_lpi_1_dfm_st_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_684_nl = MUX_s_1_2_2((or_1587_nl), or_tmp_397, or_309_cse);
  assign or_1592_nl = mul_loop_mul_if_land_8_lpi_1_dfm_st_8 | mul_loop_mul_if_land_8_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_685_nl = MUX_s_1_2_2((or_1592_nl), or_tmp_1501, or_309_cse);
  assign nor_1153_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_8_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_8_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_8_lpi_1_dfm_8 | mul_loop_mul_if_land_8_lpi_1_dfm_9);
  assign nor_1154_nl = ~(nor_1155_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_8_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_8_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_8_lpi_1_dfm_8 | mul_loop_mul_if_land_8_lpi_1_dfm_9);
  assign nor_1156_nl = ~((FpMul_8U_23U_p_mant_p1_8_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_8_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_8_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_8_lpi_1_dfm_8
      | mul_loop_mul_if_land_8_lpi_1_dfm_9);
  assign mux_687_nl = MUX_s_1_2_2((nor_1156_nl), (nor_1154_nl), nor_245_cse);
  assign and_2187_nl = mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_687_nl);
  assign nor_1157_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_70_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_8_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_8_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_8_lpi_1_dfm_8
      | mul_loop_mul_if_land_8_lpi_1_dfm_9);
  assign mux_688_nl = MUX_s_1_2_2((nor_1157_nl), (and_2187_nl), nor_53_cse);
  assign mux_689_nl = MUX_s_1_2_2((mux_688_nl), (nor_1153_nl), FpMul_8U_23U_lor_25_lpi_1_dfm_6);
  assign nor_1158_nl = ~((~ or_tmp_1469) | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_8_lpi_1_dfm_11 | mul_loop_mul_if_land_8_lpi_1_dfm_10 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_8_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_8_lpi_1_dfm_9);
  assign mux_690_nl = MUX_s_1_2_2((nor_1158_nl), (mux_689_nl), or_309_cse);
  assign nor_1636_nl = ~(IsNaN_8U_23U_1_land_9_lpi_1_dfm_8 | FpMul_8U_23U_lor_26_lpi_1_dfm_st_3
      | not_tmp_1470);
  assign or_4939_nl = IsNaN_8U_23U_1_land_9_lpi_1_dfm_8 | (~(FpMul_8U_23U_lor_26_lpi_1_dfm_st_3
      | not_tmp_1470));
  assign mux_1733_nl = MUX_s_1_2_2((or_4939_nl), (nor_1636_nl), IsNaN_8U_23U_land_9_lpi_1_dfm_st_7);
  assign nor_1131_nl = ~((~((~ (mul_loop_mul_9_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_9_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 | FpMul_8U_23U_lor_26_lpi_1_dfm_6))
      | IsNaN_8U_23U_land_9_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_9_lpi_1_dfm_8
      | mul_loop_mul_if_land_9_lpi_1_dfm_9);
  assign nor_1133_nl = ~((~ FpMul_8U_23U_lor_26_lpi_1_dfm_6) | IsNaN_8U_23U_land_9_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_9_lpi_1_dfm_8 | mul_loop_mul_if_land_9_lpi_1_dfm_9);
  assign mux_704_nl = MUX_s_1_2_2((nor_1133_nl), (nor_1131_nl), mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign nor_1134_nl = ~((~ or_tmp_1544) | IsNaN_8U_23U_land_9_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_9_lpi_1_dfm_8 | mul_loop_mul_if_land_9_lpi_1_dfm_9);
  assign mux_705_nl = MUX_s_1_2_2((nor_1134_nl), (mux_704_nl), nor_53_cse);
  assign and_2182_nl = nor_257_cse & (mux_705_nl);
  assign nor_1135_nl = ~((~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8 |
      IsNaN_8U_23U_land_9_lpi_1_dfm_11 | mul_loop_mul_if_land_9_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | mul_loop_mul_if_land_9_lpi_1_dfm_st_8 | IsNaN_8U_23U_1_land_9_lpi_1_dfm_9
      | FpMul_8U_23U_lor_26_lpi_1_dfm_st_4 | (~(mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
      & or_tmp_1549 & ((~ mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs_2) | mul_loop_mul_9_FpMantRNE_48U_24U_else_and_svs_st_2))));
  assign mux_706_nl = MUX_s_1_2_2((nor_1135_nl), (and_2182_nl), or_309_cse);
  assign or_1667_nl = FpMul_8U_23U_lor_26_lpi_1_dfm_st_4 | mul_loop_mul_if_land_9_lpi_1_dfm_st_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_708_nl = MUX_s_1_2_2((or_1667_nl), or_tmp_425, or_309_cse);
  assign or_1672_nl = mul_loop_mul_if_land_9_lpi_1_dfm_st_8 | mul_loop_mul_if_land_9_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_709_nl = MUX_s_1_2_2((or_1672_nl), or_tmp_1581, or_309_cse);
  assign nor_1121_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_9_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_9_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_9_lpi_1_dfm_8 | mul_loop_mul_if_land_9_lpi_1_dfm_9);
  assign nor_1122_nl = ~(nor_1123_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_9_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_9_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_9_lpi_1_dfm_8 | mul_loop_mul_if_land_9_lpi_1_dfm_9);
  assign nor_1124_nl = ~((FpMul_8U_23U_p_mant_p1_9_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_9_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_9_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_9_lpi_1_dfm_8
      | mul_loop_mul_if_land_9_lpi_1_dfm_9);
  assign mux_711_nl = MUX_s_1_2_2((nor_1124_nl), (nor_1122_nl), nor_261_cse);
  assign and_2181_nl = mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_711_nl);
  assign nor_1125_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_71_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_9_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_9_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_9_lpi_1_dfm_8
      | mul_loop_mul_if_land_9_lpi_1_dfm_9);
  assign mux_712_nl = MUX_s_1_2_2((nor_1125_nl), (and_2181_nl), nor_53_cse);
  assign mux_713_nl = MUX_s_1_2_2((mux_712_nl), (nor_1121_nl), FpMul_8U_23U_lor_26_lpi_1_dfm_6);
  assign nor_1126_nl = ~((~ or_tmp_1549) | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_9_lpi_1_dfm_11 | mul_loop_mul_if_land_9_lpi_1_dfm_10 |
      io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_9_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_9_lpi_1_dfm_9);
  assign mux_714_nl = MUX_s_1_2_2((nor_1126_nl), (mux_713_nl), or_309_cse);
  assign nor_1631_nl = ~(IsNaN_8U_23U_1_land_10_lpi_1_dfm_8 | FpMul_8U_23U_lor_27_lpi_1_dfm_st_3
      | not_tmp_1488);
  assign or_4936_nl = IsNaN_8U_23U_1_land_10_lpi_1_dfm_8 | (~(FpMul_8U_23U_lor_27_lpi_1_dfm_st_3
      | not_tmp_1488));
  assign mux_1738_nl = MUX_s_1_2_2((or_4936_nl), (nor_1631_nl), IsNaN_8U_23U_land_10_lpi_1_dfm_st_7);
  assign nor_1098_nl = ~((~((~ (mul_loop_mul_10_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_10_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 | FpMul_8U_23U_lor_27_lpi_1_dfm_6))
      | IsNaN_8U_23U_land_10_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_10_lpi_1_dfm_8
      | mul_loop_mul_if_land_10_lpi_1_dfm_9);
  assign nor_1100_nl = ~((~ FpMul_8U_23U_lor_27_lpi_1_dfm_6) | IsNaN_8U_23U_land_10_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_10_lpi_1_dfm_8 | mul_loop_mul_if_land_10_lpi_1_dfm_9);
  assign mux_728_nl = MUX_s_1_2_2((nor_1100_nl), (nor_1098_nl), mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign nor_1101_nl = ~((~ or_tmp_1624) | IsNaN_8U_23U_land_10_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_10_lpi_1_dfm_8 | mul_loop_mul_if_land_10_lpi_1_dfm_9);
  assign mux_729_nl = MUX_s_1_2_2((nor_1101_nl), (mux_728_nl), nor_53_cse);
  assign and_2175_nl = nor_273_cse & (mux_729_nl);
  assign and_2176_nl = or_tmp_1629 & (~(nor_1103_cse | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_10_lpi_1_dfm_11 | mul_loop_mul_if_land_10_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_10_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_10_lpi_1_dfm_9 | FpMul_8U_23U_lor_27_lpi_1_dfm_st_4 |
      (~ mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4)));
  assign mux_730_nl = MUX_s_1_2_2((and_2176_nl), (and_2175_nl), or_309_cse);
  assign or_1747_nl = FpMul_8U_23U_lor_27_lpi_1_dfm_st_4 | mul_loop_mul_if_land_10_lpi_1_dfm_st_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_732_nl = MUX_s_1_2_2((or_1747_nl), or_tmp_454, or_309_cse);
  assign or_1752_nl = mul_loop_mul_if_land_10_lpi_1_dfm_st_8 | mul_loop_mul_if_land_10_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_733_nl = MUX_s_1_2_2((or_1752_nl), or_tmp_1661, or_309_cse);
  assign nor_1088_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_10_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_10_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_10_lpi_1_dfm_8 | mul_loop_mul_if_land_10_lpi_1_dfm_9);
  assign nor_1089_nl = ~(nor_1090_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_10_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_10_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_10_lpi_1_dfm_8 | mul_loop_mul_if_land_10_lpi_1_dfm_9);
  assign nor_1091_nl = ~((FpMul_8U_23U_p_mant_p1_10_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_10_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_10_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_10_lpi_1_dfm_8
      | mul_loop_mul_if_land_10_lpi_1_dfm_9);
  assign mux_735_nl = MUX_s_1_2_2((nor_1091_nl), (nor_1089_nl), nor_277_cse);
  assign and_2174_nl = mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_735_nl);
  assign nor_1092_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_72_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_10_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_10_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_10_lpi_1_dfm_8
      | mul_loop_mul_if_land_10_lpi_1_dfm_9);
  assign mux_736_nl = MUX_s_1_2_2((nor_1092_nl), (and_2174_nl), nor_53_cse);
  assign mux_737_nl = MUX_s_1_2_2((mux_736_nl), (nor_1088_nl), FpMul_8U_23U_lor_27_lpi_1_dfm_6);
  assign nor_1093_nl = ~((~ or_tmp_1629) | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_10_lpi_1_dfm_11 | mul_loop_mul_if_land_10_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_10_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_10_lpi_1_dfm_9);
  assign mux_738_nl = MUX_s_1_2_2((nor_1093_nl), (mux_737_nl), or_309_cse);
  assign nor_1627_nl = ~(IsNaN_8U_23U_1_land_11_lpi_1_dfm_8 | FpMul_8U_23U_lor_28_lpi_1_dfm_st_3
      | not_tmp_1506);
  assign or_4935_nl = IsNaN_8U_23U_1_land_11_lpi_1_dfm_8 | (~(FpMul_8U_23U_lor_28_lpi_1_dfm_st_3
      | not_tmp_1506));
  assign mux_1745_nl = MUX_s_1_2_2((or_4935_nl), (nor_1627_nl), IsNaN_8U_23U_land_11_lpi_1_dfm_st_7);
  assign nor_1065_nl = ~((~((~ (mul_loop_mul_11_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 | FpMul_8U_23U_lor_28_lpi_1_dfm_6))
      | IsNaN_8U_23U_land_11_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_11_lpi_1_dfm_8
      | mul_loop_mul_if_land_11_lpi_1_dfm_9);
  assign nor_1067_nl = ~((~ FpMul_8U_23U_lor_28_lpi_1_dfm_6) | IsNaN_8U_23U_land_11_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_11_lpi_1_dfm_8 | mul_loop_mul_if_land_11_lpi_1_dfm_9);
  assign mux_752_nl = MUX_s_1_2_2((nor_1067_nl), (nor_1065_nl), mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign nor_1068_nl = ~((~ or_tmp_1703) | IsNaN_8U_23U_land_11_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_11_lpi_1_dfm_8 | mul_loop_mul_if_land_11_lpi_1_dfm_9);
  assign mux_753_nl = MUX_s_1_2_2((nor_1068_nl), (mux_752_nl), nor_53_cse);
  assign and_2166_nl = nor_289_cse & (mux_753_nl);
  assign and_2167_nl = or_tmp_1709 & (~(nor_1070_cse | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_11_lpi_1_dfm_11 | mul_loop_mul_if_land_11_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_11_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_11_lpi_1_dfm_9 | FpMul_8U_23U_lor_28_lpi_1_dfm_st_4 |
      (~ mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4)));
  assign mux_754_nl = MUX_s_1_2_2((and_2167_nl), (and_2166_nl), or_309_cse);
  assign or_1830_nl = FpMul_8U_23U_lor_28_lpi_1_dfm_st_4 | (~ reg_chn_mul_out_rsci_ld_core_psct_cse)
      | chn_mul_out_rsci_bawt | mul_loop_mul_if_land_11_lpi_1_dfm_st_8 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | (~ main_stage_v_4);
  assign mux_758_nl = MUX_s_1_2_2(mux_tmp_748, or_tmp_1736, FpMul_8U_23U_lor_28_lpi_1_dfm_st_4);
  assign mux_759_nl = MUX_s_1_2_2((mux_758_nl), (or_1830_nl), FpMul_8U_23U_lor_28_lpi_1_dfm_st_3);
  assign or_1835_nl = mul_loop_mul_if_land_11_lpi_1_dfm_st_8 | mul_loop_mul_if_land_11_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_760_nl = MUX_s_1_2_2((or_1835_nl), or_tmp_1744, or_309_cse);
  assign nor_1057_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_11_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_11_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_11_lpi_1_dfm_8 | mul_loop_mul_if_land_11_lpi_1_dfm_9);
  assign nor_1058_nl = ~(nor_1059_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_11_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_11_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_11_lpi_1_dfm_8 | mul_loop_mul_if_land_11_lpi_1_dfm_9);
  assign nor_1060_nl = ~((FpMul_8U_23U_p_mant_p1_11_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_11_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_11_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_11_lpi_1_dfm_8
      | mul_loop_mul_if_land_11_lpi_1_dfm_9);
  assign mux_762_nl = MUX_s_1_2_2((nor_1060_nl), (nor_1058_nl), nor_283_cse);
  assign and_2165_nl = mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_762_nl);
  assign nor_1061_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_73_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_11_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_11_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_11_lpi_1_dfm_8
      | mul_loop_mul_if_land_11_lpi_1_dfm_9);
  assign mux_763_nl = MUX_s_1_2_2((nor_1061_nl), (and_2165_nl), nor_53_cse);
  assign mux_764_nl = MUX_s_1_2_2((mux_763_nl), (nor_1057_nl), FpMul_8U_23U_lor_28_lpi_1_dfm_6);
  assign nor_1062_nl = ~((~ or_tmp_1709) | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_11_lpi_1_dfm_11 | mul_loop_mul_if_land_11_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_11_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_11_lpi_1_dfm_9);
  assign mux_765_nl = MUX_s_1_2_2((nor_1062_nl), (mux_764_nl), or_309_cse);
  assign nor_1622_nl = ~(IsNaN_8U_23U_1_land_12_lpi_1_dfm_8 | FpMul_8U_23U_lor_29_lpi_1_dfm_st_3
      | not_tmp_1524);
  assign or_4932_nl = IsNaN_8U_23U_1_land_12_lpi_1_dfm_8 | (~(FpMul_8U_23U_lor_29_lpi_1_dfm_st_3
      | not_tmp_1524));
  assign mux_1750_nl = MUX_s_1_2_2((or_4932_nl), (nor_1622_nl), IsNaN_8U_23U_land_12_lpi_1_dfm_st_7);
  assign nor_1032_nl = ~((~((~ (mul_loop_mul_12_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_12_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 | FpMul_8U_23U_lor_29_lpi_1_dfm_6))
      | IsNaN_8U_23U_land_12_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_12_lpi_1_dfm_8
      | mul_loop_mul_if_land_12_lpi_1_dfm_9);
  assign nor_1034_nl = ~((~ FpMul_8U_23U_lor_29_lpi_1_dfm_6) | IsNaN_8U_23U_land_12_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_12_lpi_1_dfm_8 | mul_loop_mul_if_land_12_lpi_1_dfm_9);
  assign mux_779_nl = MUX_s_1_2_2((nor_1034_nl), (nor_1032_nl), mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign nor_1035_nl = ~((~ or_tmp_1782) | IsNaN_8U_23U_land_12_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_12_lpi_1_dfm_8 | mul_loop_mul_if_land_12_lpi_1_dfm_9);
  assign mux_780_nl = MUX_s_1_2_2((nor_1035_nl), (mux_779_nl), nor_53_cse);
  assign and_2160_nl = nor_305_cse & (mux_780_nl);
  assign and_2161_nl = or_tmp_1786 & (~(nor_1037_cse | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_12_lpi_1_dfm_11 | mul_loop_mul_if_land_12_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_12_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_12_lpi_1_dfm_9 | FpMul_8U_23U_lor_29_lpi_1_dfm_st_4 |
      (~ mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4)));
  assign mux_781_nl = MUX_s_1_2_2((and_2161_nl), (and_2160_nl), or_309_cse);
  assign or_1905_nl = (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt
      | FpMul_8U_23U_lor_29_lpi_1_dfm_st_4 | mul_loop_mul_if_land_12_lpi_1_dfm_st_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign or_1908_nl = FpMul_8U_23U_lor_29_lpi_1_dfm_st_4 | mul_loop_mul_if_land_12_lpi_1_dfm_st_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_784_nl = MUX_s_1_2_2((or_1908_nl), or_tmp_509, or_309_cse);
  assign mux_785_nl = MUX_s_1_2_2((mux_784_nl), (or_1905_nl), FpMul_8U_23U_lor_29_lpi_1_dfm_st_3);
  assign or_1913_nl = mul_loop_mul_if_land_12_lpi_1_dfm_st_8 | mul_loop_mul_if_land_12_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_786_nl = MUX_s_1_2_2((or_1913_nl), or_tmp_1822, or_309_cse);
  assign nor_1024_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_12_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_12_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_12_lpi_1_dfm_8 | mul_loop_mul_if_land_12_lpi_1_dfm_9);
  assign nor_1025_nl = ~(nor_1026_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_12_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_12_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_12_lpi_1_dfm_8 | mul_loop_mul_if_land_12_lpi_1_dfm_9);
  assign nor_1027_nl = ~((FpMul_8U_23U_p_mant_p1_12_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_12_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_12_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_12_lpi_1_dfm_8
      | mul_loop_mul_if_land_12_lpi_1_dfm_9);
  assign mux_788_nl = MUX_s_1_2_2((nor_1027_nl), (nor_1025_nl), nor_309_cse);
  assign and_2159_nl = mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_788_nl);
  assign nor_1028_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_74_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_12_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_12_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_12_lpi_1_dfm_8
      | mul_loop_mul_if_land_12_lpi_1_dfm_9);
  assign mux_789_nl = MUX_s_1_2_2((nor_1028_nl), (and_2159_nl), nor_53_cse);
  assign mux_790_nl = MUX_s_1_2_2((mux_789_nl), (nor_1024_nl), FpMul_8U_23U_lor_29_lpi_1_dfm_6);
  assign nor_1029_nl = ~((~ or_tmp_1786) | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_12_lpi_1_dfm_11 | mul_loop_mul_if_land_12_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_12_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_12_lpi_1_dfm_9);
  assign mux_791_nl = MUX_s_1_2_2((nor_1029_nl), (mux_790_nl), or_309_cse);
  assign nor_1617_nl = ~(IsNaN_8U_23U_1_land_13_lpi_1_dfm_8 | FpMul_8U_23U_lor_30_lpi_1_dfm_st_3
      | not_tmp_1542);
  assign or_4929_nl = IsNaN_8U_23U_1_land_13_lpi_1_dfm_8 | (~(FpMul_8U_23U_lor_30_lpi_1_dfm_st_3
      | not_tmp_1542));
  assign mux_1755_nl = MUX_s_1_2_2((or_4929_nl), (nor_1617_nl), IsNaN_8U_23U_land_13_lpi_1_dfm_st_7);
  assign nor_999_nl = ~((~((~ (mul_loop_mul_13_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_13_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 | FpMul_8U_23U_lor_30_lpi_1_dfm_6))
      | IsNaN_8U_23U_land_13_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_13_lpi_1_dfm_8
      | mul_loop_mul_if_land_13_lpi_1_dfm_9);
  assign nor_1001_nl = ~((~ FpMul_8U_23U_lor_30_lpi_1_dfm_6) | IsNaN_8U_23U_land_13_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_13_lpi_1_dfm_8 | mul_loop_mul_if_land_13_lpi_1_dfm_9);
  assign mux_806_nl = MUX_s_1_2_2((nor_1001_nl), (nor_999_nl), mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign nor_1002_nl = ~((~ or_tmp_1865) | IsNaN_8U_23U_land_13_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_13_lpi_1_dfm_8 | mul_loop_mul_if_land_13_lpi_1_dfm_9);
  assign mux_807_nl = MUX_s_1_2_2((nor_1002_nl), (mux_806_nl), nor_53_cse);
  assign and_2154_nl = nor_321_cse & (mux_807_nl);
  assign and_2155_nl = or_tmp_1869 & (~(nor_1004_cse | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_13_lpi_1_dfm_11 | mul_loop_mul_if_land_13_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_13_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_13_lpi_1_dfm_9 | FpMul_8U_23U_lor_30_lpi_1_dfm_st_4 |
      (~ mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4)));
  assign mux_808_nl = MUX_s_1_2_2((and_2155_nl), (and_2154_nl), or_309_cse);
  assign or_1988_nl = (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt
      | FpMul_8U_23U_lor_30_lpi_1_dfm_st_4 | mul_loop_mul_if_land_13_lpi_1_dfm_st_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign or_1991_nl = FpMul_8U_23U_lor_30_lpi_1_dfm_st_4 | mul_loop_mul_if_land_13_lpi_1_dfm_st_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_811_nl = MUX_s_1_2_2((or_1991_nl), or_tmp_532, or_309_cse);
  assign mux_812_nl = MUX_s_1_2_2((mux_811_nl), (or_1988_nl), FpMul_8U_23U_lor_30_lpi_1_dfm_st_3);
  assign or_1996_nl = mul_loop_mul_if_land_13_lpi_1_dfm_st_8 | mul_loop_mul_if_land_13_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_813_nl = MUX_s_1_2_2((or_1996_nl), or_tmp_1905, or_309_cse);
  assign nor_991_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_13_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_13_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_13_lpi_1_dfm_8 | mul_loop_mul_if_land_13_lpi_1_dfm_9);
  assign nor_992_nl = ~(nor_993_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_13_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_13_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_13_lpi_1_dfm_8 | mul_loop_mul_if_land_13_lpi_1_dfm_9);
  assign nor_994_nl = ~((FpMul_8U_23U_p_mant_p1_13_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_13_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_13_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_13_lpi_1_dfm_8
      | mul_loop_mul_if_land_13_lpi_1_dfm_9);
  assign mux_815_nl = MUX_s_1_2_2((nor_994_nl), (nor_992_nl), nor_325_cse);
  assign and_2153_nl = mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_815_nl);
  assign nor_995_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_75_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_13_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_13_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_13_lpi_1_dfm_8
      | mul_loop_mul_if_land_13_lpi_1_dfm_9);
  assign mux_816_nl = MUX_s_1_2_2((nor_995_nl), (and_2153_nl), nor_53_cse);
  assign mux_817_nl = MUX_s_1_2_2((mux_816_nl), (nor_991_nl), FpMul_8U_23U_lor_30_lpi_1_dfm_6);
  assign nor_996_nl = ~((~ or_tmp_1869) | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_13_lpi_1_dfm_11 | mul_loop_mul_if_land_13_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_13_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_13_lpi_1_dfm_9);
  assign mux_818_nl = MUX_s_1_2_2((nor_996_nl), (mux_817_nl), or_309_cse);
  assign nor_1612_nl = ~(IsNaN_8U_23U_1_land_14_lpi_1_dfm_8 | (~ mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_31_lpi_1_dfm_st_3 | (~ mux_1758_cse));
  assign or_4928_nl = IsNaN_8U_23U_1_land_14_lpi_1_dfm_8 | (~((~ mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_31_lpi_1_dfm_st_3 | (~ mux_1758_cse)));
  assign mux_1762_nl = MUX_s_1_2_2((or_4928_nl), (nor_1612_nl), IsNaN_8U_23U_land_14_lpi_1_dfm_st_7);
  assign nor_967_nl = ~((~((~ (mul_loop_mul_14_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 | FpMul_8U_23U_lor_31_lpi_1_dfm_6))
      | IsNaN_8U_23U_land_14_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_14_lpi_1_dfm_8
      | mul_loop_mul_if_land_14_lpi_1_dfm_9);
  assign nor_969_nl = ~((~ FpMul_8U_23U_lor_31_lpi_1_dfm_6) | IsNaN_8U_23U_land_14_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_14_lpi_1_dfm_8 | mul_loop_mul_if_land_14_lpi_1_dfm_9);
  assign mux_833_nl = MUX_s_1_2_2((nor_969_nl), (nor_967_nl), mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign nor_970_nl = ~((~ or_tmp_1947) | IsNaN_8U_23U_land_14_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_14_lpi_1_dfm_8 | mul_loop_mul_if_land_14_lpi_1_dfm_9);
  assign mux_834_nl = MUX_s_1_2_2((nor_970_nl), (mux_833_nl), nor_53_cse);
  assign and_2149_nl = nor_336_cse & (mux_834_nl);
  assign and_2150_nl = or_tmp_1957 & (~(nor_972_cse | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_14_lpi_1_dfm_11 | mul_loop_mul_if_land_14_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_14_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_14_lpi_1_dfm_9 | FpMul_8U_23U_lor_31_lpi_1_dfm_st_4 |
      (~ mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4)));
  assign mux_835_nl = MUX_s_1_2_2((and_2150_nl), (and_2149_nl), or_309_cse);
  assign nor_963_nl = ~(or_tmp_1985 | (~ main_stage_v_3));
  assign nor_964_nl = ~(FpMul_8U_23U_lor_31_lpi_1_dfm_st_4 | mul_loop_mul_if_land_14_lpi_1_dfm_st_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4));
  assign mux_837_nl = MUX_s_1_2_2((nor_964_nl), (nor_963_nl), or_309_cse);
  assign or_2082_nl = mul_loop_mul_if_land_14_lpi_1_dfm_st_8 | mul_loop_mul_if_land_14_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_838_nl = MUX_s_1_2_2((or_2082_nl), or_tmp_1991, or_309_cse);
  assign nor_955_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_14_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_14_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_14_lpi_1_dfm_8 | mul_loop_mul_if_land_14_lpi_1_dfm_9);
  assign nor_956_nl = ~(nor_332_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_14_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_14_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_14_lpi_1_dfm_8 | mul_loop_mul_if_land_14_lpi_1_dfm_9);
  assign nor_958_nl = ~((FpMul_8U_23U_p_mant_p1_14_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_14_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_14_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_14_lpi_1_dfm_8
      | mul_loop_mul_if_land_14_lpi_1_dfm_9);
  assign mux_840_nl = MUX_s_1_2_2((nor_958_nl), (nor_956_nl), nor_340_cse);
  assign and_2148_nl = mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_840_nl);
  assign nor_959_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_76_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_14_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_14_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_14_lpi_1_dfm_8
      | mul_loop_mul_if_land_14_lpi_1_dfm_9);
  assign mux_841_nl = MUX_s_1_2_2((nor_959_nl), (and_2148_nl), nor_53_cse);
  assign mux_842_nl = MUX_s_1_2_2((mux_841_nl), (nor_955_nl), FpMul_8U_23U_lor_31_lpi_1_dfm_6);
  assign nor_960_nl = ~((~ or_tmp_1957) | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_14_lpi_1_dfm_11 | mul_loop_mul_if_land_14_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_14_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_14_lpi_1_dfm_9);
  assign mux_843_nl = MUX_s_1_2_2((nor_960_nl), (mux_842_nl), or_309_cse);
  assign nor_1607_nl = ~(IsNaN_8U_23U_1_land_15_lpi_1_dfm_8 | FpMul_8U_23U_lor_32_lpi_1_dfm_st_3
      | not_tmp_1578);
  assign or_4925_nl = IsNaN_8U_23U_1_land_15_lpi_1_dfm_8 | (~(FpMul_8U_23U_lor_32_lpi_1_dfm_st_3
      | not_tmp_1578));
  assign mux_1767_nl = MUX_s_1_2_2((or_4925_nl), (nor_1607_nl), IsNaN_8U_23U_land_15_lpi_1_dfm_st_7);
  assign nor_930_nl = ~((~((~ (mul_loop_mul_15_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_15_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 | FpMul_8U_23U_lor_32_lpi_1_dfm_6))
      | IsNaN_8U_23U_land_15_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_15_lpi_1_dfm_8
      | mul_loop_mul_if_land_15_lpi_1_dfm_9);
  assign nor_932_nl = ~((~ FpMul_8U_23U_lor_32_lpi_1_dfm_6) | IsNaN_8U_23U_land_15_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_15_lpi_1_dfm_8 | mul_loop_mul_if_land_15_lpi_1_dfm_9);
  assign mux_858_nl = MUX_s_1_2_2((nor_932_nl), (nor_930_nl), mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign nor_933_nl = ~((~ or_tmp_2032) | IsNaN_8U_23U_land_15_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_15_lpi_1_dfm_8 | mul_loop_mul_if_land_15_lpi_1_dfm_9);
  assign mux_859_nl = MUX_s_1_2_2((nor_933_nl), (mux_858_nl), nor_53_cse);
  assign and_2143_nl = nor_352_cse & (mux_859_nl);
  assign and_2144_nl = or_tmp_2036 & (~(nor_935_cse | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_15_lpi_1_dfm_11 | mul_loop_mul_if_land_15_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_15_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_15_lpi_1_dfm_9 | FpMul_8U_23U_lor_32_lpi_1_dfm_st_4 |
      (~ mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4)));
  assign mux_860_nl = MUX_s_1_2_2((and_2144_nl), (and_2143_nl), or_309_cse);
  assign nor_926_nl = ~(or_tmp_2065 | (~ main_stage_v_3));
  assign nor_927_nl = ~(FpMul_8U_23U_lor_32_lpi_1_dfm_st_4 | mul_loop_mul_if_land_15_lpi_1_dfm_st_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4));
  assign mux_862_nl = MUX_s_1_2_2((nor_927_nl), (nor_926_nl), or_309_cse);
  assign or_2162_nl = mul_loop_mul_if_land_15_lpi_1_dfm_st_8 | mul_loop_mul_if_land_15_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_863_nl = MUX_s_1_2_2((or_2162_nl), or_tmp_2071, or_309_cse);
  assign nor_918_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_15_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_15_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_15_lpi_1_dfm_8 | mul_loop_mul_if_land_15_lpi_1_dfm_9);
  assign nor_919_nl = ~(nor_920_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_15_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_15_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_15_lpi_1_dfm_8 | mul_loop_mul_if_land_15_lpi_1_dfm_9);
  assign nor_921_nl = ~((FpMul_8U_23U_p_mant_p1_15_sva[47]) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_15_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_15_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_15_lpi_1_dfm_8
      | mul_loop_mul_if_land_15_lpi_1_dfm_9);
  assign mux_865_nl = MUX_s_1_2_2((nor_921_nl), (nor_919_nl), nor_356_cse);
  assign and_2142_nl = mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_865_nl);
  assign nor_922_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_77_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_15_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_15_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_15_lpi_1_dfm_8
      | mul_loop_mul_if_land_15_lpi_1_dfm_9);
  assign mux_866_nl = MUX_s_1_2_2((nor_922_nl), (and_2142_nl), nor_53_cse);
  assign mux_867_nl = MUX_s_1_2_2((mux_866_nl), (nor_918_nl), FpMul_8U_23U_lor_32_lpi_1_dfm_6);
  assign nor_923_nl = ~((~ or_tmp_2036) | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_15_lpi_1_dfm_11 | mul_loop_mul_if_land_15_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | mul_loop_mul_if_land_15_lpi_1_dfm_st_8
      | IsNaN_8U_23U_1_land_15_lpi_1_dfm_9);
  assign mux_868_nl = MUX_s_1_2_2((nor_923_nl), (mux_867_nl), or_309_cse);
  assign nor_1602_nl = ~(IsNaN_8U_23U_1_land_lpi_1_dfm_8 | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3
      | not_tmp_1596);
  assign or_4922_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_8 | (~(FpMul_8U_23U_lor_1_lpi_1_dfm_st_3
      | not_tmp_1596));
  assign mux_1772_nl = MUX_s_1_2_2((or_4922_nl), (nor_1602_nl), IsNaN_8U_23U_land_lpi_1_dfm_st_7);
  assign nor_893_nl = ~((~((~ (mul_loop_mul_16_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_16_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7 | FpMul_8U_23U_lor_1_lpi_1_dfm_6))
      | IsNaN_8U_23U_land_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_lpi_1_dfm_8
      | mul_loop_mul_if_land_lpi_1_dfm_9);
  assign nor_895_nl = ~((~ FpMul_8U_23U_lor_1_lpi_1_dfm_6) | IsNaN_8U_23U_land_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_lpi_1_dfm_8 | mul_loop_mul_if_land_lpi_1_dfm_9);
  assign mux_883_nl = MUX_s_1_2_2((nor_895_nl), (nor_893_nl), mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign nor_896_nl = ~((~ or_tmp_2114) | IsNaN_8U_23U_land_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_lpi_1_dfm_8 | mul_loop_mul_if_land_lpi_1_dfm_9);
  assign mux_884_nl = MUX_s_1_2_2((nor_896_nl), (mux_883_nl), nor_53_cse);
  assign and_2137_nl = nor_368_cse & (mux_884_nl);
  assign and_2138_nl = or_tmp_2118 & (~(nor_898_cse | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_lpi_1_dfm_11 | mul_loop_mul_if_land_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | mul_loop_mul_if_land_lpi_1_dfm_st_8 | IsNaN_8U_23U_1_land_lpi_1_dfm_9 | FpMul_8U_23U_lor_1_lpi_1_dfm_st_4
      | (~ mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4)));
  assign mux_885_nl = MUX_s_1_2_2((and_2138_nl), (and_2137_nl), or_309_cse);
  assign or_2237_nl = FpMul_8U_23U_lor_1_lpi_1_dfm_st_4 | mul_loop_mul_if_land_lpi_1_dfm_st_8
      | io_read_cfg_mul_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign mux_887_nl = MUX_s_1_2_2((or_2237_nl), or_tmp_598, or_309_cse);
  assign or_2242_nl = mul_loop_mul_if_land_lpi_1_dfm_st_8 | mul_loop_mul_if_land_lpi_1_dfm_10
      | io_read_cfg_mul_bypass_rsc_svs_8 | io_read_cfg_mul_bypass_rsc_svs_st_7 |
      (~ main_stage_v_4);
  assign mux_888_nl = MUX_s_1_2_2((or_2242_nl), or_tmp_2151, or_309_cse);
  assign nor_883_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_lpi_1_dfm_8 | mul_loop_mul_if_land_lpi_1_dfm_9);
  assign nor_884_nl = ~(nor_885_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_lpi_1_dfm_8 | mul_loop_mul_if_land_lpi_1_dfm_9);
  assign nor_886_nl = ~((FpMul_8U_23U_p_mant_p1_sva[47]) | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_lpi_1_dfm_st_7 | IsNaN_8U_23U_land_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7
      | IsNaN_8U_23U_1_land_lpi_1_dfm_8 | mul_loop_mul_if_land_lpi_1_dfm_9);
  assign mux_890_nl = MUX_s_1_2_2((nor_886_nl), (nor_884_nl), nor_372_cse);
  assign and_2136_nl = mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_890_nl);
  assign nor_887_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_78_itm) | (~ main_stage_v_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_lpi_1_dfm_st_7
      | IsNaN_8U_23U_land_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_7 | IsNaN_8U_23U_1_land_lpi_1_dfm_8
      | mul_loop_mul_if_land_lpi_1_dfm_9);
  assign mux_891_nl = MUX_s_1_2_2((nor_887_nl), (and_2136_nl), nor_53_cse);
  assign mux_892_nl = MUX_s_1_2_2((mux_891_nl), (nor_883_nl), FpMul_8U_23U_lor_1_lpi_1_dfm_6);
  assign nor_888_nl = ~((~ or_tmp_2118) | (~ main_stage_v_4) | io_read_cfg_mul_bypass_rsc_svs_8
      | IsNaN_8U_23U_land_lpi_1_dfm_11 | mul_loop_mul_if_land_lpi_1_dfm_10 | io_read_cfg_mul_bypass_rsc_svs_st_7
      | mul_loop_mul_if_land_lpi_1_dfm_st_8 | IsNaN_8U_23U_1_land_lpi_1_dfm_9);
  assign mux_893_nl = MUX_s_1_2_2((nor_888_nl), (mux_892_nl), or_309_cse);
  assign or_2282_nl = nor_872_cse | (~ mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_18_lpi_1_dfm_st_3 | (mul_loop_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47])
      | mul_loop_mul_if_land_1_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign nor_873_nl = ~(nor_872_cse | (~ mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_18_lpi_1_dfm_st_3 | (~ (mul_loop_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_if_land_1_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign mux_901_nl = MUX_s_1_2_2((nor_873_nl), (or_2282_nl), mul_loop_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm);
  assign mux_902_nl = MUX_s_1_2_2((mux_901_nl), mul_loop_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      or_90_cse);
  assign mux_903_nl = MUX_s_1_2_2((~ (FpMul_8U_23U_p_mant_p1_1_sva[47])), or_cse,
      nor_133_cse);
  assign and_323_nl = mul_loop_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_903_nl);
  assign mux_904_nl = MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_itm, (and_323_nl),
      or_309_cse);
  assign or_2286_nl = (cfg_precision!=2'b10) | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_1_lpi_1_dfm_st_7;
  assign mux_905_nl = MUX_s_1_2_2((mux_904_nl), FpMul_8U_23U_FpMul_8U_23U_and_itm,
      or_2286_nl);
  assign or_2293_nl = nor_872_cse | (~ mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_19_lpi_1_dfm_st_3 | (mul_loop_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47])
      | mul_loop_mul_if_land_2_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign nor_870_nl = ~(nor_872_cse | (~ mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_19_lpi_1_dfm_st_3 | (~ (mul_loop_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_if_land_2_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign mux_906_nl = MUX_s_1_2_2((nor_870_nl), (or_2293_nl), mul_loop_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm);
  assign mux_907_nl = MUX_s_1_2_2((mux_906_nl), mul_loop_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      or_90_cse);
  assign mux_908_nl = MUX_s_1_2_2((~ (FpMul_8U_23U_p_mant_p1_2_sva[47])), or_4962_cse,
      nor_149_cse);
  assign and_324_nl = mul_loop_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_908_nl);
  assign mux_909_nl = MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_64_itm, (and_324_nl),
      or_309_cse);
  assign or_2297_nl = (cfg_precision!=2'b10) | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_2_lpi_1_dfm_st_7;
  assign mux_910_nl = MUX_s_1_2_2((mux_909_nl), FpMul_8U_23U_FpMul_8U_23U_and_64_itm,
      or_2297_nl);
  assign or_2304_nl = nor_872_cse | (~ mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_20_lpi_1_dfm_st_3 | (mul_loop_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47])
      | mul_loop_mul_if_land_3_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign nor_867_nl = ~(nor_872_cse | (~ mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_20_lpi_1_dfm_st_3 | (~ (mul_loop_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_if_land_3_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign mux_911_nl = MUX_s_1_2_2((nor_867_nl), (or_2304_nl), mul_loop_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm);
  assign mux_912_nl = MUX_s_1_2_2((mux_911_nl), mul_loop_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      or_90_cse);
  assign mux_913_nl = MUX_s_1_2_2((~ (FpMul_8U_23U_p_mant_p1_3_sva[47])), or_4959_cse,
      nor_165_cse);
  assign and_325_nl = mul_loop_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_913_nl);
  assign mux_914_nl = MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_65_itm, (and_325_nl),
      or_309_cse);
  assign or_2308_nl = (cfg_precision!=2'b10) | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_3_lpi_1_dfm_st_7;
  assign mux_915_nl = MUX_s_1_2_2((mux_914_nl), FpMul_8U_23U_FpMul_8U_23U_and_65_itm,
      or_2308_nl);
  assign or_2317_nl = (~ mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_21_lpi_1_dfm_st_3 | (mul_loop_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47])
      | or_tmp_2227;
  assign nor_865_nl = ~((~ mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_21_lpi_1_dfm_st_3 | (~ (mul_loop_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | or_tmp_2227);
  assign mux_916_nl = MUX_s_1_2_2((nor_865_nl), (or_2317_nl), mul_loop_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm);
  assign mux_917_nl = MUX_s_1_2_2((mux_916_nl), mul_loop_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      or_90_cse);
  assign mux_918_nl = MUX_s_1_2_2((~ (FpMul_8U_23U_p_mant_p1_4_sva[47])), or_4956_cse,
      nor_181_cse);
  assign and_326_nl = mul_loop_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_918_nl);
  assign mux_919_nl = MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_66_itm, (and_326_nl),
      or_309_cse);
  assign or_2318_nl = (cfg_precision!=2'b10) | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_4_lpi_1_dfm_st_7;
  assign mux_920_nl = MUX_s_1_2_2((mux_919_nl), FpMul_8U_23U_FpMul_8U_23U_and_66_itm,
      or_2318_nl);
  assign or_2325_nl = nor_872_cse | (~ mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_22_lpi_1_dfm_st_3 | (mul_loop_mul_5_FpMul_8U_23U_p_mant_p1_mul_tmp[47])
      | mul_loop_mul_if_land_5_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign nor_863_nl = ~(nor_872_cse | (~ mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_22_lpi_1_dfm_st_3 | (~ (mul_loop_mul_5_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_if_land_5_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign mux_921_nl = MUX_s_1_2_2((nor_863_nl), (or_2325_nl), mul_loop_mul_5_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm);
  assign mux_922_nl = MUX_s_1_2_2((mux_921_nl), mul_loop_mul_5_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      or_90_cse);
  assign mux_923_nl = MUX_s_1_2_2((~ (FpMul_8U_23U_p_mant_p1_5_sva[47])), or_4953_cse,
      nor_197_cse);
  assign and_327_nl = mul_loop_mul_5_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_923_nl);
  assign mux_924_nl = MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_67_itm, (and_327_nl),
      or_309_cse);
  assign or_2329_nl = (cfg_precision!=2'b10) | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_5_lpi_1_dfm_st_7;
  assign mux_925_nl = MUX_s_1_2_2((mux_924_nl), FpMul_8U_23U_FpMul_8U_23U_and_67_itm,
      or_2329_nl);
  assign or_2336_nl = nor_872_cse | (~ mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_23_lpi_1_dfm_st_3 | (mul_loop_mul_6_FpMul_8U_23U_p_mant_p1_mul_tmp[47])
      | mul_loop_mul_if_land_6_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign nor_860_nl = ~(nor_872_cse | (~ mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_23_lpi_1_dfm_st_3 | (~ (mul_loop_mul_6_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_if_land_6_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign mux_926_nl = MUX_s_1_2_2((nor_860_nl), (or_2336_nl), mul_loop_mul_6_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm);
  assign mux_927_nl = MUX_s_1_2_2((mux_926_nl), mul_loop_mul_6_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      or_90_cse);
  assign nor_385_nl = ~((FpMul_8U_23U_p_mant_p1_6_sva[47]) | (~ mul_loop_mul_6_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2));
  assign mux_928_nl = MUX_s_1_2_2(and_tmp_72, or_tmp_2254, nor_385_nl);
  assign mux_929_nl = MUX_s_1_2_2(and_tmp_72, or_tmp_2254, and_2876_cse);
  assign mux_930_nl = MUX_s_1_2_2((mux_929_nl), (mux_928_nl), or_2342_cse);
  assign mux_931_nl = MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_68_itm, (mux_930_nl),
      or_309_cse);
  assign mux_932_nl = MUX_s_1_2_2((mux_931_nl), FpMul_8U_23U_FpMul_8U_23U_and_68_itm,
      or_90_cse);
  assign or_2347_nl = nor_872_cse | (~ mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_24_lpi_1_dfm_st_3 | (mul_loop_mul_7_FpMul_8U_23U_p_mant_p1_mul_tmp[47])
      | mul_loop_mul_if_land_7_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign nor_857_nl = ~(nor_872_cse | (~ mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_24_lpi_1_dfm_st_3 | (~ (mul_loop_mul_7_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_if_land_7_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign mux_933_nl = MUX_s_1_2_2((nor_857_nl), (or_2347_nl), mul_loop_mul_7_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm);
  assign mux_934_nl = MUX_s_1_2_2((mux_933_nl), mul_loop_mul_7_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      or_90_cse);
  assign mux_935_nl = MUX_s_1_2_2((~ (FpMul_8U_23U_p_mant_p1_7_sva[47])), or_4947_cse,
      nor_229_cse);
  assign and_329_nl = mul_loop_mul_7_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_935_nl);
  assign mux_936_nl = MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_69_itm, (and_329_nl),
      or_309_cse);
  assign or_2351_nl = (cfg_precision!=2'b10) | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_7_lpi_1_dfm_st_7;
  assign mux_937_nl = MUX_s_1_2_2((mux_936_nl), FpMul_8U_23U_FpMul_8U_23U_and_69_itm,
      or_2351_nl);
  assign or_2358_nl = nor_872_cse | (~ mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_25_lpi_1_dfm_st_3 | (mul_loop_mul_8_FpMul_8U_23U_p_mant_p1_mul_tmp[47])
      | mul_loop_mul_if_land_8_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign nor_854_nl = ~(nor_872_cse | (~ mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_25_lpi_1_dfm_st_3 | (~ (mul_loop_mul_8_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_if_land_8_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign mux_938_nl = MUX_s_1_2_2((nor_854_nl), (or_2358_nl), mul_loop_mul_8_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm);
  assign mux_939_nl = MUX_s_1_2_2((mux_938_nl), mul_loop_mul_8_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      or_90_cse);
  assign mux_940_nl = MUX_s_1_2_2((~ (FpMul_8U_23U_p_mant_p1_8_sva[47])), or_4944_cse,
      nor_245_cse);
  assign and_330_nl = mul_loop_mul_8_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_940_nl);
  assign mux_941_nl = MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_70_itm, (and_330_nl),
      or_309_cse);
  assign or_2362_nl = (cfg_precision!=2'b10) | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_8_lpi_1_dfm_st_7;
  assign mux_942_nl = MUX_s_1_2_2((mux_941_nl), FpMul_8U_23U_FpMul_8U_23U_and_70_itm,
      or_2362_nl);
  assign or_2369_nl = nor_872_cse | (~ mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_26_lpi_1_dfm_st_3 | (mul_loop_mul_9_FpMul_8U_23U_p_mant_p1_mul_tmp[47])
      | mul_loop_mul_if_land_9_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign nor_851_nl = ~(nor_872_cse | (~ mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_26_lpi_1_dfm_st_3 | (~ (mul_loop_mul_9_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_if_land_9_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign mux_943_nl = MUX_s_1_2_2((nor_851_nl), (or_2369_nl), mul_loop_mul_9_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm);
  assign mux_944_nl = MUX_s_1_2_2((mux_943_nl), mul_loop_mul_9_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      or_90_cse);
  assign mux_945_nl = MUX_s_1_2_2((~ (FpMul_8U_23U_p_mant_p1_9_sva[47])), or_4941_cse,
      nor_261_cse);
  assign and_331_nl = mul_loop_mul_9_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_945_nl);
  assign mux_946_nl = MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_71_itm, (and_331_nl),
      or_309_cse);
  assign or_2373_nl = (cfg_precision!=2'b10) | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_9_lpi_1_dfm_st_7;
  assign mux_947_nl = MUX_s_1_2_2((mux_946_nl), FpMul_8U_23U_FpMul_8U_23U_and_71_itm,
      or_2373_nl);
  assign or_2380_nl = nor_872_cse | (~ mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_27_lpi_1_dfm_st_3 | (mul_loop_mul_10_FpMul_8U_23U_p_mant_p1_mul_tmp[47])
      | mul_loop_mul_if_land_10_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign nor_848_nl = ~(nor_872_cse | (~ mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_27_lpi_1_dfm_st_3 | (~ (mul_loop_mul_10_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_if_land_10_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign mux_948_nl = MUX_s_1_2_2((nor_848_nl), (or_2380_nl), mul_loop_mul_10_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm);
  assign mux_949_nl = MUX_s_1_2_2((mux_948_nl), mul_loop_mul_10_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      or_90_cse);
  assign nor_392_nl = ~((FpMul_8U_23U_p_mant_p1_10_sva[47]) | (~ mul_loop_mul_10_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2));
  assign mux_950_nl = MUX_s_1_2_2(and_tmp_76, or_tmp_2298, nor_392_nl);
  assign mux_951_nl = MUX_s_1_2_2(and_tmp_76, or_tmp_2298, and_2868_cse);
  assign mux_952_nl = MUX_s_1_2_2((mux_951_nl), (mux_950_nl), or_2386_cse);
  assign mux_953_nl = MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_72_itm, (mux_952_nl),
      or_309_cse);
  assign mux_954_nl = MUX_s_1_2_2((mux_953_nl), FpMul_8U_23U_FpMul_8U_23U_and_72_itm,
      or_90_cse);
  assign or_2391_nl = (~ mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_28_lpi_1_dfm_st_3 | (mul_loop_mul_11_FpMul_8U_23U_p_mant_p1_mul_tmp[47])
      | or_tmp_1736;
  assign nor_846_nl = ~((~ mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_28_lpi_1_dfm_st_3 | (~ (mul_loop_mul_11_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | or_tmp_1736);
  assign mux_955_nl = MUX_s_1_2_2((nor_846_nl), (or_2391_nl), mul_loop_mul_11_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm);
  assign mux_956_nl = MUX_s_1_2_2((mux_955_nl), mul_loop_mul_11_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      or_90_cse);
  assign or_4652_nl = (~ (mul_loop_mul_11_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) |
      mul_loop_mul_11_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  assign mux_957_nl = MUX_s_1_2_2((~ (FpMul_8U_23U_p_mant_p1_11_sva[47])), (or_4652_nl),
      nor_283_cse);
  assign and_333_nl = mul_loop_mul_11_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_957_nl);
  assign mux_958_nl = MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_73_itm, (and_333_nl),
      or_309_cse);
  assign or_2392_nl = (cfg_precision!=2'b10) | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_11_lpi_1_dfm_st_7;
  assign mux_959_nl = MUX_s_1_2_2((mux_958_nl), FpMul_8U_23U_FpMul_8U_23U_and_73_itm,
      or_2392_nl);
  assign or_2400_nl = (mul_loop_mul_12_FpMul_8U_23U_p_mant_p1_mul_tmp[47]) | or_tmp_2310;
  assign and_2132_nl = (mul_loop_mul_12_FpMul_8U_23U_p_mant_p1_mul_tmp[47]) & (~
      or_tmp_2310);
  assign mux_960_nl = MUX_s_1_2_2((and_2132_nl), (or_2400_nl), mul_loop_mul_12_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm);
  assign or_2396_nl = (cfg_precision!=2'b10) | (~ mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_29_lpi_1_dfm_st_3;
  assign mux_961_nl = MUX_s_1_2_2((mux_960_nl), mul_loop_mul_12_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      or_2396_nl);
  assign mux_962_nl = MUX_s_1_2_2((~ (FpMul_8U_23U_p_mant_p1_12_sva[47])), or_4934_cse,
      nor_309_cse);
  assign and_334_nl = mul_loop_mul_12_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_962_nl);
  assign mux_963_nl = MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_74_itm, (and_334_nl),
      or_309_cse);
  assign or_2401_nl = (cfg_precision!=2'b10) | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_12_lpi_1_dfm_st_7;
  assign mux_964_nl = MUX_s_1_2_2((mux_963_nl), FpMul_8U_23U_FpMul_8U_23U_and_74_itm,
      or_2401_nl);
  assign or_2409_nl = (mul_loop_mul_13_FpMul_8U_23U_p_mant_p1_mul_tmp[47]) | or_tmp_2319;
  assign and_2131_nl = (mul_loop_mul_13_FpMul_8U_23U_p_mant_p1_mul_tmp[47]) & (~
      or_tmp_2319);
  assign mux_965_nl = MUX_s_1_2_2((and_2131_nl), (or_2409_nl), mul_loop_mul_13_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm);
  assign or_2405_nl = (cfg_precision!=2'b10) | (~ mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_30_lpi_1_dfm_st_3;
  assign mux_966_nl = MUX_s_1_2_2((mux_965_nl), mul_loop_mul_13_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      or_2405_nl);
  assign mux_967_nl = MUX_s_1_2_2((~ (FpMul_8U_23U_p_mant_p1_13_sva[47])), or_4931_cse,
      nor_325_cse);
  assign and_335_nl = mul_loop_mul_13_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_967_nl);
  assign mux_968_nl = MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_75_itm, (and_335_nl),
      or_309_cse);
  assign or_2410_nl = (cfg_precision!=2'b10) | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_13_lpi_1_dfm_st_7;
  assign mux_969_nl = MUX_s_1_2_2((mux_968_nl), FpMul_8U_23U_FpMul_8U_23U_and_75_itm,
      or_2410_nl);
  assign or_2417_nl = nor_872_cse | (~ mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_31_lpi_1_dfm_st_3 | (mul_loop_mul_14_FpMul_8U_23U_p_mant_p1_mul_tmp[47])
      | mul_loop_mul_if_land_14_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign nor_844_nl = ~(nor_872_cse | (~ mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_31_lpi_1_dfm_st_3 | (~ (mul_loop_mul_14_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_if_land_14_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign mux_970_nl = MUX_s_1_2_2((nor_844_nl), (or_2417_nl), mul_loop_mul_14_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm);
  assign mux_971_nl = MUX_s_1_2_2((mux_970_nl), mul_loop_mul_14_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      or_90_cse);
  assign or_2423_nl = (~ (mul_loop_mul_14_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) |
      mul_loop_mul_14_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7;
  assign mux_972_nl = MUX_s_1_2_2((~ (FpMul_8U_23U_p_mant_p1_14_sva[47])), (or_2423_nl),
      nor_340_cse);
  assign and_336_nl = mul_loop_mul_14_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_972_nl);
  assign mux_973_nl = MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_76_itm, (and_336_nl),
      or_309_cse);
  assign or_2421_nl = (cfg_precision!=2'b10) | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_14_lpi_1_dfm_st_7;
  assign mux_974_nl = MUX_s_1_2_2((mux_973_nl), FpMul_8U_23U_FpMul_8U_23U_and_76_itm,
      or_2421_nl);
  assign or_2428_nl = nor_872_cse | (~ mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_32_lpi_1_dfm_st_3 | (mul_loop_mul_15_FpMul_8U_23U_p_mant_p1_mul_tmp[47])
      | mul_loop_mul_if_land_15_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign nor_841_nl = ~(nor_872_cse | (~ mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_32_lpi_1_dfm_st_3 | (~ (mul_loop_mul_15_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_loop_mul_if_land_15_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3));
  assign mux_975_nl = MUX_s_1_2_2((nor_841_nl), (or_2428_nl), mul_loop_mul_15_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm);
  assign mux_976_nl = MUX_s_1_2_2((mux_975_nl), mul_loop_mul_15_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      or_90_cse);
  assign mux_977_nl = MUX_s_1_2_2((~ (FpMul_8U_23U_p_mant_p1_15_sva[47])), or_4927_cse,
      nor_356_cse);
  assign and_337_nl = mul_loop_mul_15_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_977_nl);
  assign mux_978_nl = MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_77_itm, (and_337_nl),
      or_309_cse);
  assign or_2432_nl = (cfg_precision!=2'b10) | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_15_lpi_1_dfm_st_7;
  assign mux_979_nl = MUX_s_1_2_2((mux_978_nl), FpMul_8U_23U_FpMul_8U_23U_and_77_itm,
      or_2432_nl);
  assign or_2439_nl = (~ mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | (mul_loop_mul_16_FpMul_8U_23U_p_mant_p1_mul_tmp[47])
      | mul_loop_mul_if_land_lpi_1_dfm_st_7 | io_read_cfg_mul_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign nor_899_nl = ~((~ (mul_loop_mul_16_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6 | mul_loop_mul_if_land_lpi_1_dfm_st_7
      | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | (~ mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign mux_980_nl = MUX_s_1_2_2((nor_899_nl), (or_2439_nl), mul_loop_mul_16_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm);
  assign mux_981_nl = MUX_s_1_2_2(mul_loop_mul_16_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      (mux_980_nl), or_309_cse);
  assign mux_982_nl = MUX_s_1_2_2((mux_981_nl), mul_loop_mul_16_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      or_90_cse);
  assign mux_983_nl = MUX_s_1_2_2((~ (FpMul_8U_23U_p_mant_p1_sva[47])), or_4924_cse,
      nor_372_cse);
  assign and_338_nl = mul_loop_mul_16_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_983_nl);
  assign mux_984_nl = MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_78_itm, (and_338_nl),
      or_309_cse);
  assign or_2442_nl = (cfg_precision!=2'b10) | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_st_6
      | mul_loop_mul_if_land_lpi_1_dfm_st_7;
  assign mux_985_nl = MUX_s_1_2_2((mux_984_nl), FpMul_8U_23U_FpMul_8U_23U_and_78_itm,
      or_2442_nl);
  assign mux_1123_nl = MUX_s_1_2_2(or_tmp_2492, or_tmp_2490, nor_53_cse);
  assign mux_1124_nl = MUX_s_1_2_2((~ or_309_cse), (mux_1123_nl), or_2577_cse);
  assign mux_1128_nl = MUX_s_1_2_2(mux_1680_itm, or_tmp_2490, reg_FpMul_8U_23U_lor_3_lpi_1_dfm_4_cse);
  assign and_344_nl = FpMul_8U_23U_lor_3_lpi_1_dfm_st & or_309_cse;
  assign mux_1131_nl = MUX_s_1_2_2((and_344_nl), or_tmp_2492, reg_FpMul_8U_23U_lor_3_lpi_1_dfm_4_cse);
  assign mux_1132_nl = MUX_s_1_2_2((mux_1131_nl), (mux_1128_nl), nor_53_cse);
  assign mux_1135_nl = MUX_s_1_2_2(mux_1680_itm, and_tmp_86, reg_FpMul_8U_23U_lor_3_lpi_1_dfm_4_cse);
  assign nor_824_nl = ~((cfg_precision[0]) | (~((cfg_precision[1]) & (mux_1135_nl))));
  assign mux_1136_nl = MUX_s_1_2_2((nor_824_nl), (mux_1132_nl), or_2577_cse);
  assign mux_1137_nl = MUX_s_1_2_2((mux_1136_nl), (mux_1124_nl), or_2576_cse);
  assign mux_1139_nl = MUX_s_1_2_2(or_tmp_2503, (mux_1137_nl), or_2575_cse);
  assign mux_1140_nl = MUX_s_1_2_2(or_tmp_2503, (mux_1139_nl), and_2130_cse);
  assign nand_133_nl = ~(or_309_cse & (~(mul_loop_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | mul_loop_mul_if_land_1_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2) | reg_FpMul_8U_23U_lor_3_lpi_1_dfm_4_cse)));
  assign nor_822_nl = ~((~ mul_loop_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1) | mul_loop_mul_if_land_1_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_1142_nl = MUX_s_1_2_2((nor_822_nl), nor_821_cse, reg_FpMul_8U_23U_lor_3_lpi_1_dfm_4_cse);
  assign and_2129_nl = or_309_cse & (mux_1142_nl);
  assign mux_1143_nl = MUX_s_1_2_2((and_2129_nl), (nand_133_nl), FpMul_8U_23U_lor_18_lpi_1_dfm_st);
  assign mux_1144_nl = MUX_s_1_2_2((mux_1143_nl), FpMul_8U_23U_lor_18_lpi_1_dfm_st,
      or_90_cse);
  assign mux_1145_nl = MUX_s_1_2_2(or_tmp_2523, or_tmp_2521, nor_53_cse);
  assign mux_1146_nl = MUX_s_1_2_2((~ or_309_cse), (mux_1145_nl), or_2608_cse);
  assign mux_1150_nl = MUX_s_1_2_2(mux_1681_itm, or_tmp_2521, reg_FpMul_8U_23U_lor_4_lpi_1_dfm_4_cse);
  assign and_348_nl = FpMul_8U_23U_lor_4_lpi_1_dfm_st & or_309_cse;
  assign mux_1153_nl = MUX_s_1_2_2((and_348_nl), or_tmp_2523, reg_FpMul_8U_23U_lor_4_lpi_1_dfm_4_cse);
  assign mux_1154_nl = MUX_s_1_2_2((mux_1153_nl), (mux_1150_nl), nor_53_cse);
  assign mux_1157_nl = MUX_s_1_2_2(mux_1681_itm, and_tmp_90, reg_FpMul_8U_23U_lor_4_lpi_1_dfm_4_cse);
  assign nor_817_nl = ~((cfg_precision[0]) | (~((cfg_precision[1]) & (mux_1157_nl))));
  assign mux_1158_nl = MUX_s_1_2_2((nor_817_nl), (mux_1154_nl), or_2608_cse);
  assign mux_1159_nl = MUX_s_1_2_2((mux_1158_nl), (mux_1146_nl), or_2607_cse);
  assign mux_1161_nl = MUX_s_1_2_2(or_tmp_2534, (mux_1159_nl), or_2575_cse);
  assign and_2128_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_2_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt;
  assign mux_1162_nl = MUX_s_1_2_2(or_tmp_2534, (mux_1161_nl), and_2128_nl);
  assign and_350_nl = FpMul_8U_23U_lor_19_lpi_1_dfm_st & or_tmp_129;
  assign mux_1164_nl = MUX_s_1_2_2((and_350_nl), or_tmp_2538, or_2628_cse);
  assign mux_1165_nl = MUX_s_1_2_2((mux_1164_nl), or_tmp_2538, reg_FpMul_8U_23U_lor_4_lpi_1_dfm_4_cse);
  assign mux_1166_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_19_lpi_1_dfm_st, (mux_1165_nl),
      or_309_cse);
  assign mux_1167_nl = MUX_s_1_2_2((mux_1166_nl), FpMul_8U_23U_lor_19_lpi_1_dfm_st,
      or_90_cse);
  assign mux_1168_nl = MUX_s_1_2_2(or_tmp_2546, or_tmp_2544, nor_53_cse);
  assign mux_1169_nl = MUX_s_1_2_2((~ or_309_cse), (mux_1168_nl), or_2631_cse);
  assign mux_1173_nl = MUX_s_1_2_2(mux_1682_itm, or_tmp_2544, reg_FpMul_8U_23U_lor_5_lpi_1_dfm_4_cse);
  assign and_353_nl = FpMul_8U_23U_lor_5_lpi_1_dfm_st & or_309_cse;
  assign mux_1176_nl = MUX_s_1_2_2((and_353_nl), or_tmp_2546, reg_FpMul_8U_23U_lor_5_lpi_1_dfm_4_cse);
  assign mux_1177_nl = MUX_s_1_2_2((mux_1176_nl), (mux_1173_nl), nor_53_cse);
  assign mux_1180_nl = MUX_s_1_2_2(mux_1682_itm, and_tmp_95, reg_FpMul_8U_23U_lor_5_lpi_1_dfm_4_cse);
  assign nor_815_nl = ~((cfg_precision[0]) | (~((cfg_precision[1]) & (mux_1180_nl))));
  assign mux_1181_nl = MUX_s_1_2_2((nor_815_nl), (mux_1177_nl), or_2631_cse);
  assign mux_1182_nl = MUX_s_1_2_2((mux_1181_nl), (mux_1169_nl), or_2630_cse);
  assign mux_1184_nl = MUX_s_1_2_2(or_tmp_2557, (mux_1182_nl), or_2575_cse);
  assign and_2127_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_3_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt;
  assign mux_1185_nl = MUX_s_1_2_2(or_tmp_2557, (mux_1184_nl), and_2127_nl);
  assign nand_135_nl = ~(or_309_cse & (~(mul_loop_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | mul_loop_mul_if_land_3_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2) | reg_FpMul_8U_23U_lor_5_lpi_1_dfm_4_cse)));
  assign nor_813_nl = ~((~ mul_loop_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1) | mul_loop_mul_if_land_3_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_1187_nl = MUX_s_1_2_2((nor_813_nl), nor_1477_cse, reg_FpMul_8U_23U_lor_5_lpi_1_dfm_4_cse);
  assign and_2126_nl = or_309_cse & (mux_1187_nl);
  assign mux_1188_nl = MUX_s_1_2_2((and_2126_nl), (nand_135_nl), FpMul_8U_23U_lor_20_lpi_1_dfm_st);
  assign mux_1189_nl = MUX_s_1_2_2((mux_1188_nl), FpMul_8U_23U_lor_20_lpi_1_dfm_st,
      or_90_cse);
  assign or_2667_nl = nor_872_cse | reg_FpMul_8U_23U_lor_6_lpi_1_dfm_4_cse | mul_loop_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | mul_loop_mul_if_land_4_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign or_2672_nl = (~ mul_loop_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1) | mul_loop_mul_if_land_4_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign mux_1192_nl = MUX_s_1_2_2((or_2672_nl), or_tmp_142, reg_FpMul_8U_23U_lor_6_lpi_1_dfm_4_cse);
  assign nor_808_nl = ~(nor_872_cse | (mux_1192_nl));
  assign mux_1193_nl = MUX_s_1_2_2((nor_808_nl), (or_2667_nl), FpMul_8U_23U_lor_21_lpi_1_dfm_st);
  assign mux_1194_nl = MUX_s_1_2_2((mux_1193_nl), FpMul_8U_23U_lor_21_lpi_1_dfm_st,
      or_90_cse);
  assign mux_1195_nl = MUX_s_1_2_2(or_tmp_2590, or_tmp_2588, nor_53_cse);
  assign mux_1196_nl = MUX_s_1_2_2((~ or_309_cse), (mux_1195_nl), or_2675_cse);
  assign mux_1200_nl = MUX_s_1_2_2(mux_1683_itm, or_tmp_2588, reg_FpMul_8U_23U_lor_7_lpi_1_dfm_4_cse);
  assign and_357_nl = FpMul_8U_23U_lor_7_lpi_1_dfm_st & or_309_cse;
  assign mux_1203_nl = MUX_s_1_2_2((and_357_nl), or_tmp_2590, reg_FpMul_8U_23U_lor_7_lpi_1_dfm_4_cse);
  assign mux_1204_nl = MUX_s_1_2_2((mux_1203_nl), (mux_1200_nl), nor_53_cse);
  assign mux_1207_nl = MUX_s_1_2_2(mux_1683_itm, and_tmp_99, reg_FpMul_8U_23U_lor_7_lpi_1_dfm_4_cse);
  assign nor_805_nl = ~((cfg_precision[0]) | (~((cfg_precision[1]) & (mux_1207_nl))));
  assign mux_1208_nl = MUX_s_1_2_2((nor_805_nl), (mux_1204_nl), or_2675_cse);
  assign mux_1209_nl = MUX_s_1_2_2((mux_1208_nl), (mux_1196_nl), or_414_cse);
  assign mux_1211_nl = MUX_s_1_2_2(or_tmp_2601, (mux_1209_nl), or_2575_cse);
  assign and_2125_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_5_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt;
  assign mux_1212_nl = MUX_s_1_2_2(or_tmp_2601, (mux_1211_nl), and_2125_nl);
  assign and_359_nl = FpMul_8U_23U_lor_22_lpi_1_dfm_st & or_tmp_148;
  assign mux_1214_nl = MUX_s_1_2_2((and_359_nl), or_tmp_2604, mul_loop_mul_5_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_1216_nl = MUX_s_1_2_2((mux_1214_nl), or_tmp_2604, reg_FpMul_8U_23U_lor_7_lpi_1_dfm_4_cse);
  assign mux_1217_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_22_lpi_1_dfm_st, (mux_1216_nl),
      or_309_cse);
  assign mux_1218_nl = MUX_s_1_2_2((mux_1217_nl), FpMul_8U_23U_lor_22_lpi_1_dfm_st,
      or_90_cse);
  assign or_2701_nl = nor_872_cse | reg_FpMul_8U_23U_lor_8_lpi_1_dfm_4_cse | mul_loop_mul_6_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | mul_loop_mul_if_land_6_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign or_2706_nl = (~ mul_loop_mul_6_FpMul_8U_23U_oelse_1_acc_itm_9_1) | mul_loop_mul_if_land_6_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign mux_1221_nl = MUX_s_1_2_2((or_2706_nl), or_tmp_152, reg_FpMul_8U_23U_lor_8_lpi_1_dfm_4_cse);
  assign nor_803_nl = ~(nor_872_cse | (mux_1221_nl));
  assign mux_1222_nl = MUX_s_1_2_2((nor_803_nl), (or_2701_nl), FpMul_8U_23U_lor_23_lpi_1_dfm_st);
  assign mux_1223_nl = MUX_s_1_2_2((mux_1222_nl), FpMul_8U_23U_lor_23_lpi_1_dfm_st,
      or_90_cse);
  assign or_2714_nl = nor_872_cse | reg_FpMul_8U_23U_lor_9_lpi_1_dfm_4_cse | mul_loop_mul_7_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | mul_loop_mul_if_land_7_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign or_2719_nl = (~ mul_loop_mul_7_FpMul_8U_23U_oelse_1_acc_itm_9_1) | mul_loop_mul_if_land_7_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign mux_1226_nl = MUX_s_1_2_2((or_2719_nl), or_tmp_156, reg_FpMul_8U_23U_lor_9_lpi_1_dfm_4_cse);
  assign nor_800_nl = ~(nor_872_cse | (mux_1226_nl));
  assign mux_1227_nl = MUX_s_1_2_2((nor_800_nl), (or_2714_nl), FpMul_8U_23U_lor_24_lpi_1_dfm_st);
  assign mux_1228_nl = MUX_s_1_2_2((mux_1227_nl), FpMul_8U_23U_lor_24_lpi_1_dfm_st,
      or_90_cse);
  assign mux_1229_nl = MUX_s_1_2_2(or_tmp_2637, or_tmp_2635, nor_53_cse);
  assign mux_1230_nl = MUX_s_1_2_2((~ or_309_cse), (mux_1229_nl), or_2722_cse);
  assign mux_1234_nl = MUX_s_1_2_2(mux_1684_itm, or_tmp_2635, reg_FpMul_8U_23U_lor_10_lpi_1_dfm_4_cse);
  assign and_362_nl = FpMul_8U_23U_lor_10_lpi_1_dfm_st & or_309_cse;
  assign mux_1237_nl = MUX_s_1_2_2((and_362_nl), or_tmp_2637, reg_FpMul_8U_23U_lor_10_lpi_1_dfm_4_cse);
  assign mux_1238_nl = MUX_s_1_2_2((mux_1237_nl), (mux_1234_nl), nor_53_cse);
  assign mux_1241_nl = MUX_s_1_2_2(mux_1684_itm, and_tmp_104, reg_FpMul_8U_23U_lor_10_lpi_1_dfm_4_cse);
  assign nor_797_nl = ~((cfg_precision[0]) | (~((cfg_precision[1]) & (mux_1241_nl))));
  assign mux_1242_nl = MUX_s_1_2_2((nor_797_nl), (mux_1238_nl), or_2722_cse);
  assign mux_1243_nl = MUX_s_1_2_2((mux_1242_nl), (mux_1230_nl), or_2721_cse);
  assign mux_1245_nl = MUX_s_1_2_2(or_tmp_2648, (mux_1243_nl), or_2575_cse);
  assign and_2124_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_8_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt;
  assign mux_1246_nl = MUX_s_1_2_2(or_tmp_2648, (mux_1245_nl), and_2124_nl);
  assign and_364_nl = FpMul_8U_23U_lor_25_lpi_1_dfm_st & or_tmp_162;
  assign mux_1248_nl = MUX_s_1_2_2((and_364_nl), or_tmp_2652, or_2742_cse);
  assign mux_1249_nl = MUX_s_1_2_2((mux_1248_nl), or_tmp_2652, reg_FpMul_8U_23U_lor_10_lpi_1_dfm_4_cse);
  assign mux_1250_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_25_lpi_1_dfm_st, (mux_1249_nl),
      or_309_cse);
  assign mux_1251_nl = MUX_s_1_2_2((mux_1250_nl), FpMul_8U_23U_lor_25_lpi_1_dfm_st,
      or_90_cse);
  assign mux_1252_nl = MUX_s_1_2_2(or_tmp_2660, or_tmp_2658, nor_53_cse);
  assign mux_1253_nl = MUX_s_1_2_2((~ or_309_cse), (mux_1252_nl), or_2745_cse);
  assign mux_1257_nl = MUX_s_1_2_2(mux_1685_itm, or_tmp_2658, reg_FpMul_8U_23U_lor_11_lpi_1_dfm_4_cse);
  assign and_367_nl = FpMul_8U_23U_lor_11_lpi_1_dfm_st & or_309_cse;
  assign mux_1260_nl = MUX_s_1_2_2((and_367_nl), or_tmp_2660, reg_FpMul_8U_23U_lor_11_lpi_1_dfm_4_cse);
  assign mux_1261_nl = MUX_s_1_2_2((mux_1260_nl), (mux_1257_nl), nor_53_cse);
  assign mux_1264_nl = MUX_s_1_2_2(mux_1685_itm, and_tmp_109, reg_FpMul_8U_23U_lor_11_lpi_1_dfm_4_cse);
  assign nor_795_nl = ~((cfg_precision[0]) | (~((cfg_precision[1]) & (mux_1264_nl))));
  assign mux_1265_nl = MUX_s_1_2_2((nor_795_nl), (mux_1261_nl), or_2745_cse);
  assign mux_1266_nl = MUX_s_1_2_2((mux_1265_nl), (mux_1253_nl), or_517_cse);
  assign mux_1268_nl = MUX_s_1_2_2(or_tmp_2671, (mux_1266_nl), or_2575_cse);
  assign and_2123_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_9_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt;
  assign mux_1269_nl = MUX_s_1_2_2(or_tmp_2671, (mux_1268_nl), and_2123_nl);
  assign and_369_nl = FpMul_8U_23U_lor_26_lpi_1_dfm_st & or_tmp_168;
  assign mux_1271_nl = MUX_s_1_2_2((and_369_nl), or_tmp_2674, mul_loop_mul_9_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign mux_1273_nl = MUX_s_1_2_2((mux_1271_nl), or_tmp_2674, reg_FpMul_8U_23U_lor_11_lpi_1_dfm_4_cse);
  assign mux_1274_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_26_lpi_1_dfm_st, (mux_1273_nl),
      or_309_cse);
  assign mux_1275_nl = MUX_s_1_2_2((mux_1274_nl), FpMul_8U_23U_lor_26_lpi_1_dfm_st,
      or_90_cse);
  assign or_2769_nl = (~ mul_loop_mul_10_FpMul_8U_23U_oelse_1_acc_itm_9_1) | mul_loop_mul_if_land_10_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign mux_1277_nl = MUX_s_1_2_2((or_2769_nl), or_tmp_172, reg_FpMul_8U_23U_lor_12_lpi_1_dfm_4_cse);
  assign mux_1278_nl = MUX_s_1_2_2((~ (mux_1277_nl)), or_tmp_460, FpMul_8U_23U_lor_27_lpi_1_dfm_st);
  assign mux_1279_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_27_lpi_1_dfm_st, (mux_1278_nl),
      or_309_cse);
  assign mux_1280_nl = MUX_s_1_2_2((mux_1279_nl), FpMul_8U_23U_lor_27_lpi_1_dfm_st,
      or_90_cse);
  assign or_2777_nl = nor_872_cse | reg_FpMul_8U_23U_lor_13_lpi_1_dfm_4_cse | mul_loop_mul_11_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | mul_loop_mul_if_land_11_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign or_2782_nl = (~ mul_loop_mul_11_FpMul_8U_23U_oelse_1_acc_itm_9_1) | mul_loop_mul_if_land_11_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign mux_1283_nl = MUX_s_1_2_2((or_2782_nl), or_tmp_176, reg_FpMul_8U_23U_lor_13_lpi_1_dfm_4_cse);
  assign nor_793_nl = ~(nor_872_cse | (mux_1283_nl));
  assign mux_1284_nl = MUX_s_1_2_2((nor_793_nl), (or_2777_nl), FpMul_8U_23U_lor_28_lpi_1_dfm_st);
  assign mux_1285_nl = MUX_s_1_2_2((mux_1284_nl), FpMul_8U_23U_lor_28_lpi_1_dfm_st,
      or_90_cse);
  assign or_2790_nl = nor_872_cse | reg_FpMul_8U_23U_lor_14_lpi_1_dfm_4_cse | mul_loop_mul_12_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | mul_loop_mul_if_land_12_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign or_2795_nl = (~ mul_loop_mul_12_FpMul_8U_23U_oelse_1_acc_itm_9_1) | mul_loop_mul_if_land_12_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign mux_1288_nl = MUX_s_1_2_2((or_2795_nl), or_tmp_180, reg_FpMul_8U_23U_lor_14_lpi_1_dfm_4_cse);
  assign nor_790_nl = ~(nor_872_cse | (mux_1288_nl));
  assign mux_1289_nl = MUX_s_1_2_2((nor_790_nl), (or_2790_nl), FpMul_8U_23U_lor_29_lpi_1_dfm_st);
  assign mux_1290_nl = MUX_s_1_2_2((mux_1289_nl), FpMul_8U_23U_lor_29_lpi_1_dfm_st,
      or_90_cse);
  assign mux_1291_nl = MUX_s_1_2_2(or_tmp_2713, or_tmp_2711, nor_53_cse);
  assign mux_1292_nl = MUX_s_1_2_2((~ or_309_cse), (mux_1291_nl), or_2798_cse);
  assign mux_1296_nl = MUX_s_1_2_2(mux_1686_itm, or_tmp_2711, reg_FpMul_8U_23U_lor_15_lpi_1_dfm_4_cse);
  assign and_372_nl = FpMul_8U_23U_lor_15_lpi_1_dfm_st & or_309_cse;
  assign mux_1299_nl = MUX_s_1_2_2((and_372_nl), or_tmp_2713, reg_FpMul_8U_23U_lor_15_lpi_1_dfm_4_cse);
  assign mux_1300_nl = MUX_s_1_2_2((mux_1299_nl), (mux_1296_nl), nor_53_cse);
  assign mux_1303_nl = MUX_s_1_2_2(mux_1686_itm, and_tmp_114, reg_FpMul_8U_23U_lor_15_lpi_1_dfm_4_cse);
  assign nor_787_nl = ~((cfg_precision[0]) | (~((cfg_precision[1]) & (mux_1303_nl))));
  assign mux_1304_nl = MUX_s_1_2_2((nor_787_nl), (mux_1300_nl), or_2798_cse);
  assign mux_1305_nl = MUX_s_1_2_2((mux_1304_nl), (mux_1292_nl), or_2797_cse);
  assign mux_1307_nl = MUX_s_1_2_2(or_tmp_2724, (mux_1305_nl), or_2575_cse);
  assign and_2122_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_13_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt;
  assign mux_1308_nl = MUX_s_1_2_2(or_tmp_2724, (mux_1307_nl), and_2122_nl);
  assign and_374_nl = FpMul_8U_23U_lor_30_lpi_1_dfm_st & or_tmp_186;
  assign mux_1310_nl = MUX_s_1_2_2((and_374_nl), or_tmp_2728, or_616_cse);
  assign mux_1311_nl = MUX_s_1_2_2((mux_1310_nl), or_tmp_2728, reg_FpMul_8U_23U_lor_15_lpi_1_dfm_4_cse);
  assign mux_1312_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_30_lpi_1_dfm_st, (mux_1311_nl),
      or_309_cse);
  assign mux_1313_nl = MUX_s_1_2_2((mux_1312_nl), FpMul_8U_23U_lor_30_lpi_1_dfm_st,
      or_90_cse);
  assign or_2826_nl = nor_872_cse | reg_FpMul_8U_23U_lor_16_lpi_1_dfm_4_cse | mul_loop_mul_14_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | mul_loop_mul_if_land_14_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2);
  assign or_2831_nl = (~ mul_loop_mul_14_FpMul_8U_23U_oelse_1_acc_itm_9_1) | mul_loop_mul_if_land_14_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2);
  assign mux_1316_nl = MUX_s_1_2_2((or_2831_nl), or_tmp_190, reg_FpMul_8U_23U_lor_16_lpi_1_dfm_4_cse);
  assign nor_785_nl = ~(nor_872_cse | (mux_1316_nl));
  assign mux_1317_nl = MUX_s_1_2_2((nor_785_nl), (or_2826_nl), FpMul_8U_23U_lor_31_lpi_1_dfm_st);
  assign mux_1318_nl = MUX_s_1_2_2((mux_1317_nl), FpMul_8U_23U_lor_31_lpi_1_dfm_st,
      or_90_cse);
  assign mux_1319_nl = MUX_s_1_2_2(or_tmp_2749, or_tmp_2747, nor_53_cse);
  assign mux_1320_nl = MUX_s_1_2_2((~ or_309_cse), (mux_1319_nl), or_2834_cse);
  assign mux_1324_nl = MUX_s_1_2_2(mux_1687_itm, or_tmp_2747, reg_FpMul_8U_23U_lor_17_lpi_1_dfm_4_cse);
  assign and_377_nl = FpMul_8U_23U_lor_17_lpi_1_dfm_st & or_309_cse;
  assign mux_1327_nl = MUX_s_1_2_2((and_377_nl), or_tmp_2749, reg_FpMul_8U_23U_lor_17_lpi_1_dfm_4_cse);
  assign mux_1328_nl = MUX_s_1_2_2((mux_1327_nl), (mux_1324_nl), nor_53_cse);
  assign mux_1331_nl = MUX_s_1_2_2(mux_1687_itm, and_tmp_119, reg_FpMul_8U_23U_lor_17_lpi_1_dfm_4_cse);
  assign nor_782_nl = ~((cfg_precision[0]) | (~((cfg_precision[1]) & (mux_1331_nl))));
  assign mux_1332_nl = MUX_s_1_2_2((nor_782_nl), (mux_1328_nl), or_2834_cse);
  assign mux_1333_nl = MUX_s_1_2_2((mux_1332_nl), (mux_1320_nl), or_2833_cse);
  assign mux_1335_nl = MUX_s_1_2_2(or_tmp_2760, (mux_1333_nl), or_2575_cse);
  assign and_2121_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_15_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt;
  assign mux_1336_nl = MUX_s_1_2_2(or_tmp_2760, (mux_1335_nl), and_2121_nl);
  assign nand_143_nl = ~(or_309_cse & (~(mul_loop_mul_15_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | mul_loop_mul_if_land_15_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | (~ main_stage_v_2) | reg_FpMul_8U_23U_lor_17_lpi_1_dfm_4_cse)));
  assign nor_780_nl = ~((~ mul_loop_mul_15_FpMul_8U_23U_oelse_1_acc_itm_9_1) | mul_loop_mul_if_land_15_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_1338_nl = MUX_s_1_2_2((nor_780_nl), nor_1413_cse, reg_FpMul_8U_23U_lor_17_lpi_1_dfm_4_cse);
  assign and_2120_nl = or_309_cse & (mux_1338_nl);
  assign mux_1339_nl = MUX_s_1_2_2((and_2120_nl), (nand_143_nl), FpMul_8U_23U_lor_32_lpi_1_dfm_st);
  assign mux_1340_nl = MUX_s_1_2_2((mux_1339_nl), FpMul_8U_23U_lor_32_lpi_1_dfm_st,
      or_90_cse);
  assign mux_1341_nl = MUX_s_1_2_2(or_tmp_2780, or_tmp_2778, nor_53_cse);
  assign mux_1342_nl = MUX_s_1_2_2((~ or_309_cse), (mux_1341_nl), or_2865_cse);
  assign mux_1346_nl = MUX_s_1_2_2(mux_1688_itm, or_tmp_2778, reg_FpMul_8U_23U_lor_lpi_1_dfm_4_cse);
  assign and_381_nl = FpMul_8U_23U_lor_lpi_1_dfm_st & or_309_cse;
  assign mux_1349_nl = MUX_s_1_2_2((and_381_nl), or_tmp_2780, reg_FpMul_8U_23U_lor_lpi_1_dfm_4_cse);
  assign mux_1350_nl = MUX_s_1_2_2((mux_1349_nl), (mux_1346_nl), nor_53_cse);
  assign mux_1353_nl = MUX_s_1_2_2(mux_1688_itm, and_tmp_123, reg_FpMul_8U_23U_lor_lpi_1_dfm_4_cse);
  assign nor_775_nl = ~((cfg_precision[0]) | (~((cfg_precision[1]) & (mux_1353_nl))));
  assign mux_1354_nl = MUX_s_1_2_2((nor_775_nl), (mux_1350_nl), or_2865_cse);
  assign mux_1355_nl = MUX_s_1_2_2((mux_1354_nl), (mux_1342_nl), or_2864_cse);
  assign mux_1357_nl = MUX_s_1_2_2(or_tmp_2791, (mux_1355_nl), or_2575_cse);
  assign and_2119_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt &
      cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt;
  assign mux_1358_nl = MUX_s_1_2_2(or_tmp_2791, (mux_1357_nl), and_2119_nl);
  assign and_383_nl = FpMul_8U_23U_lor_1_lpi_1_dfm_st & or_tmp_202;
  assign mux_1360_nl = MUX_s_1_2_2((and_383_nl), or_tmp_2795, or_2885_cse);
  assign mux_1361_nl = MUX_s_1_2_2((mux_1360_nl), or_tmp_2795, reg_FpMul_8U_23U_lor_lpi_1_dfm_4_cse);
  assign mux_1362_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_1_lpi_1_dfm_st, (mux_1361_nl),
      or_309_cse);
  assign mux_1363_nl = MUX_s_1_2_2((mux_1362_nl), FpMul_8U_23U_lor_1_lpi_1_dfm_st,
      or_90_cse);
  assign or_2967_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_7 | IsNaN_8U_23U_land_lpi_1_dfm_9
      | mul_loop_mul_if_land_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_6 | (~
      main_stage_v_2);
  assign mux_1446_nl = MUX_s_1_2_2(or_tmp_2177, (or_2967_nl), or_309_cse);
  assign or_2970_nl = mul_loop_mul_if_land_lpi_1_dfm_st_6 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_6 | (~
      main_stage_v_2);
  assign mux_1447_nl = MUX_s_1_2_2(or_tmp_2151, (or_2970_nl), or_309_cse);
  assign or_2973_nl = io_read_cfg_mul_bypass_rsc_svs_st_5 | mul_loop_mul_if_land_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_6 | (~ main_stage_v_2);
  assign mux_1448_nl = MUX_s_1_2_2(mux_tmp_490, (or_2973_nl), or_309_cse);
  assign or_2976_nl = IsNaN_8U_23U_1_land_15_lpi_1_dfm_7 | IsNaN_8U_23U_land_15_lpi_1_dfm_9
      | mul_loop_mul_if_land_15_lpi_1_dfm_st_6 | mul_loop_mul_if_land_15_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1449_nl = MUX_s_1_2_2(or_tmp_2097, (or_2976_nl), or_309_cse);
  assign or_2979_nl = mul_loop_mul_if_land_15_lpi_1_dfm_st_6 | mul_loop_mul_if_land_15_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1450_nl = MUX_s_1_2_2(or_tmp_2071, (or_2979_nl), or_309_cse);
  assign or_2984_nl = or_tmp_2894 | (~ main_stage_v_2);
  assign mux_1452_nl = MUX_s_1_2_2(mux_tmp_484, (or_2984_nl), or_309_cse);
  assign or_2987_nl = IsNaN_8U_23U_1_land_14_lpi_1_dfm_7 | IsNaN_8U_23U_land_14_lpi_1_dfm_9
      | mul_loop_mul_if_land_14_lpi_1_dfm_st_6 | mul_loop_mul_if_land_14_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1453_nl = MUX_s_1_2_2(or_tmp_2015, (or_2987_nl), or_309_cse);
  assign or_2990_nl = mul_loop_mul_if_land_14_lpi_1_dfm_st_6 | mul_loop_mul_if_land_14_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1454_nl = MUX_s_1_2_2(or_tmp_1991, (or_2990_nl), or_309_cse);
  assign or_2995_nl = or_tmp_2905 | (~ main_stage_v_2);
  assign mux_1456_nl = MUX_s_1_2_2(mux_tmp_478, (or_2995_nl), or_309_cse);
  assign or_2998_nl = IsNaN_8U_23U_1_land_13_lpi_1_dfm_7 | IsNaN_8U_23U_land_13_lpi_1_dfm_9
      | mul_loop_mul_if_land_13_lpi_1_dfm_st_6 | mul_loop_mul_if_land_13_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1457_nl = MUX_s_1_2_2(or_tmp_1931, (or_2998_nl), or_309_cse);
  assign or_3001_nl = mul_loop_mul_if_land_13_lpi_1_dfm_st_6 | mul_loop_mul_if_land_13_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1458_nl = MUX_s_1_2_2(or_tmp_1905, (or_3001_nl), or_309_cse);
  assign or_3006_nl = or_tmp_2916 | (~ main_stage_v_2);
  assign mux_1460_nl = MUX_s_1_2_2(mux_tmp_472, (or_3006_nl), or_309_cse);
  assign or_3009_nl = IsNaN_8U_23U_1_land_12_lpi_1_dfm_7 | IsNaN_8U_23U_land_12_lpi_1_dfm_9
      | mul_loop_mul_if_land_12_lpi_1_dfm_st_6 | mul_loop_mul_if_land_12_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1461_nl = MUX_s_1_2_2(or_tmp_1848, (or_3009_nl), or_309_cse);
  assign or_3012_nl = mul_loop_mul_if_land_12_lpi_1_dfm_st_6 | mul_loop_mul_if_land_12_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1462_nl = MUX_s_1_2_2(or_tmp_1822, (or_3012_nl), or_309_cse);
  assign or_3017_nl = or_tmp_2927 | (~ main_stage_v_2);
  assign mux_1464_nl = MUX_s_1_2_2(mux_tmp_466, (or_3017_nl), or_309_cse);
  assign or_3020_nl = IsNaN_8U_23U_1_land_11_lpi_1_dfm_7 | IsNaN_8U_23U_land_11_lpi_1_dfm_9
      | mul_loop_mul_if_land_11_lpi_1_dfm_st_6 | mul_loop_mul_if_land_11_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1465_nl = MUX_s_1_2_2(or_tmp_1765, (or_3020_nl), or_309_cse);
  assign or_3023_nl = mul_loop_mul_if_land_11_lpi_1_dfm_st_6 | mul_loop_mul_if_land_11_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1466_nl = MUX_s_1_2_2(or_tmp_1744, (or_3023_nl), or_309_cse);
  assign or_3028_nl = or_tmp_2938 | (~ main_stage_v_2);
  assign mux_1468_nl = MUX_s_1_2_2(mux_tmp_460, (or_3028_nl), or_309_cse);
  assign or_3031_nl = IsNaN_8U_23U_1_land_10_lpi_1_dfm_7 | IsNaN_8U_23U_land_10_lpi_1_dfm_9
      | mul_loop_mul_if_land_10_lpi_1_dfm_st_6 | mul_loop_mul_if_land_10_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1469_nl = MUX_s_1_2_2(or_tmp_1687, (or_3031_nl), or_309_cse);
  assign or_3034_nl = mul_loop_mul_if_land_10_lpi_1_dfm_st_6 | mul_loop_mul_if_land_10_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1470_nl = MUX_s_1_2_2(or_tmp_1661, (or_3034_nl), or_309_cse);
  assign or_3039_nl = or_tmp_2949 | (~ main_stage_v_2);
  assign mux_1472_nl = MUX_s_1_2_2(mux_tmp_454, (or_3039_nl), or_309_cse);
  assign or_3042_nl = IsNaN_8U_23U_1_land_9_lpi_1_dfm_7 | IsNaN_8U_23U_land_9_lpi_1_dfm_9
      | mul_loop_mul_if_land_9_lpi_1_dfm_st_6 | mul_loop_mul_if_land_9_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1473_nl = MUX_s_1_2_2(or_tmp_1607, (or_3042_nl), or_309_cse);
  assign or_3045_nl = mul_loop_mul_if_land_9_lpi_1_dfm_st_6 | mul_loop_mul_if_land_9_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1474_nl = MUX_s_1_2_2(or_tmp_1581, (or_3045_nl), or_309_cse);
  assign or_3050_nl = or_tmp_2960 | (~ main_stage_v_2);
  assign mux_1476_nl = MUX_s_1_2_2(mux_tmp_448, (or_3050_nl), or_309_cse);
  assign or_3053_nl = IsNaN_8U_23U_1_land_8_lpi_1_dfm_7 | IsNaN_8U_23U_land_8_lpi_1_dfm_9
      | mul_loop_mul_if_land_8_lpi_1_dfm_st_6 | mul_loop_mul_if_land_8_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1477_nl = MUX_s_1_2_2(or_tmp_1527, (or_3053_nl), or_309_cse);
  assign or_3056_nl = mul_loop_mul_if_land_8_lpi_1_dfm_st_6 | mul_loop_mul_if_land_8_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1478_nl = MUX_s_1_2_2(or_tmp_1501, (or_3056_nl), or_309_cse);
  assign or_3061_nl = or_tmp_2971 | (~ main_stage_v_2);
  assign mux_1480_nl = MUX_s_1_2_2(mux_tmp_442, (or_3061_nl), or_309_cse);
  assign or_3064_nl = IsNaN_8U_23U_1_land_7_lpi_1_dfm_7 | IsNaN_8U_23U_land_7_lpi_1_dfm_9
      | mul_loop_mul_if_land_7_lpi_1_dfm_st_6 | mul_loop_mul_if_land_7_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1481_nl = MUX_s_1_2_2(or_tmp_1447, (or_3064_nl), or_309_cse);
  assign or_3067_nl = mul_loop_mul_if_land_7_lpi_1_dfm_st_6 | mul_loop_mul_if_land_7_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1482_nl = MUX_s_1_2_2(or_tmp_1421, (or_3067_nl), or_309_cse);
  assign or_3072_nl = or_tmp_2982 | (~ main_stage_v_2);
  assign mux_1484_nl = MUX_s_1_2_2(mux_tmp_436, (or_3072_nl), or_309_cse);
  assign or_3075_nl = IsNaN_8U_23U_1_land_6_lpi_1_dfm_7 | IsNaN_8U_23U_land_6_lpi_1_dfm_9
      | mul_loop_mul_if_land_6_lpi_1_dfm_st_6 | mul_loop_mul_if_land_6_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1485_nl = MUX_s_1_2_2(or_tmp_1365, (or_3075_nl), or_309_cse);
  assign or_3078_nl = mul_loop_mul_if_land_6_lpi_1_dfm_st_6 | mul_loop_mul_if_land_6_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1486_nl = MUX_s_1_2_2(or_tmp_1339, (or_3078_nl), or_309_cse);
  assign or_3083_nl = or_tmp_2993 | (~ main_stage_v_2);
  assign mux_1488_nl = MUX_s_1_2_2(mux_tmp_430, (or_3083_nl), or_309_cse);
  assign or_3086_nl = IsNaN_8U_23U_1_land_5_lpi_1_dfm_7 | IsNaN_8U_23U_land_5_lpi_1_dfm_9
      | mul_loop_mul_if_land_5_lpi_1_dfm_st_6 | mul_loop_mul_if_land_5_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1489_nl = MUX_s_1_2_2(or_tmp_1283, (or_3086_nl), or_309_cse);
  assign or_3089_nl = mul_loop_mul_if_land_5_lpi_1_dfm_st_6 | mul_loop_mul_if_land_5_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1490_nl = MUX_s_1_2_2(or_tmp_1257, (or_3089_nl), or_309_cse);
  assign or_3094_nl = or_tmp_3004 | (~ main_stage_v_2);
  assign mux_1492_nl = MUX_s_1_2_2(mux_tmp_424, (or_3094_nl), or_309_cse);
  assign or_3097_nl = IsNaN_8U_23U_1_land_4_lpi_1_dfm_7 | IsNaN_8U_23U_land_4_lpi_1_dfm_9
      | mul_loop_mul_if_land_4_lpi_1_dfm_st_6 | mul_loop_mul_if_land_4_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1493_nl = MUX_s_1_2_2(or_tmp_1203, (or_3097_nl), or_309_cse);
  assign or_3100_nl = mul_loop_mul_if_land_4_lpi_1_dfm_st_6 | mul_loop_mul_if_land_4_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1494_nl = MUX_s_1_2_2(or_tmp_1177, (or_3100_nl), or_309_cse);
  assign or_3105_nl = or_tmp_3015 | (~ main_stage_v_2);
  assign mux_1496_nl = MUX_s_1_2_2(mux_tmp_418, (or_3105_nl), or_309_cse);
  assign or_3108_nl = IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 | IsNaN_8U_23U_land_3_lpi_1_dfm_9
      | mul_loop_mul_if_land_3_lpi_1_dfm_st_6 | mul_loop_mul_if_land_3_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1497_nl = MUX_s_1_2_2(or_tmp_1120, (or_3108_nl), or_309_cse);
  assign or_3111_nl = mul_loop_mul_if_land_3_lpi_1_dfm_st_6 | mul_loop_mul_if_land_3_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1498_nl = MUX_s_1_2_2(or_tmp_1094, (or_3111_nl), or_309_cse);
  assign or_3116_nl = or_tmp_3026 | (~ main_stage_v_2);
  assign mux_1500_nl = MUX_s_1_2_2(mux_tmp_412, (or_3116_nl), or_309_cse);
  assign or_3119_nl = IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 | IsNaN_8U_23U_land_2_lpi_1_dfm_9
      | mul_loop_mul_if_land_2_lpi_1_dfm_st_6 | mul_loop_mul_if_land_2_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1501_nl = MUX_s_1_2_2(or_tmp_1038, (or_3119_nl), or_309_cse);
  assign or_3122_nl = mul_loop_mul_if_land_2_lpi_1_dfm_st_6 | mul_loop_mul_if_land_2_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1502_nl = MUX_s_1_2_2(or_tmp_1012, (or_3122_nl), or_309_cse);
  assign or_3127_nl = or_tmp_3037 | (~ main_stage_v_2);
  assign mux_1504_nl = MUX_s_1_2_2(mux_tmp_406, (or_3127_nl), or_309_cse);
  assign or_3130_nl = IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 | IsNaN_8U_23U_land_1_lpi_1_dfm_9
      | mul_loop_mul_if_land_1_lpi_1_dfm_st_6 | mul_loop_mul_if_land_1_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1505_nl = MUX_s_1_2_2(or_tmp_958, (or_3130_nl), or_309_cse);
  assign or_3133_nl = mul_loop_mul_if_land_1_lpi_1_dfm_st_6 | mul_loop_mul_if_land_1_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | io_read_cfg_mul_bypass_rsc_svs_6 |
      (~ main_stage_v_2);
  assign mux_1506_nl = MUX_s_1_2_2(or_tmp_932, (or_3133_nl), or_309_cse);
  assign or_3138_nl = or_tmp_3048 | (~ main_stage_v_2);
  assign mux_1508_nl = MUX_s_1_2_2(mux_tmp_399, (or_3138_nl), or_309_cse);
  assign or_3143_nl = mul_loop_mul_else_land_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | io_read_cfg_mul_bypass_rsc_svs_6 | (~ main_stage_v_2);
  assign mux_1510_nl = MUX_s_1_2_2(mux_tmp_493, (or_3143_nl), or_309_cse);
  assign or_4633_nl = nor_872_cse | mux_tmp_1504;
  assign mux_1512_nl = MUX_s_1_2_2(mux_tmp_403, mux_tmp_1504, or_309_cse);
  assign mux_1513_nl = MUX_s_1_2_2((mux_1512_nl), (or_4633_nl), mul_loop_mul_else_land_15_lpi_1_dfm_9);
  assign or_4632_nl = nor_872_cse | mux_tmp_1507;
  assign mux_1515_nl = MUX_s_1_2_2(mux_tmp_403, mux_tmp_1507, or_309_cse);
  assign mux_1516_nl = MUX_s_1_2_2((mux_1515_nl), (or_4632_nl), mul_loop_mul_else_land_14_lpi_1_dfm_9);
  assign or_4631_nl = nor_872_cse | mux_tmp_1510;
  assign mux_1518_nl = MUX_s_1_2_2(mux_tmp_403, mux_tmp_1510, or_309_cse);
  assign mux_1519_nl = MUX_s_1_2_2((mux_1518_nl), (or_4631_nl), mul_loop_mul_else_land_13_lpi_1_dfm_9);
  assign or_4630_nl = nor_872_cse | mux_tmp_1513;
  assign mux_1521_nl = MUX_s_1_2_2(mux_tmp_403, mux_tmp_1513, or_309_cse);
  assign mux_1522_nl = MUX_s_1_2_2((mux_1521_nl), (or_4630_nl), mul_loop_mul_else_land_12_lpi_1_dfm_9);
  assign or_4629_nl = nor_872_cse | mux_tmp_1516;
  assign mux_1524_nl = MUX_s_1_2_2(mux_tmp_403, mux_tmp_1516, or_309_cse);
  assign mux_1525_nl = MUX_s_1_2_2((mux_1524_nl), (or_4629_nl), mul_loop_mul_else_land_11_lpi_1_dfm_9);
  assign or_3178_nl = mul_loop_mul_else_land_10_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | io_read_cfg_mul_bypass_rsc_svs_6 | (~ main_stage_v_2);
  assign mux_1527_nl = MUX_s_1_2_2(mux_tmp_457, (or_3178_nl), or_309_cse);
  assign or_3183_nl = mul_loop_mul_else_land_9_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | io_read_cfg_mul_bypass_rsc_svs_6 | (~ main_stage_v_2);
  assign mux_1529_nl = MUX_s_1_2_2(mux_tmp_451, (or_3183_nl), or_309_cse);
  assign or_3188_nl = mul_loop_mul_else_land_8_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | io_read_cfg_mul_bypass_rsc_svs_6 | (~ main_stage_v_2);
  assign mux_1531_nl = MUX_s_1_2_2(mux_tmp_445, (or_3188_nl), or_309_cse);
  assign or_3193_nl = mul_loop_mul_else_land_7_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | io_read_cfg_mul_bypass_rsc_svs_6 | (~ main_stage_v_2);
  assign mux_1533_nl = MUX_s_1_2_2(mux_tmp_439, (or_3193_nl), or_309_cse);
  assign or_3198_nl = mul_loop_mul_else_land_6_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | io_read_cfg_mul_bypass_rsc_svs_6 | (~ main_stage_v_2);
  assign mux_1535_nl = MUX_s_1_2_2(mux_tmp_433, (or_3198_nl), or_309_cse);
  assign or_3203_nl = mul_loop_mul_else_land_5_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | io_read_cfg_mul_bypass_rsc_svs_6 | (~ main_stage_v_2);
  assign mux_1537_nl = MUX_s_1_2_2(mux_tmp_427, (or_3203_nl), or_309_cse);
  assign or_3208_nl = mul_loop_mul_else_land_4_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | io_read_cfg_mul_bypass_rsc_svs_6 | (~ main_stage_v_2);
  assign mux_1539_nl = MUX_s_1_2_2(mux_tmp_421, (or_3208_nl), or_309_cse);
  assign or_3213_nl = mul_loop_mul_else_land_3_lpi_1_dfm_8 | io_read_cfg_mul_bypass_rsc_svs_st_5
      | io_read_cfg_mul_bypass_rsc_svs_6 | (~ main_stage_v_2);
  assign mux_1541_nl = MUX_s_1_2_2(mux_tmp_415, (or_3213_nl), or_309_cse);
  assign or_4628_nl = nor_872_cse | mux_tmp_1535;
  assign mux_1543_nl = MUX_s_1_2_2(mux_tmp_403, mux_tmp_1535, or_309_cse);
  assign mux_1544_nl = MUX_s_1_2_2((mux_1543_nl), (or_4628_nl), mul_loop_mul_else_land_2_lpi_1_dfm_9);
  assign or_4627_nl = nor_872_cse | mux_tmp_1538;
  assign mux_1546_nl = MUX_s_1_2_2(mux_tmp_403, mux_tmp_1538, or_309_cse);
  assign mux_1547_nl = MUX_s_1_2_2((mux_1546_nl), (or_4627_nl), mul_loop_mul_else_land_1_lpi_1_dfm_9);
  assign mux_1430_nl = MUX_s_1_2_2(and_384_cse, or_2577_cse, FpMul_8U_23U_lor_3_lpi_1_dfm_st);
  assign and_385_nl = FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_tmp & mux_tmp_1427;
  assign mux_1438_nl = MUX_s_1_2_2(mux_tmp_1430, (and_385_nl), or_2575_cse);
  assign mux_1439_nl = MUX_s_1_2_2(mux_tmp_1430, (mux_1438_nl), and_2130_cse);
  assign mux_1440_nl = MUX_s_1_2_2((mux_1439_nl), (mux_1430_nl), or_90_cse);
  assign or_2963_nl = reg_FpMul_8U_23U_lor_3_lpi_1_dfm_4_cse | mul_loop_mul_if_land_1_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5;
  assign mux_1441_nl = MUX_s_1_2_2(not_tmp_845, or_2577_cse, or_2963_nl);
  assign and_2500_nl = and_384_cse & reg_FpMul_8U_23U_lor_3_lpi_1_dfm_4_cse;
  assign mux_1444_nl = MUX_s_1_2_2((and_2500_nl), (mux_1441_nl), FpMul_8U_23U_lor_3_lpi_1_dfm_st);
  assign mux_1445_nl = MUX_s_1_2_2((mux_1444_nl), (mux_1440_nl), or_309_cse);
  assign and_2099_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_1_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~(((io_read_cfg_mul_bypass_rsc_svs_5 | mul_loop_mul_if_land_1_lpi_1_dfm_7)
      & IsNaN_8U_23U_land_1_lpi_1_dfm_8) | nor_749_cse));
  assign nor_750_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_1_lpi_1_dfm_st_6 | (or_tmp_3048 & IsNaN_8U_23U_land_1_lpi_1_dfm_9));
  assign mux_1548_nl = MUX_s_1_2_2((nor_750_nl), (and_2099_nl), or_309_cse);
  assign and_2096_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_2_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~(((io_read_cfg_mul_bypass_rsc_svs_5 | mul_loop_mul_if_land_2_lpi_1_dfm_7)
      & IsNaN_8U_23U_land_2_lpi_1_dfm_8) | nor_749_cse));
  assign nor_747_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_2_lpi_1_dfm_st_6 | (or_tmp_3037 & IsNaN_8U_23U_land_2_lpi_1_dfm_9));
  assign mux_1549_nl = MUX_s_1_2_2((nor_747_nl), (and_2096_nl), or_309_cse);
  assign and_2093_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_3_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~(((io_read_cfg_mul_bypass_rsc_svs_5 | mul_loop_mul_if_land_3_lpi_1_dfm_7)
      & IsNaN_8U_23U_land_3_lpi_1_dfm_8) | nor_749_cse));
  assign nor_744_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_3_lpi_1_dfm_st_6 | (or_tmp_3026 & IsNaN_8U_23U_land_3_lpi_1_dfm_9));
  assign mux_1550_nl = MUX_s_1_2_2((nor_744_nl), (and_2093_nl), or_309_cse);
  assign and_2090_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_4_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~(((io_read_cfg_mul_bypass_rsc_svs_5 | mul_loop_mul_if_land_4_lpi_1_dfm_7)
      & IsNaN_8U_23U_land_4_lpi_1_dfm_8) | nor_749_cse));
  assign nor_741_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_4_lpi_1_dfm_st_6 | (or_tmp_3015 & IsNaN_8U_23U_land_4_lpi_1_dfm_9));
  assign mux_1551_nl = MUX_s_1_2_2((nor_741_nl), (and_2090_nl), or_309_cse);
  assign and_2087_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_5_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~(((io_read_cfg_mul_bypass_rsc_svs_5 | mul_loop_mul_if_land_5_lpi_1_dfm_7)
      & IsNaN_8U_23U_land_5_lpi_1_dfm_8) | nor_749_cse));
  assign nor_738_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_5_lpi_1_dfm_st_6 | (or_tmp_3004 & IsNaN_8U_23U_land_5_lpi_1_dfm_9));
  assign mux_1552_nl = MUX_s_1_2_2((nor_738_nl), (and_2087_nl), or_309_cse);
  assign and_2084_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_6_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~(((io_read_cfg_mul_bypass_rsc_svs_5 | mul_loop_mul_if_land_6_lpi_1_dfm_7)
      & IsNaN_8U_23U_land_6_lpi_1_dfm_8) | nor_749_cse));
  assign nor_735_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_6_lpi_1_dfm_st_6 | (or_tmp_2993 & IsNaN_8U_23U_land_6_lpi_1_dfm_9));
  assign mux_1553_nl = MUX_s_1_2_2((nor_735_nl), (and_2084_nl), or_309_cse);
  assign and_2081_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_7_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~(((io_read_cfg_mul_bypass_rsc_svs_5 | mul_loop_mul_if_land_7_lpi_1_dfm_7)
      & IsNaN_8U_23U_land_7_lpi_1_dfm_8) | nor_749_cse));
  assign nor_732_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_7_lpi_1_dfm_st_6 | (or_tmp_2982 & IsNaN_8U_23U_land_7_lpi_1_dfm_9));
  assign mux_1554_nl = MUX_s_1_2_2((nor_732_nl), (and_2081_nl), or_309_cse);
  assign and_2078_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_8_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~(((io_read_cfg_mul_bypass_rsc_svs_5 | mul_loop_mul_if_land_8_lpi_1_dfm_7)
      & IsNaN_8U_23U_land_8_lpi_1_dfm_8) | nor_749_cse));
  assign nor_729_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_8_lpi_1_dfm_st_6 | (or_tmp_2971 & IsNaN_8U_23U_land_8_lpi_1_dfm_9));
  assign mux_1555_nl = MUX_s_1_2_2((nor_729_nl), (and_2078_nl), or_309_cse);
  assign and_2075_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_9_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~(((io_read_cfg_mul_bypass_rsc_svs_5 | mul_loop_mul_if_land_9_lpi_1_dfm_7)
      & IsNaN_8U_23U_land_9_lpi_1_dfm_8) | nor_749_cse));
  assign nor_726_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_9_lpi_1_dfm_st_6 | (or_tmp_2960 & IsNaN_8U_23U_land_9_lpi_1_dfm_9));
  assign mux_1556_nl = MUX_s_1_2_2((nor_726_nl), (and_2075_nl), or_309_cse);
  assign and_2072_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_10_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~(((io_read_cfg_mul_bypass_rsc_svs_5 | mul_loop_mul_if_land_10_lpi_1_dfm_7)
      & IsNaN_8U_23U_land_10_lpi_1_dfm_8) | nor_749_cse));
  assign nor_723_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_10_lpi_1_dfm_st_6 | (or_tmp_2949 & IsNaN_8U_23U_land_10_lpi_1_dfm_9));
  assign mux_1557_nl = MUX_s_1_2_2((nor_723_nl), (and_2072_nl), or_309_cse);
  assign and_2069_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_11_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~(((io_read_cfg_mul_bypass_rsc_svs_5 | mul_loop_mul_if_land_11_lpi_1_dfm_7)
      & IsNaN_8U_23U_land_11_lpi_1_dfm_8) | nor_749_cse));
  assign nor_720_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_11_lpi_1_dfm_st_6 | (or_tmp_2938 & IsNaN_8U_23U_land_11_lpi_1_dfm_9));
  assign mux_1558_nl = MUX_s_1_2_2((nor_720_nl), (and_2069_nl), or_309_cse);
  assign and_2066_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_12_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~(((io_read_cfg_mul_bypass_rsc_svs_5 | mul_loop_mul_if_land_12_lpi_1_dfm_7)
      & IsNaN_8U_23U_land_12_lpi_1_dfm_8) | nor_749_cse));
  assign nor_717_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_12_lpi_1_dfm_st_6 | (or_tmp_2927 & IsNaN_8U_23U_land_12_lpi_1_dfm_9));
  assign mux_1559_nl = MUX_s_1_2_2((nor_717_nl), (and_2066_nl), or_309_cse);
  assign and_2063_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_13_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~(((io_read_cfg_mul_bypass_rsc_svs_5 | mul_loop_mul_if_land_13_lpi_1_dfm_7)
      & IsNaN_8U_23U_land_13_lpi_1_dfm_8) | nor_749_cse));
  assign nor_714_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_13_lpi_1_dfm_st_6 | (or_tmp_2916 & IsNaN_8U_23U_land_13_lpi_1_dfm_9));
  assign mux_1560_nl = MUX_s_1_2_2((nor_714_nl), (and_2063_nl), or_309_cse);
  assign and_2060_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_14_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~(((io_read_cfg_mul_bypass_rsc_svs_5 | mul_loop_mul_if_land_14_lpi_1_dfm_7)
      & IsNaN_8U_23U_land_14_lpi_1_dfm_8) | nor_749_cse));
  assign nor_711_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_14_lpi_1_dfm_st_6 | (or_tmp_2905 & IsNaN_8U_23U_land_14_lpi_1_dfm_9));
  assign mux_1561_nl = MUX_s_1_2_2((nor_711_nl), (and_2060_nl), or_309_cse);
  assign and_2057_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_15_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~(((io_read_cfg_mul_bypass_rsc_svs_5 | mul_loop_mul_if_land_15_lpi_1_dfm_7)
      & IsNaN_8U_23U_land_15_lpi_1_dfm_8) | nor_749_cse));
  assign nor_708_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_15_lpi_1_dfm_st_6 | (or_tmp_2894 & IsNaN_8U_23U_land_15_lpi_1_dfm_9));
  assign mux_1562_nl = MUX_s_1_2_2((nor_708_nl), (and_2057_nl), or_309_cse);
  assign and_2054_nl = main_stage_v_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1) &
      (~ mul_loop_mul_if_land_lpi_1_dfm_st_5) & cfg_mul_op_rsc_triosy_obj_bawt &
      cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt
      & (~(((io_read_cfg_mul_bypass_rsc_svs_5 | mul_loop_mul_if_land_lpi_1_dfm_7)
      & IsNaN_8U_23U_land_lpi_1_dfm_8) | nor_749_cse));
  assign nor_705_nl = ~((~ main_stage_v_2) | io_read_cfg_mul_bypass_rsc_svs_st_5
      | mul_loop_mul_if_land_lpi_1_dfm_st_6 | ((io_read_cfg_mul_bypass_rsc_svs_6
      | mul_loop_mul_if_land_lpi_1_dfm_8) & IsNaN_8U_23U_land_lpi_1_dfm_9));
  assign mux_1563_nl = MUX_s_1_2_2((nor_705_nl), (and_2054_nl), or_309_cse);
  assign and_2052_nl = main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt & cfg_mul_bypass_rsc_triosy_obj_bawt
      & cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt & (~
      io_read_cfg_mul_bypass_rsc_svs_5) & (~ mul_loop_mul_else_land_lpi_1_dfm_7);
  assign and_2053_nl = or_2575_cse & main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~ io_read_cfg_mul_bypass_rsc_svs_5) & (~
      mul_loop_mul_else_land_lpi_1_dfm_7);
  assign mux_1564_nl = MUX_s_1_2_2((and_2053_nl), (and_2052_nl), io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign nor_702_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_6 | mul_loop_mul_else_land_lpi_1_dfm_8);
  assign mux_1565_nl = MUX_s_1_2_2((nor_702_nl), (mux_1564_nl), or_309_cse);
  assign and_2050_nl = main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt & cfg_mul_bypass_rsc_triosy_obj_bawt
      & cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt & (~
      io_read_cfg_mul_bypass_rsc_svs_5) & (~ mul_loop_mul_else_land_15_lpi_1_dfm_7);
  assign and_2051_nl = or_2575_cse & main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~ io_read_cfg_mul_bypass_rsc_svs_5) & (~
      mul_loop_mul_else_land_15_lpi_1_dfm_7);
  assign mux_1566_nl = MUX_s_1_2_2((and_2051_nl), (and_2050_nl), io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign nor_701_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_6 | mul_loop_mul_else_land_15_lpi_1_dfm_8);
  assign mux_1567_nl = MUX_s_1_2_2((nor_701_nl), (mux_1566_nl), or_309_cse);
  assign and_2048_nl = main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt & cfg_mul_bypass_rsc_triosy_obj_bawt
      & cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt & (~
      io_read_cfg_mul_bypass_rsc_svs_5) & (~ mul_loop_mul_else_land_14_lpi_1_dfm_7);
  assign and_2049_nl = or_2575_cse & main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~ io_read_cfg_mul_bypass_rsc_svs_5) & (~
      mul_loop_mul_else_land_14_lpi_1_dfm_7);
  assign mux_1568_nl = MUX_s_1_2_2((and_2049_nl), (and_2048_nl), io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign nor_700_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_6 | mul_loop_mul_else_land_14_lpi_1_dfm_8);
  assign mux_1569_nl = MUX_s_1_2_2((nor_700_nl), (mux_1568_nl), or_309_cse);
  assign and_2046_nl = main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt & cfg_mul_bypass_rsc_triosy_obj_bawt
      & cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt & (~
      io_read_cfg_mul_bypass_rsc_svs_5) & (~ mul_loop_mul_else_land_13_lpi_1_dfm_7);
  assign and_2047_nl = or_2575_cse & main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~ io_read_cfg_mul_bypass_rsc_svs_5) & (~
      mul_loop_mul_else_land_13_lpi_1_dfm_7);
  assign mux_1570_nl = MUX_s_1_2_2((and_2047_nl), (and_2046_nl), io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign nor_699_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_6 | mul_loop_mul_else_land_13_lpi_1_dfm_8);
  assign mux_1571_nl = MUX_s_1_2_2((nor_699_nl), (mux_1570_nl), or_309_cse);
  assign and_2044_nl = main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt & cfg_mul_bypass_rsc_triosy_obj_bawt
      & cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt & (~
      io_read_cfg_mul_bypass_rsc_svs_5) & (~ mul_loop_mul_else_land_12_lpi_1_dfm_7);
  assign and_2045_nl = or_2575_cse & main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~ io_read_cfg_mul_bypass_rsc_svs_5) & (~
      mul_loop_mul_else_land_12_lpi_1_dfm_7);
  assign mux_1572_nl = MUX_s_1_2_2((and_2045_nl), (and_2044_nl), io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign nor_698_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_6 | mul_loop_mul_else_land_12_lpi_1_dfm_8);
  assign mux_1573_nl = MUX_s_1_2_2((nor_698_nl), (mux_1572_nl), or_309_cse);
  assign and_2042_nl = main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt & cfg_mul_bypass_rsc_triosy_obj_bawt
      & cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt & (~
      io_read_cfg_mul_bypass_rsc_svs_5) & (~ mul_loop_mul_else_land_11_lpi_1_dfm_7);
  assign and_2043_nl = or_2575_cse & main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~ io_read_cfg_mul_bypass_rsc_svs_5) & (~
      mul_loop_mul_else_land_11_lpi_1_dfm_7);
  assign mux_1574_nl = MUX_s_1_2_2((and_2043_nl), (and_2042_nl), io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign nor_697_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_6 | mul_loop_mul_else_land_11_lpi_1_dfm_8);
  assign mux_1575_nl = MUX_s_1_2_2((nor_697_nl), (mux_1574_nl), or_309_cse);
  assign and_2040_nl = main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt & cfg_mul_bypass_rsc_triosy_obj_bawt
      & cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt & (~
      io_read_cfg_mul_bypass_rsc_svs_5) & (~ mul_loop_mul_else_land_10_lpi_1_dfm_7);
  assign and_2041_nl = or_2575_cse & main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~ io_read_cfg_mul_bypass_rsc_svs_5) & (~
      mul_loop_mul_else_land_10_lpi_1_dfm_7);
  assign mux_1576_nl = MUX_s_1_2_2((and_2041_nl), (and_2040_nl), io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign nor_696_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_6 | mul_loop_mul_else_land_10_lpi_1_dfm_8);
  assign mux_1577_nl = MUX_s_1_2_2((nor_696_nl), (mux_1576_nl), or_309_cse);
  assign and_2038_nl = main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt & cfg_mul_bypass_rsc_triosy_obj_bawt
      & cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt & (~
      io_read_cfg_mul_bypass_rsc_svs_5) & (~ mul_loop_mul_else_land_9_lpi_1_dfm_7);
  assign and_2039_nl = or_2575_cse & main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~ io_read_cfg_mul_bypass_rsc_svs_5) & (~
      mul_loop_mul_else_land_9_lpi_1_dfm_7);
  assign mux_1578_nl = MUX_s_1_2_2((and_2039_nl), (and_2038_nl), io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign nor_695_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_6 | mul_loop_mul_else_land_9_lpi_1_dfm_8);
  assign mux_1579_nl = MUX_s_1_2_2((nor_695_nl), (mux_1578_nl), or_309_cse);
  assign and_2036_nl = main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt & cfg_mul_bypass_rsc_triosy_obj_bawt
      & cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt & (~
      io_read_cfg_mul_bypass_rsc_svs_5) & (~ mul_loop_mul_else_land_8_lpi_1_dfm_7);
  assign and_2037_nl = or_2575_cse & main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~ io_read_cfg_mul_bypass_rsc_svs_5) & (~
      mul_loop_mul_else_land_8_lpi_1_dfm_7);
  assign mux_1580_nl = MUX_s_1_2_2((and_2037_nl), (and_2036_nl), io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign nor_694_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_6 | mul_loop_mul_else_land_8_lpi_1_dfm_8);
  assign mux_1581_nl = MUX_s_1_2_2((nor_694_nl), (mux_1580_nl), or_309_cse);
  assign and_2034_nl = main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt & cfg_mul_bypass_rsc_triosy_obj_bawt
      & cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt & (~
      io_read_cfg_mul_bypass_rsc_svs_5) & (~ mul_loop_mul_else_land_7_lpi_1_dfm_7);
  assign and_2035_nl = or_2575_cse & main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~ io_read_cfg_mul_bypass_rsc_svs_5) & (~
      mul_loop_mul_else_land_7_lpi_1_dfm_7);
  assign mux_1582_nl = MUX_s_1_2_2((and_2035_nl), (and_2034_nl), io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign nor_693_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_6 | mul_loop_mul_else_land_7_lpi_1_dfm_8);
  assign mux_1583_nl = MUX_s_1_2_2((nor_693_nl), (mux_1582_nl), or_309_cse);
  assign and_2032_nl = main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt & cfg_mul_bypass_rsc_triosy_obj_bawt
      & cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt & (~
      io_read_cfg_mul_bypass_rsc_svs_5) & (~ mul_loop_mul_else_land_6_lpi_1_dfm_7);
  assign and_2033_nl = or_2575_cse & main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~ io_read_cfg_mul_bypass_rsc_svs_5) & (~
      mul_loop_mul_else_land_6_lpi_1_dfm_7);
  assign mux_1584_nl = MUX_s_1_2_2((and_2033_nl), (and_2032_nl), io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign nor_692_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_6 | mul_loop_mul_else_land_6_lpi_1_dfm_8);
  assign mux_1585_nl = MUX_s_1_2_2((nor_692_nl), (mux_1584_nl), or_309_cse);
  assign and_2030_nl = main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt & cfg_mul_bypass_rsc_triosy_obj_bawt
      & cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt & (~
      io_read_cfg_mul_bypass_rsc_svs_5) & (~ mul_loop_mul_else_land_5_lpi_1_dfm_7);
  assign and_2031_nl = or_2575_cse & main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~ io_read_cfg_mul_bypass_rsc_svs_5) & (~
      mul_loop_mul_else_land_5_lpi_1_dfm_7);
  assign mux_1586_nl = MUX_s_1_2_2((and_2031_nl), (and_2030_nl), io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign nor_691_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_6 | mul_loop_mul_else_land_5_lpi_1_dfm_8);
  assign mux_1587_nl = MUX_s_1_2_2((nor_691_nl), (mux_1586_nl), or_309_cse);
  assign and_2028_nl = main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt & cfg_mul_bypass_rsc_triosy_obj_bawt
      & cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt & (~
      io_read_cfg_mul_bypass_rsc_svs_5) & (~ mul_loop_mul_else_land_4_lpi_1_dfm_7);
  assign and_2029_nl = or_2575_cse & main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~ io_read_cfg_mul_bypass_rsc_svs_5) & (~
      mul_loop_mul_else_land_4_lpi_1_dfm_7);
  assign mux_1588_nl = MUX_s_1_2_2((and_2029_nl), (and_2028_nl), io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign nor_690_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_6 | mul_loop_mul_else_land_4_lpi_1_dfm_8);
  assign mux_1589_nl = MUX_s_1_2_2((nor_690_nl), (mux_1588_nl), or_309_cse);
  assign and_2026_nl = main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt & cfg_mul_bypass_rsc_triosy_obj_bawt
      & cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt & (~
      io_read_cfg_mul_bypass_rsc_svs_5) & (~ mul_loop_mul_else_land_3_lpi_1_dfm_7);
  assign and_2027_nl = or_2575_cse & main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~ io_read_cfg_mul_bypass_rsc_svs_5) & (~
      mul_loop_mul_else_land_3_lpi_1_dfm_7);
  assign mux_1590_nl = MUX_s_1_2_2((and_2027_nl), (and_2026_nl), io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign nor_689_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_6 | mul_loop_mul_else_land_3_lpi_1_dfm_8);
  assign mux_1591_nl = MUX_s_1_2_2((nor_689_nl), (mux_1590_nl), or_309_cse);
  assign and_2024_nl = main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt & cfg_mul_bypass_rsc_triosy_obj_bawt
      & cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt & (~
      io_read_cfg_mul_bypass_rsc_svs_5) & (~ mul_loop_mul_else_land_2_lpi_1_dfm_7);
  assign and_2025_nl = or_2575_cse & main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~ io_read_cfg_mul_bypass_rsc_svs_5) & (~
      mul_loop_mul_else_land_2_lpi_1_dfm_7);
  assign mux_1592_nl = MUX_s_1_2_2((and_2025_nl), (and_2024_nl), io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign nor_688_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_6 | mul_loop_mul_else_land_2_lpi_1_dfm_8);
  assign mux_1593_nl = MUX_s_1_2_2((nor_688_nl), (mux_1592_nl), or_309_cse);
  assign and_2022_nl = main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt & cfg_mul_bypass_rsc_triosy_obj_bawt
      & cfg_mul_prelu_rsc_triosy_obj_bawt & cfg_mul_src_rsc_triosy_obj_bawt & (~
      io_read_cfg_mul_bypass_rsc_svs_5) & (~ mul_loop_mul_else_land_1_lpi_1_dfm_7);
  assign and_2023_nl = or_2575_cse & main_stage_v_1 & cfg_mul_op_rsc_triosy_obj_bawt
      & cfg_mul_bypass_rsc_triosy_obj_bawt & cfg_mul_prelu_rsc_triosy_obj_bawt &
      cfg_mul_src_rsc_triosy_obj_bawt & (~ io_read_cfg_mul_bypass_rsc_svs_5) & (~
      mul_loop_mul_else_land_1_lpi_1_dfm_7);
  assign mux_1594_nl = MUX_s_1_2_2((and_2023_nl), (and_2022_nl), io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign nor_687_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2)
      | io_read_cfg_mul_bypass_rsc_svs_6 | mul_loop_mul_else_land_1_lpi_1_dfm_8);
  assign mux_1595_nl = MUX_s_1_2_2((nor_687_nl), (mux_1594_nl), or_309_cse);
  assign nor_684_nl = ~(nor_749_cse | mul_loop_mul_if_land_1_lpi_1_dfm_st_5 | IsNaN_8U_23U_land_1_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | not_tmp_30);
  assign nor_686_nl = ~(IsNaN_8U_23U_land_1_lpi_1_dfm_9 | mul_loop_mul_if_land_1_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_1596_nl = MUX_s_1_2_2((nor_686_nl), (nor_684_nl), or_309_cse);
  assign nor_681_nl = ~(nor_749_cse | IsNaN_8U_23U_land_2_lpi_1_dfm_8 | mul_loop_mul_if_land_2_lpi_1_dfm_st_5
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | not_tmp_30);
  assign nor_683_nl = ~(IsNaN_8U_23U_land_2_lpi_1_dfm_9 | mul_loop_mul_if_land_2_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_1597_nl = MUX_s_1_2_2((nor_683_nl), (nor_681_nl), or_309_cse);
  assign nor_678_nl = ~(nor_749_cse | mul_loop_mul_if_land_3_lpi_1_dfm_st_5 | IsNaN_8U_23U_land_3_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | not_tmp_30);
  assign nor_680_nl = ~(IsNaN_8U_23U_land_3_lpi_1_dfm_9 | mul_loop_mul_if_land_3_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_1598_nl = MUX_s_1_2_2((nor_680_nl), (nor_678_nl), or_309_cse);
  assign nor_675_nl = ~(mul_loop_mul_if_land_4_lpi_1_dfm_st_5 | nor_749_cse | IsNaN_8U_23U_land_4_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | not_tmp_30);
  assign nor_677_nl = ~(IsNaN_8U_23U_land_4_lpi_1_dfm_9 | mul_loop_mul_if_land_4_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_1599_nl = MUX_s_1_2_2((nor_677_nl), (nor_675_nl), or_309_cse);
  assign nor_672_nl = ~(nor_749_cse | IsNaN_8U_23U_land_5_lpi_1_dfm_8 | mul_loop_mul_if_land_5_lpi_1_dfm_st_5
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | not_tmp_30);
  assign nor_674_nl = ~(IsNaN_8U_23U_land_5_lpi_1_dfm_9 | mul_loop_mul_if_land_5_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_1600_nl = MUX_s_1_2_2((nor_674_nl), (nor_672_nl), or_309_cse);
  assign nor_669_nl = ~(mul_loop_mul_if_land_6_lpi_1_dfm_st_5 | nor_749_cse | IsNaN_8U_23U_land_6_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | not_tmp_30);
  assign nor_671_nl = ~(IsNaN_8U_23U_land_6_lpi_1_dfm_9 | mul_loop_mul_if_land_6_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_1601_nl = MUX_s_1_2_2((nor_671_nl), (nor_669_nl), or_309_cse);
  assign nor_666_nl = ~(mul_loop_mul_if_land_7_lpi_1_dfm_st_5 | nor_749_cse | IsNaN_8U_23U_land_7_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | not_tmp_30);
  assign nor_668_nl = ~(IsNaN_8U_23U_land_7_lpi_1_dfm_9 | mul_loop_mul_if_land_7_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_1602_nl = MUX_s_1_2_2((nor_668_nl), (nor_666_nl), or_309_cse);
  assign nor_663_nl = ~(nor_749_cse | mul_loop_mul_if_land_8_lpi_1_dfm_st_5 | IsNaN_8U_23U_land_8_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | not_tmp_30);
  assign nor_665_nl = ~(IsNaN_8U_23U_land_8_lpi_1_dfm_9 | mul_loop_mul_if_land_8_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_1603_nl = MUX_s_1_2_2((nor_665_nl), (nor_663_nl), or_309_cse);
  assign nor_660_nl = ~(nor_749_cse | mul_loop_mul_if_land_9_lpi_1_dfm_st_5 | IsNaN_8U_23U_land_9_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | not_tmp_30);
  assign nor_662_nl = ~(IsNaN_8U_23U_land_9_lpi_1_dfm_9 | mul_loop_mul_if_land_9_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_1604_nl = MUX_s_1_2_2((nor_662_nl), (nor_660_nl), or_309_cse);
  assign nor_657_nl = ~(mul_loop_mul_if_land_10_lpi_1_dfm_st_5 | nor_749_cse | IsNaN_8U_23U_land_10_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | not_tmp_30);
  assign nor_659_nl = ~(IsNaN_8U_23U_land_10_lpi_1_dfm_9 | mul_loop_mul_if_land_10_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_1605_nl = MUX_s_1_2_2((nor_659_nl), (nor_657_nl), or_309_cse);
  assign nor_654_nl = ~(mul_loop_mul_if_land_11_lpi_1_dfm_st_5 | nor_749_cse | IsNaN_8U_23U_land_11_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | not_tmp_30);
  assign nor_656_nl = ~(IsNaN_8U_23U_land_11_lpi_1_dfm_9 | mul_loop_mul_if_land_11_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_1606_nl = MUX_s_1_2_2((nor_656_nl), (nor_654_nl), or_309_cse);
  assign nor_651_nl = ~(mul_loop_mul_if_land_12_lpi_1_dfm_st_5 | nor_749_cse | IsNaN_8U_23U_land_12_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | not_tmp_30);
  assign nor_653_nl = ~(IsNaN_8U_23U_land_12_lpi_1_dfm_9 | mul_loop_mul_if_land_12_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_1607_nl = MUX_s_1_2_2((nor_653_nl), (nor_651_nl), or_309_cse);
  assign nor_648_nl = ~(nor_749_cse | mul_loop_mul_if_land_13_lpi_1_dfm_st_5 | IsNaN_8U_23U_land_13_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | not_tmp_30);
  assign nor_650_nl = ~(IsNaN_8U_23U_land_13_lpi_1_dfm_9 | mul_loop_mul_if_land_13_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_1608_nl = MUX_s_1_2_2((nor_650_nl), (nor_648_nl), or_309_cse);
  assign nor_645_nl = ~(mul_loop_mul_if_land_14_lpi_1_dfm_st_5 | nor_749_cse | IsNaN_8U_23U_land_14_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | not_tmp_30);
  assign nor_647_nl = ~(IsNaN_8U_23U_land_14_lpi_1_dfm_9 | mul_loop_mul_if_land_14_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_1609_nl = MUX_s_1_2_2((nor_647_nl), (nor_645_nl), or_309_cse);
  assign nor_642_nl = ~(nor_749_cse | mul_loop_mul_if_land_15_lpi_1_dfm_st_5 | IsNaN_8U_23U_land_15_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | not_tmp_30);
  assign nor_644_nl = ~(IsNaN_8U_23U_land_15_lpi_1_dfm_9 | mul_loop_mul_if_land_15_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_1610_nl = MUX_s_1_2_2((nor_644_nl), (nor_642_nl), or_309_cse);
  assign nor_639_nl = ~(nor_749_cse | mul_loop_mul_if_land_lpi_1_dfm_st_5 | IsNaN_8U_23U_land_lpi_1_dfm_8
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | not_tmp_30);
  assign nor_641_nl = ~(IsNaN_8U_23U_land_lpi_1_dfm_9 | mul_loop_mul_if_land_lpi_1_dfm_st_6
      | io_read_cfg_mul_bypass_rsc_svs_st_5 | (~ main_stage_v_2));
  assign mux_1611_nl = MUX_s_1_2_2((nor_641_nl), (nor_639_nl), or_309_cse);
  function [0:0] MUX1HOT_s_1_1_2;
    input [0:0] input_0;
    input [0:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction
  function [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction
  function [9:0] MUX1HOT_v_10_3_2;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [2:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    MUX1HOT_v_10_3_2 = result;
  end
  endfunction
  function [9:0] MUX1HOT_v_10_4_2;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [3:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    result = result | ( input_3 & {10{sel[3]}});
    MUX1HOT_v_10_4_2 = result;
  end
  endfunction
  function [17:0] MUX1HOT_v_18_3_2;
    input [17:0] input_2;
    input [17:0] input_1;
    input [17:0] input_0;
    input [2:0] sel;
    reg [17:0] result;
  begin
    result = input_0 & {18{sel[0]}};
    result = result | ( input_1 & {18{sel[1]}});
    result = result | ( input_2 & {18{sel[2]}});
    MUX1HOT_v_18_3_2 = result;
  end
  endfunction
  function [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    result = result | ( input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction
  function [2:0] MUX1HOT_v_3_4_2;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [3:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    result = result | ( input_3 & {3{sel[3]}});
    MUX1HOT_v_3_4_2 = result;
  end
  endfunction
  function [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction
  function [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction
  function [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction
  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction
  function [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction
  function [22:0] MUX_v_23_2_2;
    input [22:0] input_0;
    input [22:0] input_1;
    input [0:0] sel;
    reg [22:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_23_2_2 = result;
  end
  endfunction
  function [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction
  function [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction
  function [45:0] MUX_v_46_2_2;
    input [45:0] input_0;
    input [45:0] input_1;
    input [0:0] sel;
    reg [45:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_46_2_2 = result;
  end
  endfunction
  function [47:0] MUX_v_48_2_2;
    input [47:0] input_0;
    input [47:0] input_1;
    input [0:0] sel;
    reg [47:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_48_2_2 = result;
  end
  endfunction
  function [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction
  function [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction
  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction
  function [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction
  function [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction
  function [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction
  function [7:0] readslicef_9_8_1;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_9_8_1 = tmp[7:0];
  end
  endfunction
  function [17:0] signext_18_2;
    input [1:0] vector;
  begin
    signext_18_2= {{16{vector[1]}}, vector};
  end
  endfunction
  function [9:0] conv_s2s_9_10 ;
    input [8:0] vector ;
  begin
    conv_s2s_9_10 = {vector[8], vector};
  end
  endfunction
  function [48:0] conv_s2u_49_49 ;
    input [48:0] vector ;
  begin
    conv_s2u_49_49 = vector;
  end
  endfunction
  function [8:0] conv_u2s_8_9 ;
    input [7:0] vector ;
  begin
    conv_u2s_8_9 = {1'b0, vector};
  end
  endfunction
  function [9:0] conv_u2s_8_10 ;
    input [7:0] vector ;
  begin
    conv_u2s_8_10 = {{2{1'b0}}, vector};
  end
  endfunction
  function [22:0] conv_u2u_1_23 ;
    input [0:0] vector ;
  begin
    conv_u2u_1_23 = {{22{1'b0}}, vector};
  end
  endfunction
  function [3:0] conv_u2u_3_4 ;
    input [2:0] vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction
  function [5:0] conv_u2u_5_6 ;
    input [4:0] vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction
  function [8:0] conv_u2u_8_9 ;
    input [7:0] vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction
  function [47:0] conv_u2u_48_48 ;
    input [47:0] vector ;
  begin
    conv_u2u_48_48 = vector;
  end
  endfunction
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_trt_core
// ------------------------------------------------------------------
module SDP_X_X_trt_core (
  nvdla_core_clk, nvdla_core_rstn, chn_trt_in_rsc_slz, chn_trt_in_rsc_sz, chn_trt_in_rsc_z,
      chn_trt_in_rsc_vz, chn_trt_in_rsc_lz, cfg_mul_shift_value_rsc_triosy_lz, cfg_precision,
      chn_trt_out_rsc_z, chn_trt_out_rsc_vz, chn_trt_out_rsc_lz, chn_trt_in_rsci_oswt,
      chn_trt_in_rsci_oswt_unreg, cfg_mul_shift_value_rsci_d, chn_trt_out_rsci_oswt,
      cfg_mul_shift_value_rsc_triosy_obj_oswt, chn_trt_out_rsci_oswt_unreg_pff
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output chn_trt_in_rsc_slz;
  input chn_trt_in_rsc_sz;
  input [799:0] chn_trt_in_rsc_z;
  input chn_trt_in_rsc_vz;
  output chn_trt_in_rsc_lz;
  output cfg_mul_shift_value_rsc_triosy_lz;
  input [1:0] cfg_precision;
  output [511:0] chn_trt_out_rsc_z;
  input chn_trt_out_rsc_vz;
  output chn_trt_out_rsc_lz;
  input chn_trt_in_rsci_oswt;
  output chn_trt_in_rsci_oswt_unreg;
  input [5:0] cfg_mul_shift_value_rsci_d;
  input chn_trt_out_rsci_oswt;
  input cfg_mul_shift_value_rsc_triosy_obj_oswt;
  output chn_trt_out_rsci_oswt_unreg_pff;
// Interconnect Declarations
  wire core_wen;
  reg chn_trt_in_rsci_iswt0;
  wire chn_trt_in_rsci_bawt;
  wire chn_trt_in_rsci_wen_comp;
  reg chn_trt_in_rsci_ld_core_psct;
  wire [799:0] chn_trt_in_rsci_d_mxwt;
  wire core_wten;
  wire chn_trt_out_rsci_bawt;
  wire chn_trt_out_rsci_wen_comp;
  wire cfg_mul_shift_value_rsc_triosy_obj_bawt;
  reg chn_trt_out_rsci_d_511;
  reg [29:0] chn_trt_out_rsci_d_510_481;
  reg chn_trt_out_rsci_d_480;
  reg chn_trt_out_rsci_d_479;
  reg [29:0] chn_trt_out_rsci_d_478_449;
  reg chn_trt_out_rsci_d_448;
  reg chn_trt_out_rsci_d_447;
  reg [29:0] chn_trt_out_rsci_d_446_417;
  reg chn_trt_out_rsci_d_416;
  reg chn_trt_out_rsci_d_415;
  reg [29:0] chn_trt_out_rsci_d_414_385;
  reg chn_trt_out_rsci_d_384;
  reg chn_trt_out_rsci_d_383;
  reg [29:0] chn_trt_out_rsci_d_382_353;
  reg chn_trt_out_rsci_d_352;
  reg chn_trt_out_rsci_d_351;
  reg [29:0] chn_trt_out_rsci_d_350_321;
  reg chn_trt_out_rsci_d_320;
  reg chn_trt_out_rsci_d_319;
  reg [29:0] chn_trt_out_rsci_d_318_289;
  reg chn_trt_out_rsci_d_288;
  reg chn_trt_out_rsci_d_287;
  reg [29:0] chn_trt_out_rsci_d_286_257;
  reg chn_trt_out_rsci_d_256;
  reg chn_trt_out_rsci_d_255;
  reg [29:0] chn_trt_out_rsci_d_254_225;
  reg chn_trt_out_rsci_d_224;
  reg chn_trt_out_rsci_d_223;
  reg [29:0] chn_trt_out_rsci_d_222_193;
  reg chn_trt_out_rsci_d_192;
  reg chn_trt_out_rsci_d_191;
  reg [29:0] chn_trt_out_rsci_d_190_161;
  reg chn_trt_out_rsci_d_160;
  reg chn_trt_out_rsci_d_159;
  reg [29:0] chn_trt_out_rsci_d_158_129;
  reg chn_trt_out_rsci_d_128;
  reg chn_trt_out_rsci_d_127;
  reg [29:0] chn_trt_out_rsci_d_126_97;
  reg chn_trt_out_rsci_d_96;
  reg chn_trt_out_rsci_d_95;
  reg [29:0] chn_trt_out_rsci_d_94_65;
  reg chn_trt_out_rsci_d_64;
  reg chn_trt_out_rsci_d_63;
  reg [29:0] chn_trt_out_rsci_d_62_33;
  reg chn_trt_out_rsci_d_32;
  reg chn_trt_out_rsci_d_31;
  reg [29:0] chn_trt_out_rsci_d_30_1;
  reg chn_trt_out_rsci_d_0;
  wire [1:0] fsm_output;
  wire and_dcpl_1;
  wire or_dcpl;
  wire and_dcpl_3;
  wire or_dcpl_3;
  wire and_dcpl_7;
  wire and_dcpl_11;
  wire and_dcpl_15;
  wire and_dcpl_17;
  wire and_dcpl_19;
  wire not_tmp_9;
  wire and_dcpl_23;
  wire and_dcpl_24;
  wire and_dcpl_134;
  wire or_tmp_150;
  wire and_148_cse;
  wire and_150_cse;
  wire and_4_mdf;
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_sva;
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_15_sva;
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_14_sva;
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_13_sva;
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_12_sva;
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_11_sva;
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_10_sva;
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_9_sva;
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_8_sva;
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_7_sva;
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_6_sva;
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_5_sva;
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_4_sva;
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_3_sva;
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_2_sva;
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_1_sva;
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva;
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva;
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva;
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva;
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva;
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva;
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva;
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva;
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva;
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva;
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva;
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva;
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva;
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva;
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva;
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva;
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva;
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva;
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva;
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva;
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva;
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva;
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva;
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva;
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva;
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva;
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva;
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva;
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva;
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva;
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva;
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva;
  wire chn_trt_out_and_2_cse;
  reg reg_cfg_mul_shift_value_rsc_triosy_obj_ld_core_psct_cse;
  reg reg_chn_trt_out_rsci_ld_core_psct_cse;
  wire chn_trt_in_rsci_ld_core_psct_mx0c0;
  wire chn_trt_out_rsci_d_0_mx0c1;
  wire chn_trt_out_rsci_d_30_1_mx0c1;
  wire chn_trt_out_rsci_d_62_33_mx0c1;
  wire chn_trt_out_rsci_d_94_65_mx0c1;
  wire chn_trt_out_rsci_d_126_97_mx0c1;
  wire chn_trt_out_rsci_d_158_129_mx0c1;
  wire chn_trt_out_rsci_d_190_161_mx0c1;
  wire chn_trt_out_rsci_d_222_193_mx0c1;
  wire chn_trt_out_rsci_d_254_225_mx0c1;
  wire chn_trt_out_rsci_d_286_257_mx0c1;
  wire chn_trt_out_rsci_d_318_289_mx0c1;
  wire chn_trt_out_rsci_d_350_321_mx0c1;
  wire chn_trt_out_rsci_d_382_353_mx0c1;
  wire chn_trt_out_rsci_d_414_385_mx0c1;
  wire chn_trt_out_rsci_d_446_417_mx0c1;
  wire chn_trt_out_rsci_d_478_449_mx0c1;
  wire chn_trt_out_rsci_d_510_481_mx0c1;
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_1_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_1_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_2_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_2_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_3_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_3_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_4_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_4_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_5_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_5_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_6_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_6_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_7_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_7_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_8_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_8_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_9_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_9_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_10_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_10_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_11_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_11_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_12_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_12_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_13_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_13_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_14_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_14_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_15_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_15_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_sva;
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_sva;
  wire[0:0] trt_loop_else_mux_112_nl;
  wire[0:0] trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  wire[29:0] trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  wire[29:0] trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_113_nl;
  wire[0:0] trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_114_nl;
  wire[0:0] trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  wire[29:0] trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  wire[29:0] trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_115_nl;
  wire[0:0] trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_116_nl;
  wire[0:0] trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  wire[29:0] trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  wire[29:0] trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_117_nl;
  wire[0:0] trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_118_nl;
  wire[0:0] trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  wire[29:0] trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  wire[29:0] trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_119_nl;
  wire[0:0] trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_120_nl;
  wire[0:0] trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  wire[29:0] trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  wire[29:0] trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_121_nl;
  wire[0:0] trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_122_nl;
  wire[0:0] trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  wire[29:0] trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  wire[29:0] trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_123_nl;
  wire[0:0] trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_124_nl;
  wire[0:0] trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  wire[29:0] trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  wire[29:0] trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_125_nl;
  wire[0:0] trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_126_nl;
  wire[0:0] trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  wire[29:0] trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  wire[29:0] trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_127_nl;
  wire[0:0] trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_128_nl;
  wire[0:0] trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  wire[29:0] trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  wire[29:0] trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_129_nl;
  wire[0:0] trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_130_nl;
  wire[0:0] trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  wire[29:0] trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  wire[29:0] trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_131_nl;
  wire[0:0] trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_132_nl;
  wire[0:0] trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  wire[29:0] trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  wire[29:0] trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_133_nl;
  wire[0:0] trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_134_nl;
  wire[0:0] trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  wire[29:0] trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  wire[29:0] trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_135_nl;
  wire[0:0] trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_136_nl;
  wire[0:0] trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  wire[29:0] trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  wire[29:0] trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_137_nl;
  wire[0:0] trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_138_nl;
  wire[0:0] trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  wire[29:0] trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  wire[29:0] trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_139_nl;
  wire[0:0] trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_140_nl;
  wire[0:0] trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  wire[29:0] trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  wire[29:0] trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_141_nl;
  wire[0:0] trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_142_nl;
  wire[0:0] trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  wire[29:0] trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  wire[29:0] trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_else_mux_143_nl;
  wire[0:0] trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  wire[0:0] trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  wire[0:0] trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  wire[0:0] trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  wire[0:0] trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  wire[0:0] trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  wire[0:0] trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  wire[0:0] trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  wire[0:0] trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  wire[0:0] trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  wire[0:0] trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  wire[0:0] trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  wire[0:0] trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  wire[0:0] trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  wire[0:0] trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  wire[0:0] trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  wire[0:0] trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  wire[0:0] mux_4_nl;
  wire[0:0] mux_5_nl;
  wire[0:0] mux_6_nl;
  wire[0:0] mux_7_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] mux_9_nl;
  wire[0:0] mux_10_nl;
  wire[0:0] mux_11_nl;
  wire[0:0] mux_12_nl;
  wire[0:0] mux_13_nl;
  wire[0:0] mux_14_nl;
  wire[0:0] mux_15_nl;
  wire[0:0] mux_16_nl;
  wire[0:0] mux_17_nl;
  wire[0:0] mux_18_nl;
  wire[0:0] mux_19_nl;
// Interconnect Declarations for Component Instantiations
  wire [111:0] nl_trt_loop_1_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  assign nl_trt_loop_1_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = {(chn_trt_in_rsci_d_mxwt[48:0])
      , 63'b0};
  wire [111:0] nl_trt_loop_2_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  assign nl_trt_loop_2_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = {(chn_trt_in_rsci_d_mxwt[97:49])
      , 63'b0};
  wire [111:0] nl_trt_loop_3_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  assign nl_trt_loop_3_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = {(chn_trt_in_rsci_d_mxwt[146:98])
      , 63'b0};
  wire [111:0] nl_trt_loop_4_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  assign nl_trt_loop_4_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = {(chn_trt_in_rsci_d_mxwt[195:147])
      , 63'b0};
  wire [111:0] nl_trt_loop_5_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  assign nl_trt_loop_5_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = {(chn_trt_in_rsci_d_mxwt[244:196])
      , 63'b0};
  wire [111:0] nl_trt_loop_6_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  assign nl_trt_loop_6_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = {(chn_trt_in_rsci_d_mxwt[293:245])
      , 63'b0};
  wire [111:0] nl_trt_loop_7_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  assign nl_trt_loop_7_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = {(chn_trt_in_rsci_d_mxwt[342:294])
      , 63'b0};
  wire [111:0] nl_trt_loop_8_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  assign nl_trt_loop_8_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = {(chn_trt_in_rsci_d_mxwt[391:343])
      , 63'b0};
  wire [111:0] nl_trt_loop_9_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  assign nl_trt_loop_9_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = {(chn_trt_in_rsci_d_mxwt[440:392])
      , 63'b0};
  wire [111:0] nl_trt_loop_10_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  assign nl_trt_loop_10_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = {(chn_trt_in_rsci_d_mxwt[489:441])
      , 63'b0};
  wire [111:0] nl_trt_loop_11_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  assign nl_trt_loop_11_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = {(chn_trt_in_rsci_d_mxwt[538:490])
      , 63'b0};
  wire [111:0] nl_trt_loop_12_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  assign nl_trt_loop_12_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = {(chn_trt_in_rsci_d_mxwt[587:539])
      , 63'b0};
  wire [111:0] nl_trt_loop_13_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  assign nl_trt_loop_13_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = {(chn_trt_in_rsci_d_mxwt[636:588])
      , 63'b0};
  wire [111:0] nl_trt_loop_14_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  assign nl_trt_loop_14_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = {(chn_trt_in_rsci_d_mxwt[685:637])
      , 63'b0};
  wire [111:0] nl_trt_loop_15_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  assign nl_trt_loop_15_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = {(chn_trt_in_rsci_d_mxwt[734:686])
      , 63'b0};
  wire [111:0] nl_trt_loop_16_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  assign nl_trt_loop_16_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = {(chn_trt_in_rsci_d_mxwt[783:735])
      , 63'b0};
  wire [511:0] nl_X_trt_core_chn_trt_out_rsci_inst_chn_trt_out_rsci_d;
  assign nl_X_trt_core_chn_trt_out_rsci_inst_chn_trt_out_rsci_d = {chn_trt_out_rsci_d_511
      , chn_trt_out_rsci_d_510_481 , chn_trt_out_rsci_d_480 , chn_trt_out_rsci_d_479
      , chn_trt_out_rsci_d_478_449 , chn_trt_out_rsci_d_448 , chn_trt_out_rsci_d_447
      , chn_trt_out_rsci_d_446_417 , chn_trt_out_rsci_d_416 , chn_trt_out_rsci_d_415
      , chn_trt_out_rsci_d_414_385 , chn_trt_out_rsci_d_384 , chn_trt_out_rsci_d_383
      , chn_trt_out_rsci_d_382_353 , chn_trt_out_rsci_d_352 , chn_trt_out_rsci_d_351
      , chn_trt_out_rsci_d_350_321 , chn_trt_out_rsci_d_320 , chn_trt_out_rsci_d_319
      , chn_trt_out_rsci_d_318_289 , chn_trt_out_rsci_d_288 , chn_trt_out_rsci_d_287
      , chn_trt_out_rsci_d_286_257 , chn_trt_out_rsci_d_256 , chn_trt_out_rsci_d_255
      , chn_trt_out_rsci_d_254_225 , chn_trt_out_rsci_d_224 , chn_trt_out_rsci_d_223
      , chn_trt_out_rsci_d_222_193 , chn_trt_out_rsci_d_192 , chn_trt_out_rsci_d_191
      , chn_trt_out_rsci_d_190_161 , chn_trt_out_rsci_d_160 , chn_trt_out_rsci_d_159
      , chn_trt_out_rsci_d_158_129 , chn_trt_out_rsci_d_128 , chn_trt_out_rsci_d_127
      , chn_trt_out_rsci_d_126_97 , chn_trt_out_rsci_d_96 , chn_trt_out_rsci_d_95
      , chn_trt_out_rsci_d_94_65 , chn_trt_out_rsci_d_64 , chn_trt_out_rsci_d_63
      , chn_trt_out_rsci_d_62_33 , chn_trt_out_rsci_d_32 , chn_trt_out_rsci_d_31
      , chn_trt_out_rsci_d_30_1 , chn_trt_out_rsci_d_0};
  SDP_X_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) trt_loop_1_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
      .a(nl_trt_loop_1_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a[111:0]),
      .s(cfg_mul_shift_value_rsci_d),
      .z(IntShiftRight_49U_6U_32U_mbits_fixed_1_sva)
    );
  SDP_X_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) trt_loop_2_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
      .a(nl_trt_loop_2_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a[111:0]),
      .s(cfg_mul_shift_value_rsci_d),
      .z(IntShiftRight_49U_6U_32U_mbits_fixed_2_sva)
    );
  SDP_X_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) trt_loop_3_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
      .a(nl_trt_loop_3_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a[111:0]),
      .s(cfg_mul_shift_value_rsci_d),
      .z(IntShiftRight_49U_6U_32U_mbits_fixed_3_sva)
    );
  SDP_X_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) trt_loop_4_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
      .a(nl_trt_loop_4_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a[111:0]),
      .s(cfg_mul_shift_value_rsci_d),
      .z(IntShiftRight_49U_6U_32U_mbits_fixed_4_sva)
    );
  SDP_X_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) trt_loop_5_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
      .a(nl_trt_loop_5_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a[111:0]),
      .s(cfg_mul_shift_value_rsci_d),
      .z(IntShiftRight_49U_6U_32U_mbits_fixed_5_sva)
    );
  SDP_X_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) trt_loop_6_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
      .a(nl_trt_loop_6_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a[111:0]),
      .s(cfg_mul_shift_value_rsci_d),
      .z(IntShiftRight_49U_6U_32U_mbits_fixed_6_sva)
    );
  SDP_X_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) trt_loop_7_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
      .a(nl_trt_loop_7_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a[111:0]),
      .s(cfg_mul_shift_value_rsci_d),
      .z(IntShiftRight_49U_6U_32U_mbits_fixed_7_sva)
    );
  SDP_X_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) trt_loop_8_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
      .a(nl_trt_loop_8_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a[111:0]),
      .s(cfg_mul_shift_value_rsci_d),
      .z(IntShiftRight_49U_6U_32U_mbits_fixed_8_sva)
    );
  SDP_X_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) trt_loop_9_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
      .a(nl_trt_loop_9_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a[111:0]),
      .s(cfg_mul_shift_value_rsci_d),
      .z(IntShiftRight_49U_6U_32U_mbits_fixed_9_sva)
    );
  SDP_X_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) trt_loop_10_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg
      (
      .a(nl_trt_loop_10_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a[111:0]),
      .s(cfg_mul_shift_value_rsci_d),
      .z(IntShiftRight_49U_6U_32U_mbits_fixed_10_sva)
    );
  SDP_X_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) trt_loop_11_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg
      (
      .a(nl_trt_loop_11_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a[111:0]),
      .s(cfg_mul_shift_value_rsci_d),
      .z(IntShiftRight_49U_6U_32U_mbits_fixed_11_sva)
    );
  SDP_X_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) trt_loop_12_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg
      (
      .a(nl_trt_loop_12_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a[111:0]),
      .s(cfg_mul_shift_value_rsci_d),
      .z(IntShiftRight_49U_6U_32U_mbits_fixed_12_sva)
    );
  SDP_X_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) trt_loop_13_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg
      (
      .a(nl_trt_loop_13_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a[111:0]),
      .s(cfg_mul_shift_value_rsci_d),
      .z(IntShiftRight_49U_6U_32U_mbits_fixed_13_sva)
    );
  SDP_X_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) trt_loop_14_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg
      (
      .a(nl_trt_loop_14_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a[111:0]),
      .s(cfg_mul_shift_value_rsci_d),
      .z(IntShiftRight_49U_6U_32U_mbits_fixed_14_sva)
    );
  SDP_X_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) trt_loop_15_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg
      (
      .a(nl_trt_loop_15_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a[111:0]),
      .s(cfg_mul_shift_value_rsci_d),
      .z(IntShiftRight_49U_6U_32U_mbits_fixed_15_sva)
    );
  SDP_X_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) trt_loop_16_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg
      (
      .a(nl_trt_loop_16_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a[111:0]),
      .s(cfg_mul_shift_value_rsci_d),
      .z(IntShiftRight_49U_6U_32U_mbits_fixed_sva)
    );
  SDP_X_X_trt_core_chn_trt_in_rsci X_trt_core_chn_trt_in_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_trt_in_rsc_slz(chn_trt_in_rsc_slz),
      .chn_trt_in_rsc_sz(chn_trt_in_rsc_sz),
      .chn_trt_in_rsc_z(chn_trt_in_rsc_z),
      .chn_trt_in_rsc_vz(chn_trt_in_rsc_vz),
      .chn_trt_in_rsc_lz(chn_trt_in_rsc_lz),
      .chn_trt_in_rsci_oswt(chn_trt_in_rsci_oswt),
      .core_wen(core_wen),
      .chn_trt_in_rsci_iswt0(chn_trt_in_rsci_iswt0),
      .chn_trt_in_rsci_bawt(chn_trt_in_rsci_bawt),
      .chn_trt_in_rsci_wen_comp(chn_trt_in_rsci_wen_comp),
      .chn_trt_in_rsci_ld_core_psct(chn_trt_in_rsci_ld_core_psct),
      .chn_trt_in_rsci_d_mxwt(chn_trt_in_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  SDP_X_X_trt_core_chn_trt_out_rsci X_trt_core_chn_trt_out_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_trt_out_rsc_z(chn_trt_out_rsc_z),
      .chn_trt_out_rsc_vz(chn_trt_out_rsc_vz),
      .chn_trt_out_rsc_lz(chn_trt_out_rsc_lz),
      .chn_trt_out_rsci_oswt(chn_trt_out_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_trt_out_rsci_iswt0(reg_cfg_mul_shift_value_rsc_triosy_obj_ld_core_psct_cse),
      .chn_trt_out_rsci_bawt(chn_trt_out_rsci_bawt),
      .chn_trt_out_rsci_wen_comp(chn_trt_out_rsci_wen_comp),
      .chn_trt_out_rsci_ld_core_psct(reg_chn_trt_out_rsci_ld_core_psct_cse),
      .chn_trt_out_rsci_d(nl_X_trt_core_chn_trt_out_rsci_inst_chn_trt_out_rsci_d[511:0])
    );
  SDP_X_X_trt_core_cfg_mul_shift_value_rsc_triosy_obj X_trt_core_cfg_mul_shift_value_rsc_triosy_obj_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_mul_shift_value_rsc_triosy_lz(cfg_mul_shift_value_rsc_triosy_lz),
      .cfg_mul_shift_value_rsc_triosy_obj_oswt(cfg_mul_shift_value_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_mul_shift_value_rsc_triosy_obj_iswt0(reg_cfg_mul_shift_value_rsc_triosy_obj_ld_core_psct_cse),
      .cfg_mul_shift_value_rsc_triosy_obj_bawt(cfg_mul_shift_value_rsc_triosy_obj_bawt)
    );
  SDP_X_X_trt_core_staller X_trt_core_staller_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .chn_trt_in_rsci_wen_comp(chn_trt_in_rsci_wen_comp),
      .core_wten(core_wten),
      .chn_trt_out_rsci_wen_comp(chn_trt_out_rsci_wen_comp)
    );
  SDP_X_X_trt_core_core_fsm X_trt_core_core_fsm_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign chn_trt_out_and_2_cse = core_wen & (and_148_cse | and_150_cse);
  assign trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[62])
      & ((IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[0]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[1])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[2]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[3])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[4]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[5])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[6]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[7])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[8]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[9])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[10]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[11])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[12]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[13])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[14]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[15])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[16]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[17])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[18]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[19])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[20]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[21])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[22]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[23])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[24]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[25])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[26]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[27])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[28]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[29])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[30]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[31])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[32]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[33])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[34]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[35])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[36]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[37])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[38]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[39])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[40]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[41])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[42]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[43])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[44]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[45])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[46]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[47])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[48]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[49])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[50]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[51])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[52]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[53])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[54]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[55])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[56]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[57])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[58]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[59])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[60]) | (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[61])
      | (~ (IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[111])));
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva = conv_s2s_49_50(IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[111:63])
      + conv_u2s_1_50(trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_and_nl);
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva = nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva[49:0];
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_1_sva = ~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva[49])
      | (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva[48:31]!=18'b000000000000000000))));
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_1_sva = (IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva[49])
      & (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva[48:31]==18'b111111111111111111)));
  assign trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[62])
      & ((IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[0]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[1])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[2]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[3])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[4]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[5])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[6]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[7])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[8]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[9])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[10]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[11])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[12]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[13])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[14]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[15])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[16]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[17])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[18]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[19])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[20]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[21])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[22]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[23])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[24]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[25])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[26]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[27])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[28]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[29])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[30]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[31])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[32]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[33])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[34]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[35])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[36]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[37])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[38]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[39])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[40]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[41])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[42]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[43])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[44]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[45])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[46]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[47])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[48]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[49])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[50]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[51])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[52]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[53])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[54]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[55])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[56]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[57])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[58]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[59])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[60]) | (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[61])
      | (~ (IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[111])));
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva = conv_s2s_49_50(IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[111:63])
      + conv_u2s_1_50(trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_and_nl);
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva = nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva[49:0];
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_2_sva = ~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva[49])
      | (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva[48:31]!=18'b000000000000000000))));
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_2_sva = (IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva[49])
      & (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva[48:31]==18'b111111111111111111)));
  assign trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[62])
      & ((IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[0]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[1])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[2]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[3])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[4]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[5])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[6]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[7])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[8]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[9])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[10]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[11])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[12]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[13])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[14]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[15])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[16]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[17])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[18]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[19])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[20]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[21])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[22]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[23])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[24]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[25])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[26]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[27])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[28]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[29])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[30]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[31])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[32]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[33])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[34]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[35])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[36]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[37])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[38]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[39])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[40]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[41])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[42]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[43])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[44]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[45])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[46]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[47])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[48]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[49])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[50]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[51])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[52]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[53])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[54]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[55])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[56]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[57])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[58]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[59])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[60]) | (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[61])
      | (~ (IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[111])));
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva = conv_s2s_49_50(IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[111:63])
      + conv_u2s_1_50(trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_and_nl);
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva = nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva[49:0];
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_3_sva = ~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva[49])
      | (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva[48:31]!=18'b000000000000000000))));
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_3_sva = (IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva[49])
      & (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva[48:31]==18'b111111111111111111)));
  assign trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[62])
      & ((IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[0]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[1])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[2]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[3])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[4]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[5])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[6]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[7])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[8]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[9])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[10]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[11])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[12]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[13])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[14]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[15])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[16]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[17])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[18]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[19])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[20]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[21])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[22]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[23])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[24]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[25])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[26]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[27])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[28]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[29])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[30]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[31])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[32]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[33])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[34]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[35])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[36]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[37])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[38]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[39])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[40]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[41])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[42]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[43])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[44]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[45])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[46]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[47])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[48]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[49])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[50]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[51])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[52]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[53])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[54]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[55])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[56]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[57])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[58]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[59])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[60]) | (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[61])
      | (~ (IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[111])));
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva = conv_s2s_49_50(IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[111:63])
      + conv_u2s_1_50(trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_and_nl);
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva = nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva[49:0];
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_4_sva = ~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva[49])
      | (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva[48:31]!=18'b000000000000000000))));
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_4_sva = (IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva[49])
      & (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva[48:31]==18'b111111111111111111)));
  assign trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[62])
      & ((IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[0]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[1])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[2]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[3])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[4]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[5])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[6]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[7])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[8]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[9])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[10]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[11])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[12]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[13])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[14]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[15])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[16]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[17])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[18]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[19])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[20]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[21])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[22]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[23])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[24]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[25])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[26]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[27])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[28]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[29])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[30]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[31])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[32]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[33])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[34]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[35])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[36]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[37])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[38]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[39])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[40]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[41])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[42]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[43])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[44]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[45])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[46]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[47])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[48]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[49])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[50]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[51])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[52]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[53])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[54]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[55])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[56]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[57])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[58]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[59])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[60]) | (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[61])
      | (~ (IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[111])));
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva = conv_s2s_49_50(IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[111:63])
      + conv_u2s_1_50(trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_and_nl);
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva = nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva[49:0];
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_5_sva = ~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva[49])
      | (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva[48:31]!=18'b000000000000000000))));
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_5_sva = (IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva[49])
      & (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva[48:31]==18'b111111111111111111)));
  assign trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[62])
      & ((IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[0]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[1])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[2]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[3])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[4]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[5])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[6]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[7])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[8]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[9])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[10]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[11])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[12]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[13])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[14]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[15])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[16]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[17])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[18]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[19])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[20]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[21])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[22]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[23])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[24]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[25])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[26]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[27])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[28]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[29])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[30]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[31])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[32]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[33])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[34]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[35])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[36]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[37])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[38]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[39])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[40]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[41])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[42]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[43])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[44]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[45])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[46]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[47])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[48]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[49])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[50]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[51])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[52]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[53])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[54]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[55])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[56]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[57])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[58]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[59])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[60]) | (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[61])
      | (~ (IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[111])));
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva = conv_s2s_49_50(IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[111:63])
      + conv_u2s_1_50(trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_and_nl);
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva = nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva[49:0];
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_6_sva = ~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva[49])
      | (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva[48:31]!=18'b000000000000000000))));
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_6_sva = (IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva[49])
      & (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva[48:31]==18'b111111111111111111)));
  assign trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[62])
      & ((IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[0]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[1])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[2]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[3])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[4]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[5])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[6]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[7])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[8]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[9])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[10]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[11])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[12]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[13])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[14]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[15])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[16]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[17])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[18]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[19])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[20]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[21])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[22]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[23])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[24]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[25])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[26]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[27])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[28]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[29])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[30]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[31])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[32]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[33])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[34]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[35])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[36]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[37])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[38]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[39])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[40]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[41])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[42]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[43])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[44]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[45])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[46]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[47])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[48]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[49])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[50]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[51])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[52]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[53])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[54]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[55])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[56]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[57])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[58]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[59])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[60]) | (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[61])
      | (~ (IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[111])));
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva = conv_s2s_49_50(IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[111:63])
      + conv_u2s_1_50(trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_and_nl);
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva = nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva[49:0];
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_7_sva = ~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva[49])
      | (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva[48:31]!=18'b000000000000000000))));
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_7_sva = (IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva[49])
      & (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva[48:31]==18'b111111111111111111)));
  assign trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[62])
      & ((IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[0]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[1])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[2]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[3])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[4]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[5])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[6]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[7])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[8]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[9])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[10]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[11])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[12]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[13])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[14]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[15])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[16]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[17])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[18]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[19])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[20]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[21])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[22]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[23])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[24]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[25])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[26]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[27])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[28]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[29])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[30]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[31])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[32]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[33])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[34]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[35])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[36]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[37])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[38]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[39])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[40]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[41])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[42]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[43])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[44]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[45])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[46]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[47])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[48]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[49])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[50]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[51])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[52]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[53])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[54]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[55])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[56]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[57])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[58]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[59])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[60]) | (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[61])
      | (~ (IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[111])));
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva = conv_s2s_49_50(IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[111:63])
      + conv_u2s_1_50(trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_and_nl);
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva = nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva[49:0];
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_8_sva = ~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva[49])
      | (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva[48:31]!=18'b000000000000000000))));
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_8_sva = (IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva[49])
      & (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva[48:31]==18'b111111111111111111)));
  assign trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[62])
      & ((IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[0]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[1])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[2]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[3])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[4]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[5])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[6]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[7])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[8]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[9])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[10]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[11])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[12]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[13])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[14]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[15])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[16]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[17])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[18]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[19])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[20]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[21])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[22]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[23])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[24]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[25])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[26]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[27])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[28]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[29])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[30]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[31])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[32]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[33])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[34]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[35])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[36]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[37])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[38]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[39])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[40]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[41])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[42]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[43])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[44]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[45])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[46]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[47])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[48]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[49])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[50]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[51])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[52]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[53])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[54]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[55])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[56]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[57])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[58]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[59])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[60]) | (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[61])
      | (~ (IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[111])));
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva = conv_s2s_49_50(IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[111:63])
      + conv_u2s_1_50(trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_and_nl);
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva = nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva[49:0];
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_9_sva = ~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva[49])
      | (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva[48:31]!=18'b000000000000000000))));
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_9_sva = (IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva[49])
      & (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva[48:31]==18'b111111111111111111)));
  assign trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[62])
      & ((IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[0]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[1])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[2]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[3])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[4]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[5])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[6]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[7])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[8]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[9])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[10]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[11])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[12]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[13])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[14]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[15])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[16]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[17])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[18]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[19])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[20]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[21])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[22]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[23])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[24]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[25])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[26]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[27])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[28]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[29])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[30]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[31])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[32]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[33])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[34]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[35])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[36]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[37])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[38]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[39])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[40]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[41])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[42]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[43])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[44]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[45])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[46]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[47])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[48]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[49])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[50]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[51])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[52]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[53])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[54]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[55])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[56]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[57])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[58]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[59])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[60]) | (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[61])
      | (~ (IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[111])));
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva = conv_s2s_49_50(IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[111:63])
      + conv_u2s_1_50(trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_and_nl);
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva = nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva[49:0];
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_10_sva = ~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva[49])
      | (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva[48:31]!=18'b000000000000000000))));
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_10_sva = (IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva[49])
      & (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva[48:31]==18'b111111111111111111)));
  assign trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[62])
      & ((IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[0]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[1])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[2]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[3])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[4]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[5])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[6]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[7])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[8]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[9])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[10]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[11])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[12]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[13])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[14]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[15])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[16]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[17])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[18]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[19])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[20]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[21])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[22]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[23])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[24]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[25])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[26]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[27])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[28]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[29])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[30]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[31])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[32]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[33])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[34]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[35])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[36]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[37])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[38]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[39])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[40]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[41])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[42]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[43])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[44]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[45])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[46]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[47])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[48]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[49])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[50]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[51])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[52]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[53])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[54]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[55])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[56]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[57])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[58]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[59])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[60]) | (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[61])
      | (~ (IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[111])));
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva = conv_s2s_49_50(IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[111:63])
      + conv_u2s_1_50(trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_and_nl);
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva = nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva[49:0];
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_11_sva = ~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva[49])
      | (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva[48:31]!=18'b000000000000000000))));
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_11_sva = (IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva[49])
      & (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva[48:31]==18'b111111111111111111)));
  assign trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[62])
      & ((IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[0]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[1])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[2]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[3])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[4]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[5])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[6]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[7])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[8]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[9])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[10]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[11])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[12]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[13])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[14]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[15])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[16]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[17])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[18]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[19])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[20]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[21])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[22]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[23])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[24]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[25])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[26]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[27])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[28]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[29])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[30]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[31])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[32]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[33])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[34]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[35])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[36]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[37])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[38]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[39])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[40]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[41])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[42]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[43])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[44]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[45])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[46]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[47])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[48]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[49])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[50]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[51])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[52]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[53])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[54]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[55])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[56]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[57])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[58]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[59])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[60]) | (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[61])
      | (~ (IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[111])));
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva = conv_s2s_49_50(IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[111:63])
      + conv_u2s_1_50(trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_and_nl);
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva = nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva[49:0];
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_12_sva = ~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva[49])
      | (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva[48:31]!=18'b000000000000000000))));
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_12_sva = (IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva[49])
      & (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva[48:31]==18'b111111111111111111)));
  assign trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[62])
      & ((IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[0]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[1])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[2]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[3])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[4]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[5])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[6]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[7])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[8]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[9])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[10]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[11])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[12]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[13])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[14]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[15])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[16]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[17])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[18]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[19])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[20]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[21])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[22]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[23])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[24]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[25])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[26]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[27])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[28]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[29])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[30]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[31])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[32]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[33])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[34]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[35])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[36]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[37])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[38]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[39])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[40]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[41])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[42]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[43])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[44]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[45])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[46]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[47])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[48]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[49])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[50]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[51])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[52]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[53])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[54]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[55])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[56]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[57])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[58]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[59])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[60]) | (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[61])
      | (~ (IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[111])));
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva = conv_s2s_49_50(IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[111:63])
      + conv_u2s_1_50(trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_and_nl);
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva = nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva[49:0];
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_13_sva = ~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva[49])
      | (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva[48:31]!=18'b000000000000000000))));
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_13_sva = (IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva[49])
      & (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva[48:31]==18'b111111111111111111)));
  assign trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[62])
      & ((IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[0]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[1])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[2]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[3])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[4]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[5])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[6]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[7])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[8]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[9])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[10]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[11])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[12]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[13])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[14]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[15])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[16]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[17])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[18]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[19])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[20]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[21])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[22]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[23])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[24]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[25])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[26]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[27])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[28]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[29])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[30]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[31])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[32]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[33])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[34]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[35])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[36]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[37])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[38]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[39])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[40]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[41])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[42]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[43])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[44]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[45])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[46]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[47])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[48]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[49])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[50]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[51])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[52]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[53])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[54]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[55])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[56]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[57])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[58]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[59])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[60]) | (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[61])
      | (~ (IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[111])));
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva = conv_s2s_49_50(IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[111:63])
      + conv_u2s_1_50(trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_and_nl);
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva = nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva[49:0];
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_14_sva = ~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva[49])
      | (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva[48:31]!=18'b000000000000000000))));
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_14_sva = (IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva[49])
      & (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva[48:31]==18'b111111111111111111)));
  assign trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[62])
      & ((IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[0]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[1])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[2]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[3])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[4]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[5])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[6]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[7])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[8]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[9])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[10]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[11])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[12]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[13])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[14]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[15])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[16]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[17])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[18]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[19])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[20]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[21])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[22]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[23])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[24]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[25])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[26]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[27])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[28]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[29])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[30]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[31])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[32]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[33])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[34]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[35])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[36]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[37])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[38]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[39])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[40]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[41])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[42]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[43])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[44]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[45])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[46]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[47])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[48]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[49])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[50]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[51])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[52]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[53])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[54]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[55])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[56]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[57])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[58]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[59])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[60]) | (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[61])
      | (~ (IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[111])));
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva = conv_s2s_49_50(IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[111:63])
      + conv_u2s_1_50(trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_and_nl);
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva = nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva[49:0];
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_15_sva = ~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva[49])
      | (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva[48:31]!=18'b000000000000000000))));
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_15_sva = (IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva[49])
      & (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva[48:31]==18'b111111111111111111)));
  assign trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = (IntShiftRight_49U_6U_32U_mbits_fixed_sva[62])
      & ((IntShiftRight_49U_6U_32U_mbits_fixed_sva[0]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[1])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[2]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[3])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[4]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[5])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[6]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[7])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[8]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[9])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[10]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[11])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[12]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[13])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[14]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[15])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[16]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[17])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[18]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[19])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[20]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[21])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[22]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[23])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[24]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[25])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[26]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[27])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[28]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[29])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[30]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[31])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[32]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[33])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[34]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[35])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[36]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[37])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[38]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[39])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[40]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[41])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[42]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[43])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[44]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[45])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[46]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[47])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[48]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[49])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[50]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[51])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[52]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[53])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[54]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[55])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[56]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[57])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[58]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[59])
      | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[60]) | (IntShiftRight_49U_6U_32U_mbits_fixed_sva[61])
      | (~ (IntShiftRight_49U_6U_32U_mbits_fixed_sva[111])));
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva = conv_s2s_49_50(IntShiftRight_49U_6U_32U_mbits_fixed_sva[111:63])
      + conv_u2s_1_50(trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_and_nl);
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva = nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva[49:0];
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_sva = ~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva[49])
      | (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva[48:31]!=18'b000000000000000000))));
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_sva = (IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva[49])
      & (~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva[48:31]==18'b111111111111111111)));
  assign and_4_mdf = chn_trt_in_rsci_bawt & (chn_trt_out_rsci_bawt | (~ reg_chn_trt_out_rsci_ld_core_psct_cse))
      & (cfg_mul_shift_value_rsc_triosy_obj_bawt | (~ reg_chn_trt_out_rsci_ld_core_psct_cse));
  assign and_dcpl_1 = chn_trt_out_rsci_bawt & cfg_mul_shift_value_rsc_triosy_obj_bawt;
  assign or_dcpl = and_dcpl_1 | (~ reg_chn_trt_out_rsci_ld_core_psct_cse);
  assign and_dcpl_3 = and_dcpl_1 & reg_chn_trt_out_rsci_ld_core_psct_cse;
  assign or_dcpl_3 = (cfg_precision!=2'b10);
  assign and_dcpl_7 = or_dcpl_3 & chn_trt_in_rsci_bawt;
  assign and_dcpl_11 = chn_trt_in_rsci_bawt & (cfg_precision==2'b10);
  assign and_dcpl_15 = or_dcpl & or_dcpl_3;
  assign and_dcpl_17 = reg_chn_trt_out_rsci_ld_core_psct_cse & chn_trt_in_rsci_bawt;
  assign and_dcpl_19 = and_dcpl_1 & or_dcpl_3;
  assign not_tmp_9 = ~((cfg_precision[0]) | (~((cfg_precision[1]) & or_dcpl)));
  assign and_dcpl_23 = cfg_mul_shift_value_rsc_triosy_obj_bawt & reg_chn_trt_out_rsci_ld_core_psct_cse
      & chn_trt_in_rsci_bawt;
  assign and_dcpl_24 = (cfg_precision==2'b10);
  assign and_dcpl_134 = and_dcpl_1 & reg_chn_trt_out_rsci_ld_core_psct_cse & (~ chn_trt_in_rsci_bawt);
  assign and_148_cse = or_dcpl & and_dcpl_7 & (fsm_output[1]);
  assign and_150_cse = or_dcpl & and_dcpl_11 & (fsm_output[1]);
  assign or_tmp_150 = or_dcpl & chn_trt_in_rsci_bawt & (fsm_output[1]);
  assign chn_trt_in_rsci_ld_core_psct_mx0c0 = and_4_mdf | (fsm_output[0]);
  assign chn_trt_out_rsci_d_0_mx0c1 = and_150_cse | (and_dcpl_3 & and_dcpl_11);
  assign mux_4_nl = MUX_s_1_2_2(not_tmp_9, or_dcpl, chn_trt_in_rsci_d_mxwt[784]);
  assign chn_trt_out_rsci_d_30_1_mx0c1 = ((mux_4_nl) & chn_trt_in_rsci_bawt & (fsm_output[1]))
      | ((and_dcpl_24 | (chn_trt_in_rsci_d_mxwt[784])) & chn_trt_out_rsci_bawt &
      and_dcpl_23);
  assign mux_5_nl = MUX_s_1_2_2(not_tmp_9, or_dcpl, chn_trt_in_rsci_d_mxwt[785]);
  assign chn_trt_out_rsci_d_62_33_mx0c1 = ((mux_5_nl) & chn_trt_in_rsci_bawt & (fsm_output[1]))
      | ((and_dcpl_24 | (chn_trt_in_rsci_d_mxwt[785])) & chn_trt_out_rsci_bawt &
      and_dcpl_23);
  assign mux_6_nl = MUX_s_1_2_2(not_tmp_9, or_dcpl, chn_trt_in_rsci_d_mxwt[786]);
  assign chn_trt_out_rsci_d_94_65_mx0c1 = ((mux_6_nl) & chn_trt_in_rsci_bawt & (fsm_output[1]))
      | ((and_dcpl_24 | (chn_trt_in_rsci_d_mxwt[786])) & chn_trt_out_rsci_bawt &
      and_dcpl_23);
  assign mux_7_nl = MUX_s_1_2_2(not_tmp_9, or_dcpl, chn_trt_in_rsci_d_mxwt[787]);
  assign chn_trt_out_rsci_d_126_97_mx0c1 = ((mux_7_nl) & chn_trt_in_rsci_bawt & (fsm_output[1]))
      | ((and_dcpl_24 | (chn_trt_in_rsci_d_mxwt[787])) & chn_trt_out_rsci_bawt &
      and_dcpl_23);
  assign mux_8_nl = MUX_s_1_2_2(not_tmp_9, or_dcpl, chn_trt_in_rsci_d_mxwt[788]);
  assign chn_trt_out_rsci_d_158_129_mx0c1 = ((mux_8_nl) & chn_trt_in_rsci_bawt &
      (fsm_output[1])) | ((and_dcpl_24 | (chn_trt_in_rsci_d_mxwt[788])) & chn_trt_out_rsci_bawt
      & and_dcpl_23);
  assign mux_9_nl = MUX_s_1_2_2(not_tmp_9, or_dcpl, chn_trt_in_rsci_d_mxwt[789]);
  assign chn_trt_out_rsci_d_190_161_mx0c1 = ((mux_9_nl) & chn_trt_in_rsci_bawt &
      (fsm_output[1])) | ((and_dcpl_24 | (chn_trt_in_rsci_d_mxwt[789])) & chn_trt_out_rsci_bawt
      & and_dcpl_23);
  assign mux_10_nl = MUX_s_1_2_2(not_tmp_9, or_dcpl, chn_trt_in_rsci_d_mxwt[790]);
  assign chn_trt_out_rsci_d_222_193_mx0c1 = ((mux_10_nl) & chn_trt_in_rsci_bawt &
      (fsm_output[1])) | ((and_dcpl_24 | (chn_trt_in_rsci_d_mxwt[790])) & chn_trt_out_rsci_bawt
      & and_dcpl_23);
  assign mux_11_nl = MUX_s_1_2_2(not_tmp_9, or_dcpl, chn_trt_in_rsci_d_mxwt[791]);
  assign chn_trt_out_rsci_d_254_225_mx0c1 = ((mux_11_nl) & chn_trt_in_rsci_bawt &
      (fsm_output[1])) | ((and_dcpl_24 | (chn_trt_in_rsci_d_mxwt[791])) & chn_trt_out_rsci_bawt
      & and_dcpl_23);
  assign mux_12_nl = MUX_s_1_2_2(not_tmp_9, or_dcpl, chn_trt_in_rsci_d_mxwt[792]);
  assign chn_trt_out_rsci_d_286_257_mx0c1 = ((mux_12_nl) & chn_trt_in_rsci_bawt &
      (fsm_output[1])) | ((and_dcpl_24 | (chn_trt_in_rsci_d_mxwt[792])) & chn_trt_out_rsci_bawt
      & and_dcpl_23);
  assign mux_13_nl = MUX_s_1_2_2(not_tmp_9, or_dcpl, chn_trt_in_rsci_d_mxwt[793]);
  assign chn_trt_out_rsci_d_318_289_mx0c1 = ((mux_13_nl) & chn_trt_in_rsci_bawt &
      (fsm_output[1])) | ((and_dcpl_24 | (chn_trt_in_rsci_d_mxwt[793])) & chn_trt_out_rsci_bawt
      & and_dcpl_23);
  assign mux_14_nl = MUX_s_1_2_2(not_tmp_9, or_dcpl, chn_trt_in_rsci_d_mxwt[794]);
  assign chn_trt_out_rsci_d_350_321_mx0c1 = ((mux_14_nl) & chn_trt_in_rsci_bawt &
      (fsm_output[1])) | ((and_dcpl_24 | (chn_trt_in_rsci_d_mxwt[794])) & chn_trt_out_rsci_bawt
      & and_dcpl_23);
  assign mux_15_nl = MUX_s_1_2_2(not_tmp_9, or_dcpl, chn_trt_in_rsci_d_mxwt[795]);
  assign chn_trt_out_rsci_d_382_353_mx0c1 = ((mux_15_nl) & chn_trt_in_rsci_bawt &
      (fsm_output[1])) | ((and_dcpl_24 | (chn_trt_in_rsci_d_mxwt[795])) & chn_trt_out_rsci_bawt
      & and_dcpl_23);
  assign mux_16_nl = MUX_s_1_2_2(not_tmp_9, or_dcpl, chn_trt_in_rsci_d_mxwt[796]);
  assign chn_trt_out_rsci_d_414_385_mx0c1 = ((mux_16_nl) & chn_trt_in_rsci_bawt &
      (fsm_output[1])) | ((and_dcpl_24 | (chn_trt_in_rsci_d_mxwt[796])) & chn_trt_out_rsci_bawt
      & and_dcpl_23);
  assign mux_17_nl = MUX_s_1_2_2(not_tmp_9, or_dcpl, chn_trt_in_rsci_d_mxwt[797]);
  assign chn_trt_out_rsci_d_446_417_mx0c1 = ((mux_17_nl) & chn_trt_in_rsci_bawt &
      (fsm_output[1])) | ((and_dcpl_24 | (chn_trt_in_rsci_d_mxwt[797])) & chn_trt_out_rsci_bawt
      & and_dcpl_23);
  assign mux_18_nl = MUX_s_1_2_2(not_tmp_9, or_dcpl, chn_trt_in_rsci_d_mxwt[798]);
  assign chn_trt_out_rsci_d_478_449_mx0c1 = ((mux_18_nl) & chn_trt_in_rsci_bawt &
      (fsm_output[1])) | ((and_dcpl_24 | (chn_trt_in_rsci_d_mxwt[798])) & chn_trt_out_rsci_bawt
      & and_dcpl_23);
  assign mux_19_nl = MUX_s_1_2_2(not_tmp_9, or_dcpl, chn_trt_in_rsci_d_mxwt[799]);
  assign chn_trt_out_rsci_d_510_481_mx0c1 = ((mux_19_nl) & chn_trt_in_rsci_bawt &
      (fsm_output[1])) | ((and_dcpl_24 | (chn_trt_in_rsci_d_mxwt[799])) & chn_trt_out_rsci_bawt
      & and_dcpl_23);
  assign chn_trt_in_rsci_oswt_unreg = or_tmp_150;
  assign chn_trt_out_rsci_oswt_unreg_pff = and_dcpl_3;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_in_rsci_iswt0 <= 1'b0;
      reg_cfg_mul_shift_value_rsc_triosy_obj_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen ) begin
      chn_trt_in_rsci_iswt0 <= ~((~ and_4_mdf) & (fsm_output[1]));
      reg_cfg_mul_shift_value_rsc_triosy_obj_ld_core_psct_cse <= or_tmp_150;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_in_rsci_ld_core_psct <= 1'b0;
    end
    else if ( core_wen & chn_trt_in_rsci_ld_core_psct_mx0c0 ) begin
      chn_trt_in_rsci_ld_core_psct <= chn_trt_in_rsci_ld_core_psct_mx0c0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_out_rsci_d_0 <= 1'b0;
    end
    else if ( core_wen & (and_148_cse | (and_dcpl_3 & and_dcpl_7) | chn_trt_out_rsci_d_0_mx0c1)
        ) begin
      chn_trt_out_rsci_d_0 <= MUX_s_1_2_2((trt_loop_else_mux_112_nl), (chn_trt_in_rsci_d_mxwt[0]),
          chn_trt_out_rsci_d_0_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_out_rsci_d_30_1 <= 30'b0;
    end
    else if ( core_wen & ((and_dcpl_15 & chn_trt_in_rsci_bawt & (~ (chn_trt_in_rsci_d_mxwt[784]))
        & (fsm_output[1])) | (and_dcpl_19 & and_dcpl_17 & (~ (chn_trt_in_rsci_d_mxwt[784])))
        | chn_trt_out_rsci_d_30_1_mx0c1) ) begin
      chn_trt_out_rsci_d_30_1 <= MUX_v_30_2_2((trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl),
          (chn_trt_in_rsci_d_mxwt[30:1]), chn_trt_out_rsci_d_30_1_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_out_rsci_d_31 <= 1'b0;
      chn_trt_out_rsci_d_32 <= 1'b0;
      chn_trt_out_rsci_d_63 <= 1'b0;
      chn_trt_out_rsci_d_64 <= 1'b0;
      chn_trt_out_rsci_d_95 <= 1'b0;
      chn_trt_out_rsci_d_96 <= 1'b0;
      chn_trt_out_rsci_d_127 <= 1'b0;
      chn_trt_out_rsci_d_128 <= 1'b0;
      chn_trt_out_rsci_d_159 <= 1'b0;
      chn_trt_out_rsci_d_160 <= 1'b0;
      chn_trt_out_rsci_d_191 <= 1'b0;
      chn_trt_out_rsci_d_192 <= 1'b0;
      chn_trt_out_rsci_d_223 <= 1'b0;
      chn_trt_out_rsci_d_224 <= 1'b0;
      chn_trt_out_rsci_d_255 <= 1'b0;
      chn_trt_out_rsci_d_256 <= 1'b0;
      chn_trt_out_rsci_d_287 <= 1'b0;
      chn_trt_out_rsci_d_288 <= 1'b0;
      chn_trt_out_rsci_d_319 <= 1'b0;
      chn_trt_out_rsci_d_320 <= 1'b0;
      chn_trt_out_rsci_d_351 <= 1'b0;
      chn_trt_out_rsci_d_352 <= 1'b0;
      chn_trt_out_rsci_d_383 <= 1'b0;
      chn_trt_out_rsci_d_384 <= 1'b0;
      chn_trt_out_rsci_d_415 <= 1'b0;
      chn_trt_out_rsci_d_416 <= 1'b0;
      chn_trt_out_rsci_d_447 <= 1'b0;
      chn_trt_out_rsci_d_448 <= 1'b0;
      chn_trt_out_rsci_d_479 <= 1'b0;
      chn_trt_out_rsci_d_480 <= 1'b0;
      chn_trt_out_rsci_d_511 <= 1'b0;
    end
    else if ( chn_trt_out_and_2_cse ) begin
      chn_trt_out_rsci_d_31 <= MUX_s_1_2_2((trt_loop_else_mux_113_nl), (chn_trt_in_rsci_d_mxwt[31]),
          and_150_cse);
      chn_trt_out_rsci_d_32 <= MUX_s_1_2_2((trt_loop_else_mux_114_nl), (chn_trt_in_rsci_d_mxwt[49]),
          and_150_cse);
      chn_trt_out_rsci_d_63 <= MUX_s_1_2_2((trt_loop_else_mux_115_nl), (chn_trt_in_rsci_d_mxwt[80]),
          and_150_cse);
      chn_trt_out_rsci_d_64 <= MUX_s_1_2_2((trt_loop_else_mux_116_nl), (chn_trt_in_rsci_d_mxwt[98]),
          and_150_cse);
      chn_trt_out_rsci_d_95 <= MUX_s_1_2_2((trt_loop_else_mux_117_nl), (chn_trt_in_rsci_d_mxwt[129]),
          and_150_cse);
      chn_trt_out_rsci_d_96 <= MUX_s_1_2_2((trt_loop_else_mux_118_nl), (chn_trt_in_rsci_d_mxwt[147]),
          and_150_cse);
      chn_trt_out_rsci_d_127 <= MUX_s_1_2_2((trt_loop_else_mux_119_nl), (chn_trt_in_rsci_d_mxwt[178]),
          and_150_cse);
      chn_trt_out_rsci_d_128 <= MUX_s_1_2_2((trt_loop_else_mux_120_nl), (chn_trt_in_rsci_d_mxwt[196]),
          and_150_cse);
      chn_trt_out_rsci_d_159 <= MUX_s_1_2_2((trt_loop_else_mux_121_nl), (chn_trt_in_rsci_d_mxwt[227]),
          and_150_cse);
      chn_trt_out_rsci_d_160 <= MUX_s_1_2_2((trt_loop_else_mux_122_nl), (chn_trt_in_rsci_d_mxwt[245]),
          and_150_cse);
      chn_trt_out_rsci_d_191 <= MUX_s_1_2_2((trt_loop_else_mux_123_nl), (chn_trt_in_rsci_d_mxwt[276]),
          and_150_cse);
      chn_trt_out_rsci_d_192 <= MUX_s_1_2_2((trt_loop_else_mux_124_nl), (chn_trt_in_rsci_d_mxwt[294]),
          and_150_cse);
      chn_trt_out_rsci_d_223 <= MUX_s_1_2_2((trt_loop_else_mux_125_nl), (chn_trt_in_rsci_d_mxwt[325]),
          and_150_cse);
      chn_trt_out_rsci_d_224 <= MUX_s_1_2_2((trt_loop_else_mux_126_nl), (chn_trt_in_rsci_d_mxwt[343]),
          and_150_cse);
      chn_trt_out_rsci_d_255 <= MUX_s_1_2_2((trt_loop_else_mux_127_nl), (chn_trt_in_rsci_d_mxwt[374]),
          and_150_cse);
      chn_trt_out_rsci_d_256 <= MUX_s_1_2_2((trt_loop_else_mux_128_nl), (chn_trt_in_rsci_d_mxwt[392]),
          and_150_cse);
      chn_trt_out_rsci_d_287 <= MUX_s_1_2_2((trt_loop_else_mux_129_nl), (chn_trt_in_rsci_d_mxwt[423]),
          and_150_cse);
      chn_trt_out_rsci_d_288 <= MUX_s_1_2_2((trt_loop_else_mux_130_nl), (chn_trt_in_rsci_d_mxwt[441]),
          and_150_cse);
      chn_trt_out_rsci_d_319 <= MUX_s_1_2_2((trt_loop_else_mux_131_nl), (chn_trt_in_rsci_d_mxwt[472]),
          and_150_cse);
      chn_trt_out_rsci_d_320 <= MUX_s_1_2_2((trt_loop_else_mux_132_nl), (chn_trt_in_rsci_d_mxwt[490]),
          and_150_cse);
      chn_trt_out_rsci_d_351 <= MUX_s_1_2_2((trt_loop_else_mux_133_nl), (chn_trt_in_rsci_d_mxwt[521]),
          and_150_cse);
      chn_trt_out_rsci_d_352 <= MUX_s_1_2_2((trt_loop_else_mux_134_nl), (chn_trt_in_rsci_d_mxwt[539]),
          and_150_cse);
      chn_trt_out_rsci_d_383 <= MUX_s_1_2_2((trt_loop_else_mux_135_nl), (chn_trt_in_rsci_d_mxwt[570]),
          and_150_cse);
      chn_trt_out_rsci_d_384 <= MUX_s_1_2_2((trt_loop_else_mux_136_nl), (chn_trt_in_rsci_d_mxwt[588]),
          and_150_cse);
      chn_trt_out_rsci_d_415 <= MUX_s_1_2_2((trt_loop_else_mux_137_nl), (chn_trt_in_rsci_d_mxwt[619]),
          and_150_cse);
      chn_trt_out_rsci_d_416 <= MUX_s_1_2_2((trt_loop_else_mux_138_nl), (chn_trt_in_rsci_d_mxwt[637]),
          and_150_cse);
      chn_trt_out_rsci_d_447 <= MUX_s_1_2_2((trt_loop_else_mux_139_nl), (chn_trt_in_rsci_d_mxwt[668]),
          and_150_cse);
      chn_trt_out_rsci_d_448 <= MUX_s_1_2_2((trt_loop_else_mux_140_nl), (chn_trt_in_rsci_d_mxwt[686]),
          and_150_cse);
      chn_trt_out_rsci_d_479 <= MUX_s_1_2_2((trt_loop_else_mux_141_nl), (chn_trt_in_rsci_d_mxwt[717]),
          and_150_cse);
      chn_trt_out_rsci_d_480 <= MUX_s_1_2_2((trt_loop_else_mux_142_nl), (chn_trt_in_rsci_d_mxwt[735]),
          and_150_cse);
      chn_trt_out_rsci_d_511 <= MUX_s_1_2_2((trt_loop_else_mux_143_nl), (chn_trt_in_rsci_d_mxwt[766]),
          and_150_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_out_rsci_d_62_33 <= 30'b0;
    end
    else if ( core_wen & ((and_dcpl_15 & chn_trt_in_rsci_bawt & (~ (chn_trt_in_rsci_d_mxwt[785]))
        & (fsm_output[1])) | (and_dcpl_19 & and_dcpl_17 & (~ (chn_trt_in_rsci_d_mxwt[785])))
        | chn_trt_out_rsci_d_62_33_mx0c1) ) begin
      chn_trt_out_rsci_d_62_33 <= MUX_v_30_2_2((trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl),
          (chn_trt_in_rsci_d_mxwt[79:50]), chn_trt_out_rsci_d_62_33_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_out_rsci_d_94_65 <= 30'b0;
    end
    else if ( core_wen & ((and_dcpl_15 & chn_trt_in_rsci_bawt & (~ (chn_trt_in_rsci_d_mxwt[786]))
        & (fsm_output[1])) | (and_dcpl_19 & and_dcpl_17 & (~ (chn_trt_in_rsci_d_mxwt[786])))
        | chn_trt_out_rsci_d_94_65_mx0c1) ) begin
      chn_trt_out_rsci_d_94_65 <= MUX_v_30_2_2((trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl),
          (chn_trt_in_rsci_d_mxwt[128:99]), chn_trt_out_rsci_d_94_65_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_out_rsci_d_126_97 <= 30'b0;
    end
    else if ( core_wen & ((and_dcpl_15 & chn_trt_in_rsci_bawt & (~ (chn_trt_in_rsci_d_mxwt[787]))
        & (fsm_output[1])) | (and_dcpl_19 & and_dcpl_17 & (~ (chn_trt_in_rsci_d_mxwt[787])))
        | chn_trt_out_rsci_d_126_97_mx0c1) ) begin
      chn_trt_out_rsci_d_126_97 <= MUX_v_30_2_2((trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl),
          (chn_trt_in_rsci_d_mxwt[177:148]), chn_trt_out_rsci_d_126_97_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_out_rsci_d_158_129 <= 30'b0;
    end
    else if ( core_wen & ((and_dcpl_15 & chn_trt_in_rsci_bawt & (~ (chn_trt_in_rsci_d_mxwt[788]))
        & (fsm_output[1])) | (and_dcpl_19 & and_dcpl_17 & (~ (chn_trt_in_rsci_d_mxwt[788])))
        | chn_trt_out_rsci_d_158_129_mx0c1) ) begin
      chn_trt_out_rsci_d_158_129 <= MUX_v_30_2_2((trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl),
          (chn_trt_in_rsci_d_mxwt[226:197]), chn_trt_out_rsci_d_158_129_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_out_rsci_d_190_161 <= 30'b0;
    end
    else if ( core_wen & ((and_dcpl_15 & chn_trt_in_rsci_bawt & (~ (chn_trt_in_rsci_d_mxwt[789]))
        & (fsm_output[1])) | (and_dcpl_19 & and_dcpl_17 & (~ (chn_trt_in_rsci_d_mxwt[789])))
        | chn_trt_out_rsci_d_190_161_mx0c1) ) begin
      chn_trt_out_rsci_d_190_161 <= MUX_v_30_2_2((trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl),
          (chn_trt_in_rsci_d_mxwt[275:246]), chn_trt_out_rsci_d_190_161_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_out_rsci_d_222_193 <= 30'b0;
    end
    else if ( core_wen & ((and_dcpl_15 & chn_trt_in_rsci_bawt & (~ (chn_trt_in_rsci_d_mxwt[790]))
        & (fsm_output[1])) | (and_dcpl_19 & and_dcpl_17 & (~ (chn_trt_in_rsci_d_mxwt[790])))
        | chn_trt_out_rsci_d_222_193_mx0c1) ) begin
      chn_trt_out_rsci_d_222_193 <= MUX_v_30_2_2((trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl),
          (chn_trt_in_rsci_d_mxwt[324:295]), chn_trt_out_rsci_d_222_193_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_out_rsci_d_254_225 <= 30'b0;
    end
    else if ( core_wen & ((and_dcpl_15 & chn_trt_in_rsci_bawt & (~ (chn_trt_in_rsci_d_mxwt[791]))
        & (fsm_output[1])) | (and_dcpl_19 & and_dcpl_17 & (~ (chn_trt_in_rsci_d_mxwt[791])))
        | chn_trt_out_rsci_d_254_225_mx0c1) ) begin
      chn_trt_out_rsci_d_254_225 <= MUX_v_30_2_2((trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl),
          (chn_trt_in_rsci_d_mxwt[373:344]), chn_trt_out_rsci_d_254_225_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_out_rsci_d_286_257 <= 30'b0;
    end
    else if ( core_wen & ((and_dcpl_15 & chn_trt_in_rsci_bawt & (~ (chn_trt_in_rsci_d_mxwt[792]))
        & (fsm_output[1])) | (and_dcpl_19 & and_dcpl_17 & (~ (chn_trt_in_rsci_d_mxwt[792])))
        | chn_trt_out_rsci_d_286_257_mx0c1) ) begin
      chn_trt_out_rsci_d_286_257 <= MUX_v_30_2_2((trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl),
          (chn_trt_in_rsci_d_mxwt[422:393]), chn_trt_out_rsci_d_286_257_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_out_rsci_d_318_289 <= 30'b0;
    end
    else if ( core_wen & ((and_dcpl_15 & chn_trt_in_rsci_bawt & (~ (chn_trt_in_rsci_d_mxwt[793]))
        & (fsm_output[1])) | (and_dcpl_19 & and_dcpl_17 & (~ (chn_trt_in_rsci_d_mxwt[793])))
        | chn_trt_out_rsci_d_318_289_mx0c1) ) begin
      chn_trt_out_rsci_d_318_289 <= MUX_v_30_2_2((trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl),
          (chn_trt_in_rsci_d_mxwt[471:442]), chn_trt_out_rsci_d_318_289_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_out_rsci_d_350_321 <= 30'b0;
    end
    else if ( core_wen & ((and_dcpl_15 & chn_trt_in_rsci_bawt & (~ (chn_trt_in_rsci_d_mxwt[794]))
        & (fsm_output[1])) | (and_dcpl_19 & and_dcpl_17 & (~ (chn_trt_in_rsci_d_mxwt[794])))
        | chn_trt_out_rsci_d_350_321_mx0c1) ) begin
      chn_trt_out_rsci_d_350_321 <= MUX_v_30_2_2((trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl),
          (chn_trt_in_rsci_d_mxwt[520:491]), chn_trt_out_rsci_d_350_321_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_out_rsci_d_382_353 <= 30'b0;
    end
    else if ( core_wen & ((and_dcpl_15 & chn_trt_in_rsci_bawt & (~ (chn_trt_in_rsci_d_mxwt[795]))
        & (fsm_output[1])) | (and_dcpl_19 & and_dcpl_17 & (~ (chn_trt_in_rsci_d_mxwt[795])))
        | chn_trt_out_rsci_d_382_353_mx0c1) ) begin
      chn_trt_out_rsci_d_382_353 <= MUX_v_30_2_2((trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl),
          (chn_trt_in_rsci_d_mxwt[569:540]), chn_trt_out_rsci_d_382_353_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_out_rsci_d_414_385 <= 30'b0;
    end
    else if ( core_wen & ((and_dcpl_15 & chn_trt_in_rsci_bawt & (~ (chn_trt_in_rsci_d_mxwt[796]))
        & (fsm_output[1])) | (and_dcpl_19 & and_dcpl_17 & (~ (chn_trt_in_rsci_d_mxwt[796])))
        | chn_trt_out_rsci_d_414_385_mx0c1) ) begin
      chn_trt_out_rsci_d_414_385 <= MUX_v_30_2_2((trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl),
          (chn_trt_in_rsci_d_mxwt[618:589]), chn_trt_out_rsci_d_414_385_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_out_rsci_d_446_417 <= 30'b0;
    end
    else if ( core_wen & ((and_dcpl_15 & chn_trt_in_rsci_bawt & (~ (chn_trt_in_rsci_d_mxwt[797]))
        & (fsm_output[1])) | (and_dcpl_19 & and_dcpl_17 & (~ (chn_trt_in_rsci_d_mxwt[797])))
        | chn_trt_out_rsci_d_446_417_mx0c1) ) begin
      chn_trt_out_rsci_d_446_417 <= MUX_v_30_2_2((trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl),
          (chn_trt_in_rsci_d_mxwt[667:638]), chn_trt_out_rsci_d_446_417_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_out_rsci_d_478_449 <= 30'b0;
    end
    else if ( core_wen & ((and_dcpl_15 & chn_trt_in_rsci_bawt & (~ (chn_trt_in_rsci_d_mxwt[798]))
        & (fsm_output[1])) | (and_dcpl_19 & and_dcpl_17 & (~ (chn_trt_in_rsci_d_mxwt[798])))
        | chn_trt_out_rsci_d_478_449_mx0c1) ) begin
      chn_trt_out_rsci_d_478_449 <= MUX_v_30_2_2((trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl),
          (chn_trt_in_rsci_d_mxwt[716:687]), chn_trt_out_rsci_d_478_449_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_trt_out_rsci_d_510_481 <= 30'b0;
    end
    else if ( core_wen & ((and_dcpl_15 & chn_trt_in_rsci_bawt & (~ (chn_trt_in_rsci_d_mxwt[799]))
        & (fsm_output[1])) | (and_dcpl_19 & and_dcpl_17 & (~ (chn_trt_in_rsci_d_mxwt[799])))
        | chn_trt_out_rsci_d_510_481_mx0c1) ) begin
      chn_trt_out_rsci_d_510_481 <= MUX_v_30_2_2((trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl),
          (chn_trt_in_rsci_d_mxwt[765:736]), chn_trt_out_rsci_d_510_481_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_trt_out_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (or_tmp_150 | and_dcpl_134) ) begin
      reg_chn_trt_out_rsci_ld_core_psct_cse <= ~ and_dcpl_134;
    end
  end
  assign trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva[0]) | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_1_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_1_sva);
  assign trt_loop_else_mux_112_nl = MUX_s_1_2_2((trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl),
      (chn_trt_in_rsci_d_mxwt[0]), chn_trt_in_rsci_d_mxwt[784]);
  assign trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_1_sva));
  assign trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl
      = ~(MUX_v_30_2_2((trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_1_sva));
  assign trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva[31]) | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_1_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_1_sva);
  assign trt_loop_else_mux_113_nl = MUX_s_1_2_2((trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      (chn_trt_in_rsci_d_mxwt[31]), chn_trt_in_rsci_d_mxwt[784]);
  assign trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva[0]) | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_2_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_2_sva);
  assign trt_loop_else_mux_114_nl = MUX_s_1_2_2((trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl),
      (chn_trt_in_rsci_d_mxwt[49]), chn_trt_in_rsci_d_mxwt[785]);
  assign trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva[31]) | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_2_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_2_sva);
  assign trt_loop_else_mux_115_nl = MUX_s_1_2_2((trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      (chn_trt_in_rsci_d_mxwt[80]), chn_trt_in_rsci_d_mxwt[785]);
  assign trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva[0]) | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_3_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_3_sva);
  assign trt_loop_else_mux_116_nl = MUX_s_1_2_2((trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl),
      (chn_trt_in_rsci_d_mxwt[98]), chn_trt_in_rsci_d_mxwt[786]);
  assign trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva[31]) | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_3_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_3_sva);
  assign trt_loop_else_mux_117_nl = MUX_s_1_2_2((trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      (chn_trt_in_rsci_d_mxwt[129]), chn_trt_in_rsci_d_mxwt[786]);
  assign trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva[0]) | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_4_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_4_sva);
  assign trt_loop_else_mux_118_nl = MUX_s_1_2_2((trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl),
      (chn_trt_in_rsci_d_mxwt[147]), chn_trt_in_rsci_d_mxwt[787]);
  assign trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva[31]) | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_4_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_4_sva);
  assign trt_loop_else_mux_119_nl = MUX_s_1_2_2((trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      (chn_trt_in_rsci_d_mxwt[178]), chn_trt_in_rsci_d_mxwt[787]);
  assign trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva[0]) | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_5_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_5_sva);
  assign trt_loop_else_mux_120_nl = MUX_s_1_2_2((trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl),
      (chn_trt_in_rsci_d_mxwt[196]), chn_trt_in_rsci_d_mxwt[788]);
  assign trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva[31]) | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_5_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_5_sva);
  assign trt_loop_else_mux_121_nl = MUX_s_1_2_2((trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      (chn_trt_in_rsci_d_mxwt[227]), chn_trt_in_rsci_d_mxwt[788]);
  assign trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva[0]) | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_6_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_6_sva);
  assign trt_loop_else_mux_122_nl = MUX_s_1_2_2((trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl),
      (chn_trt_in_rsci_d_mxwt[245]), chn_trt_in_rsci_d_mxwt[789]);
  assign trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva[31]) | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_6_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_6_sva);
  assign trt_loop_else_mux_123_nl = MUX_s_1_2_2((trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      (chn_trt_in_rsci_d_mxwt[276]), chn_trt_in_rsci_d_mxwt[789]);
  assign trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva[0]) | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_7_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_7_sva);
  assign trt_loop_else_mux_124_nl = MUX_s_1_2_2((trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl),
      (chn_trt_in_rsci_d_mxwt[294]), chn_trt_in_rsci_d_mxwt[790]);
  assign trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva[31]) | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_7_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_7_sva);
  assign trt_loop_else_mux_125_nl = MUX_s_1_2_2((trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      (chn_trt_in_rsci_d_mxwt[325]), chn_trt_in_rsci_d_mxwt[790]);
  assign trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva[0]) | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_8_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_8_sva);
  assign trt_loop_else_mux_126_nl = MUX_s_1_2_2((trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl),
      (chn_trt_in_rsci_d_mxwt[343]), chn_trt_in_rsci_d_mxwt[791]);
  assign trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva[31]) | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_8_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_8_sva);
  assign trt_loop_else_mux_127_nl = MUX_s_1_2_2((trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      (chn_trt_in_rsci_d_mxwt[374]), chn_trt_in_rsci_d_mxwt[791]);
  assign trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva[0]) | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_9_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_9_sva);
  assign trt_loop_else_mux_128_nl = MUX_s_1_2_2((trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl),
      (chn_trt_in_rsci_d_mxwt[392]), chn_trt_in_rsci_d_mxwt[792]);
  assign trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva[31]) | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_9_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_9_sva);
  assign trt_loop_else_mux_129_nl = MUX_s_1_2_2((trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      (chn_trt_in_rsci_d_mxwt[423]), chn_trt_in_rsci_d_mxwt[792]);
  assign trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva[0]) | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_10_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_10_sva);
  assign trt_loop_else_mux_130_nl = MUX_s_1_2_2((trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl),
      (chn_trt_in_rsci_d_mxwt[441]), chn_trt_in_rsci_d_mxwt[793]);
  assign trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva[31]) | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_10_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_10_sva);
  assign trt_loop_else_mux_131_nl = MUX_s_1_2_2((trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      (chn_trt_in_rsci_d_mxwt[472]), chn_trt_in_rsci_d_mxwt[793]);
  assign trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva[0]) | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_11_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_11_sva);
  assign trt_loop_else_mux_132_nl = MUX_s_1_2_2((trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl),
      (chn_trt_in_rsci_d_mxwt[490]), chn_trt_in_rsci_d_mxwt[794]);
  assign trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva[31]) | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_11_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_11_sva);
  assign trt_loop_else_mux_133_nl = MUX_s_1_2_2((trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      (chn_trt_in_rsci_d_mxwt[521]), chn_trt_in_rsci_d_mxwt[794]);
  assign trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva[0]) | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_12_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_12_sva);
  assign trt_loop_else_mux_134_nl = MUX_s_1_2_2((trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl),
      (chn_trt_in_rsci_d_mxwt[539]), chn_trt_in_rsci_d_mxwt[795]);
  assign trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva[31]) | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_12_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_12_sva);
  assign trt_loop_else_mux_135_nl = MUX_s_1_2_2((trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      (chn_trt_in_rsci_d_mxwt[570]), chn_trt_in_rsci_d_mxwt[795]);
  assign trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva[0]) | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_13_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_13_sva);
  assign trt_loop_else_mux_136_nl = MUX_s_1_2_2((trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl),
      (chn_trt_in_rsci_d_mxwt[588]), chn_trt_in_rsci_d_mxwt[796]);
  assign trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva[31]) | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_13_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_13_sva);
  assign trt_loop_else_mux_137_nl = MUX_s_1_2_2((trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      (chn_trt_in_rsci_d_mxwt[619]), chn_trt_in_rsci_d_mxwt[796]);
  assign trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva[0]) | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_14_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_14_sva);
  assign trt_loop_else_mux_138_nl = MUX_s_1_2_2((trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl),
      (chn_trt_in_rsci_d_mxwt[637]), chn_trt_in_rsci_d_mxwt[797]);
  assign trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva[31]) | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_14_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_14_sva);
  assign trt_loop_else_mux_139_nl = MUX_s_1_2_2((trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      (chn_trt_in_rsci_d_mxwt[668]), chn_trt_in_rsci_d_mxwt[797]);
  assign trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva[0]) | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_15_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_15_sva);
  assign trt_loop_else_mux_140_nl = MUX_s_1_2_2((trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl),
      (chn_trt_in_rsci_d_mxwt[686]), chn_trt_in_rsci_d_mxwt[798]);
  assign trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva[31]) | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_15_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_15_sva);
  assign trt_loop_else_mux_141_nl = MUX_s_1_2_2((trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      (chn_trt_in_rsci_d_mxwt[717]), chn_trt_in_rsci_d_mxwt[798]);
  assign trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva[0]) | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_sva);
  assign trt_loop_else_mux_142_nl = MUX_s_1_2_2((trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl),
      (chn_trt_in_rsci_d_mxwt[735]), chn_trt_in_rsci_d_mxwt[799]);
  assign trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl
      = ~((~((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva[31]) | IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_sva))
      | IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_sva);
  assign trt_loop_else_mux_143_nl = MUX_s_1_2_2((trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      (chn_trt_in_rsci_d_mxwt[766]), chn_trt_in_rsci_d_mxwt[799]);
  assign trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_2_sva));
  assign trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl
      = ~(MUX_v_30_2_2((trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_2_sva));
  assign trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_3_sva));
  assign trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl
      = ~(MUX_v_30_2_2((trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_3_sva));
  assign trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_4_sva));
  assign trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl
      = ~(MUX_v_30_2_2((trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_4_sva));
  assign trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_5_sva));
  assign trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl
      = ~(MUX_v_30_2_2((trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_5_sva));
  assign trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_6_sva));
  assign trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl
      = ~(MUX_v_30_2_2((trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_6_sva));
  assign trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_7_sva));
  assign trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl
      = ~(MUX_v_30_2_2((trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_7_sva));
  assign trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_8_sva));
  assign trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl
      = ~(MUX_v_30_2_2((trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_8_sva));
  assign trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_9_sva));
  assign trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl
      = ~(MUX_v_30_2_2((trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_9_sva));
  assign trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_10_sva));
  assign trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl
      = ~(MUX_v_30_2_2((trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_10_sva));
  assign trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_11_sva));
  assign trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl
      = ~(MUX_v_30_2_2((trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_11_sva));
  assign trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_12_sva));
  assign trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl
      = ~(MUX_v_30_2_2((trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_12_sva));
  assign trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_13_sva));
  assign trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl
      = ~(MUX_v_30_2_2((trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_13_sva));
  assign trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_14_sva));
  assign trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl
      = ~(MUX_v_30_2_2((trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_14_sva));
  assign trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_15_sva));
  assign trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl
      = ~(MUX_v_30_2_2((trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_15_sva));
  assign trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva[30:1]),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_sva));
  assign trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl
      = ~(MUX_v_30_2_2((trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl),
      30'b111111111111111111111111111111, IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_sva));
  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction
  function [29:0] MUX_v_30_2_2;
    input [29:0] input_0;
    input [29:0] input_1;
    input [0:0] sel;
    reg [29:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_30_2_2 = result;
  end
  endfunction
  function [49:0] conv_s2s_49_50 ;
    input [48:0] vector ;
  begin
    conv_s2s_49_50 = {vector[48], vector};
  end
  endfunction
  function [49:0] conv_u2s_1_50 ;
    input [0:0] vector ;
  begin
    conv_u2s_1_50 = {{49{1'b0}}, vector};
  end
  endfunction
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_relu_core
// ------------------------------------------------------------------
module SDP_X_X_relu_core (
  nvdla_core_clk, nvdla_core_rstn, chn_relu_in_rsc_z, chn_relu_in_rsc_vz, chn_relu_in_rsc_lz,
      cfg_relu_bypass_rsc_triosy_lz, cfg_precision, chn_relu_out_rsc_z, chn_relu_out_rsc_vz,
      chn_relu_out_rsc_lz, chn_relu_in_rsci_oswt, chn_relu_in_rsci_oswt_unreg, cfg_relu_bypass_rsci_d,
      chn_relu_out_rsci_oswt, cfg_relu_bypass_rsc_triosy_obj_oswt, chn_relu_out_rsci_oswt_unreg_pff
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [511:0] chn_relu_in_rsc_z;
  input chn_relu_in_rsc_vz;
  output chn_relu_in_rsc_lz;
  output cfg_relu_bypass_rsc_triosy_lz;
  input [1:0] cfg_precision;
  output [511:0] chn_relu_out_rsc_z;
  input chn_relu_out_rsc_vz;
  output chn_relu_out_rsc_lz;
  input chn_relu_in_rsci_oswt;
  output chn_relu_in_rsci_oswt_unreg;
  input cfg_relu_bypass_rsci_d;
  input chn_relu_out_rsci_oswt;
  input cfg_relu_bypass_rsc_triosy_obj_oswt;
  output chn_relu_out_rsci_oswt_unreg_pff;
// Interconnect Declarations
  wire core_wen;
  reg chn_relu_in_rsci_iswt0;
  wire chn_relu_in_rsci_bawt;
  wire chn_relu_in_rsci_wen_comp;
  reg chn_relu_in_rsci_ld_core_psct;
  wire [511:0] chn_relu_in_rsci_d_mxwt;
  wire core_wten;
  wire chn_relu_out_rsci_bawt;
  wire chn_relu_out_rsci_wen_comp;
  wire cfg_relu_bypass_rsc_triosy_obj_bawt;
  reg chn_relu_out_rsci_d_511;
  reg [7:0] chn_relu_out_rsci_d_510_503;
  reg [22:0] chn_relu_out_rsci_d_502_480;
  reg chn_relu_out_rsci_d_479;
  reg [7:0] chn_relu_out_rsci_d_478_471;
  reg [22:0] chn_relu_out_rsci_d_470_448;
  reg chn_relu_out_rsci_d_447;
  reg [7:0] chn_relu_out_rsci_d_446_439;
  reg [22:0] chn_relu_out_rsci_d_438_416;
  reg chn_relu_out_rsci_d_415;
  reg [7:0] chn_relu_out_rsci_d_414_407;
  reg [22:0] chn_relu_out_rsci_d_406_384;
  reg chn_relu_out_rsci_d_383;
  reg [7:0] chn_relu_out_rsci_d_382_375;
  reg [22:0] chn_relu_out_rsci_d_374_352;
  reg chn_relu_out_rsci_d_351;
  reg [7:0] chn_relu_out_rsci_d_350_343;
  reg [22:0] chn_relu_out_rsci_d_342_320;
  reg chn_relu_out_rsci_d_319;
  reg [7:0] chn_relu_out_rsci_d_318_311;
  reg [22:0] chn_relu_out_rsci_d_310_288;
  reg chn_relu_out_rsci_d_287;
  reg [7:0] chn_relu_out_rsci_d_286_279;
  reg [22:0] chn_relu_out_rsci_d_278_256;
  reg chn_relu_out_rsci_d_255;
  reg [7:0] chn_relu_out_rsci_d_254_247;
  reg [22:0] chn_relu_out_rsci_d_246_224;
  reg chn_relu_out_rsci_d_223;
  reg [7:0] chn_relu_out_rsci_d_222_215;
  reg [22:0] chn_relu_out_rsci_d_214_192;
  reg chn_relu_out_rsci_d_191;
  reg [7:0] chn_relu_out_rsci_d_190_183;
  reg [22:0] chn_relu_out_rsci_d_182_160;
  reg chn_relu_out_rsci_d_159;
  reg [7:0] chn_relu_out_rsci_d_158_151;
  reg [22:0] chn_relu_out_rsci_d_150_128;
  reg chn_relu_out_rsci_d_127;
  reg [7:0] chn_relu_out_rsci_d_126_119;
  reg [22:0] chn_relu_out_rsci_d_118_96;
  reg chn_relu_out_rsci_d_95;
  reg [7:0] chn_relu_out_rsci_d_94_87;
  reg [22:0] chn_relu_out_rsci_d_86_64;
  reg chn_relu_out_rsci_d_63;
  reg [7:0] chn_relu_out_rsci_d_62_55;
  reg [22:0] chn_relu_out_rsci_d_54_32;
  reg chn_relu_out_rsci_d_31;
  reg [7:0] chn_relu_out_rsci_d_30_23;
  reg [22:0] chn_relu_out_rsci_d_22_0;
  wire [1:0] fsm_output;
  wire and_dcpl_1;
  wire or_dcpl;
  wire and_dcpl_3;
  wire or_dcpl_1;
  wire or_dcpl_2;
  wire and_dcpl_7;
  wire and_dcpl_10;
  wire and_dcpl_15;
  wire or_dcpl_10;
  wire or_tmp_85;
  reg FpRelu_8U_23U_lor_1_lpi_1_dfm;
  reg FpRelu_8U_23U_lor_2_lpi_1_dfm;
  reg FpRelu_8U_23U_lor_3_lpi_1_dfm;
  reg FpRelu_8U_23U_lor_4_lpi_1_dfm;
  reg FpRelu_8U_23U_lor_5_lpi_1_dfm;
  reg FpRelu_8U_23U_lor_6_lpi_1_dfm;
  reg FpRelu_8U_23U_lor_7_lpi_1_dfm;
  reg FpRelu_8U_23U_lor_8_lpi_1_dfm;
  reg FpRelu_8U_23U_lor_9_lpi_1_dfm;
  reg FpRelu_8U_23U_lor_10_lpi_1_dfm;
  reg FpRelu_8U_23U_lor_11_lpi_1_dfm;
  reg FpRelu_8U_23U_lor_12_lpi_1_dfm;
  reg FpRelu_8U_23U_lor_13_lpi_1_dfm;
  reg FpRelu_8U_23U_lor_14_lpi_1_dfm;
  reg FpRelu_8U_23U_lor_15_lpi_1_dfm;
  reg FpRelu_8U_23U_lor_lpi_1_dfm;
  wire and_32_cse;
  wire and_34_cse;
  wire and_4_mdf;
  wire relu_loop_else_unequal_tmp;
  wire chn_relu_out_and_1_cse;
  wire chn_relu_out_and_5_cse;
  reg reg_cfg_relu_bypass_rsc_triosy_obj_ld_core_psct_cse;
  wire FpRelu_8U_23U_oelse_and_cse;
  reg reg_chn_relu_out_rsci_ld_core_psct_cse;
  wire or_dcpl_12;
  wire or_dcpl_13;
  wire or_dcpl_14;
  wire or_dcpl_15;
  wire or_dcpl_16;
  wire or_dcpl_17;
  wire or_dcpl_18;
  wire or_dcpl_19;
  wire or_dcpl_20;
  wire or_dcpl_21;
  wire or_dcpl_22;
  wire or_dcpl_23;
  wire or_dcpl_24;
  wire or_dcpl_25;
  wire or_dcpl_26;
  wire or_dcpl_27;
  wire relu_loop_asn_113;
  wire FpRelu_8U_23U_lor_1_lpi_1_dfm_mx0w0;
  wire FpRelu_8U_23U_lor_2_lpi_1_dfm_mx0w0;
  wire FpRelu_8U_23U_lor_3_lpi_1_dfm_mx0w0;
  wire FpRelu_8U_23U_lor_4_lpi_1_dfm_mx0w0;
  wire FpRelu_8U_23U_lor_5_lpi_1_dfm_mx0w0;
  wire FpRelu_8U_23U_lor_6_lpi_1_dfm_mx0w0;
  wire FpRelu_8U_23U_lor_7_lpi_1_dfm_mx0w0;
  wire FpRelu_8U_23U_lor_8_lpi_1_dfm_mx0w0;
  wire FpRelu_8U_23U_lor_9_lpi_1_dfm_mx0w0;
  wire FpRelu_8U_23U_lor_10_lpi_1_dfm_mx0w0;
  wire FpRelu_8U_23U_lor_11_lpi_1_dfm_mx0w0;
  wire FpRelu_8U_23U_lor_12_lpi_1_dfm_mx0w0;
  wire FpRelu_8U_23U_lor_13_lpi_1_dfm_mx0w0;
  wire FpRelu_8U_23U_lor_14_lpi_1_dfm_mx0w0;
  wire FpRelu_8U_23U_lor_15_lpi_1_dfm_mx0w0;
  wire FpRelu_8U_23U_lor_lpi_1_dfm_mx0w0;
  wire [30:0] relu_loop_else_else_qr_30_0_1_lpi_1_dfm;
  wire relu_loop_asn_115;
  wire [30:0] relu_loop_else_else_qr_30_0_2_lpi_1_dfm;
  wire [30:0] relu_loop_else_else_qr_30_0_3_lpi_1_dfm;
  wire [30:0] relu_loop_else_else_qr_30_0_4_lpi_1_dfm;
  wire [30:0] relu_loop_else_else_qr_30_0_5_lpi_1_dfm;
  wire [30:0] relu_loop_else_else_qr_30_0_6_lpi_1_dfm;
  wire [30:0] relu_loop_else_else_qr_30_0_7_lpi_1_dfm;
  wire [30:0] relu_loop_else_else_qr_30_0_8_lpi_1_dfm;
  wire [30:0] relu_loop_else_else_qr_30_0_9_lpi_1_dfm;
  wire [30:0] relu_loop_else_else_qr_30_0_10_lpi_1_dfm;
  wire [30:0] relu_loop_else_else_qr_30_0_11_lpi_1_dfm;
  wire [30:0] relu_loop_else_else_qr_30_0_12_lpi_1_dfm;
  wire [30:0] relu_loop_else_else_qr_30_0_13_lpi_1_dfm;
  wire [30:0] relu_loop_else_else_qr_30_0_14_lpi_1_dfm;
  wire [30:0] relu_loop_else_else_qr_30_0_15_lpi_1_dfm;
  wire [30:0] relu_loop_else_else_qr_30_0_lpi_1_dfm;
  wire nor_cse;
  wire nor_2_cse;
  wire nor_4_cse;
  wire nor_6_cse;
  wire nor_8_cse;
  wire nor_10_cse;
  wire nor_12_cse;
  wire nor_14_cse;
  wire nor_16_cse;
  wire nor_18_cse;
  wire nor_20_cse;
  wire nor_22_cse;
  wire nor_24_cse;
  wire nor_26_cse;
  wire nor_28_cse;
  wire nor_30_cse;
  wire chn_relu_in_rsci_ld_core_psct_mx0c0;
  wire chn_relu_out_rsci_d_31_mx0c1;
  wire[0:0] relu_loop_else_relu_loop_else_and_16_nl;
  wire[0:0] FpRelu_8U_23U_oelse_mux_32_nl;
  wire[0:0] relu_loop_else_relu_loop_else_and_17_nl;
  wire[0:0] FpRelu_8U_23U_oelse_mux_30_nl;
  wire[0:0] relu_loop_else_relu_loop_else_and_18_nl;
  wire[0:0] FpRelu_8U_23U_oelse_mux_28_nl;
  wire[0:0] relu_loop_else_relu_loop_else_and_19_nl;
  wire[0:0] FpRelu_8U_23U_oelse_mux_26_nl;
  wire[0:0] relu_loop_else_relu_loop_else_and_20_nl;
  wire[0:0] FpRelu_8U_23U_oelse_mux_24_nl;
  wire[0:0] relu_loop_else_relu_loop_else_and_21_nl;
  wire[0:0] FpRelu_8U_23U_oelse_mux_22_nl;
  wire[0:0] relu_loop_else_relu_loop_else_and_22_nl;
  wire[0:0] FpRelu_8U_23U_oelse_mux_20_nl;
  wire[0:0] relu_loop_else_relu_loop_else_and_23_nl;
  wire[0:0] FpRelu_8U_23U_oelse_mux_18_nl;
  wire[0:0] relu_loop_else_relu_loop_else_and_24_nl;
  wire[0:0] FpRelu_8U_23U_oelse_mux_16_nl;
  wire[0:0] relu_loop_else_relu_loop_else_and_25_nl;
  wire[0:0] FpRelu_8U_23U_oelse_mux_14_nl;
  wire[0:0] relu_loop_else_relu_loop_else_and_26_nl;
  wire[0:0] FpRelu_8U_23U_oelse_mux_12_nl;
  wire[0:0] relu_loop_else_relu_loop_else_and_27_nl;
  wire[0:0] FpRelu_8U_23U_oelse_mux_10_nl;
  wire[0:0] relu_loop_else_relu_loop_else_and_28_nl;
  wire[0:0] FpRelu_8U_23U_oelse_mux_8_nl;
  wire[0:0] relu_loop_else_relu_loop_else_and_29_nl;
  wire[0:0] FpRelu_8U_23U_oelse_mux_6_nl;
  wire[0:0] relu_loop_else_relu_loop_else_and_30_nl;
  wire[0:0] FpRelu_8U_23U_oelse_mux_4_nl;
  wire[0:0] relu_loop_else_relu_loop_else_and_31_nl;
  wire[0:0] FpRelu_8U_23U_oelse_mux_2_nl;
  wire[32:0] relu_loop_16_else_else_acc_nl;
  wire[33:0] nl_relu_loop_16_else_else_acc_nl;
  wire[32:0] relu_loop_15_else_else_acc_nl;
  wire[33:0] nl_relu_loop_15_else_else_acc_nl;
  wire[32:0] relu_loop_14_else_else_acc_nl;
  wire[33:0] nl_relu_loop_14_else_else_acc_nl;
  wire[32:0] relu_loop_13_else_else_acc_nl;
  wire[33:0] nl_relu_loop_13_else_else_acc_nl;
  wire[32:0] relu_loop_12_else_else_acc_nl;
  wire[33:0] nl_relu_loop_12_else_else_acc_nl;
  wire[32:0] relu_loop_11_else_else_acc_nl;
  wire[33:0] nl_relu_loop_11_else_else_acc_nl;
  wire[32:0] relu_loop_10_else_else_acc_nl;
  wire[33:0] nl_relu_loop_10_else_else_acc_nl;
  wire[32:0] relu_loop_9_else_else_acc_nl;
  wire[33:0] nl_relu_loop_9_else_else_acc_nl;
  wire[32:0] relu_loop_8_else_else_acc_nl;
  wire[33:0] nl_relu_loop_8_else_else_acc_nl;
  wire[32:0] relu_loop_7_else_else_acc_nl;
  wire[33:0] nl_relu_loop_7_else_else_acc_nl;
  wire[32:0] relu_loop_6_else_else_acc_nl;
  wire[33:0] nl_relu_loop_6_else_else_acc_nl;
  wire[32:0] relu_loop_5_else_else_acc_nl;
  wire[33:0] nl_relu_loop_5_else_else_acc_nl;
  wire[32:0] relu_loop_4_else_else_acc_nl;
  wire[33:0] nl_relu_loop_4_else_else_acc_nl;
  wire[32:0] relu_loop_3_else_else_acc_nl;
  wire[33:0] nl_relu_loop_3_else_else_acc_nl;
  wire[32:0] relu_loop_2_else_else_acc_nl;
  wire[33:0] nl_relu_loop_2_else_else_acc_nl;
  wire[32:0] relu_loop_1_else_else_acc_nl;
  wire[33:0] nl_relu_loop_1_else_else_acc_nl;
// Interconnect Declarations for Component Instantiations
  wire [511:0] nl_X_relu_core_chn_relu_out_rsci_inst_chn_relu_out_rsci_d;
  assign nl_X_relu_core_chn_relu_out_rsci_inst_chn_relu_out_rsci_d = {chn_relu_out_rsci_d_511
      , chn_relu_out_rsci_d_510_503 , chn_relu_out_rsci_d_502_480 , chn_relu_out_rsci_d_479
      , chn_relu_out_rsci_d_478_471 , chn_relu_out_rsci_d_470_448 , chn_relu_out_rsci_d_447
      , chn_relu_out_rsci_d_446_439 , chn_relu_out_rsci_d_438_416 , chn_relu_out_rsci_d_415
      , chn_relu_out_rsci_d_414_407 , chn_relu_out_rsci_d_406_384 , chn_relu_out_rsci_d_383
      , chn_relu_out_rsci_d_382_375 , chn_relu_out_rsci_d_374_352 , chn_relu_out_rsci_d_351
      , chn_relu_out_rsci_d_350_343 , chn_relu_out_rsci_d_342_320 , chn_relu_out_rsci_d_319
      , chn_relu_out_rsci_d_318_311 , chn_relu_out_rsci_d_310_288 , chn_relu_out_rsci_d_287
      , chn_relu_out_rsci_d_286_279 , chn_relu_out_rsci_d_278_256 , chn_relu_out_rsci_d_255
      , chn_relu_out_rsci_d_254_247 , chn_relu_out_rsci_d_246_224 , chn_relu_out_rsci_d_223
      , chn_relu_out_rsci_d_222_215 , chn_relu_out_rsci_d_214_192 , chn_relu_out_rsci_d_191
      , chn_relu_out_rsci_d_190_183 , chn_relu_out_rsci_d_182_160 , chn_relu_out_rsci_d_159
      , chn_relu_out_rsci_d_158_151 , chn_relu_out_rsci_d_150_128 , chn_relu_out_rsci_d_127
      , chn_relu_out_rsci_d_126_119 , chn_relu_out_rsci_d_118_96 , chn_relu_out_rsci_d_95
      , chn_relu_out_rsci_d_94_87 , chn_relu_out_rsci_d_86_64 , chn_relu_out_rsci_d_63
      , chn_relu_out_rsci_d_62_55 , chn_relu_out_rsci_d_54_32 , chn_relu_out_rsci_d_31
      , chn_relu_out_rsci_d_30_23 , chn_relu_out_rsci_d_22_0};
  SDP_X_X_relu_core_chn_relu_in_rsci X_relu_core_chn_relu_in_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_relu_in_rsc_z(chn_relu_in_rsc_z),
      .chn_relu_in_rsc_vz(chn_relu_in_rsc_vz),
      .chn_relu_in_rsc_lz(chn_relu_in_rsc_lz),
      .chn_relu_in_rsci_oswt(chn_relu_in_rsci_oswt),
      .core_wen(core_wen),
      .chn_relu_in_rsci_iswt0(chn_relu_in_rsci_iswt0),
      .chn_relu_in_rsci_bawt(chn_relu_in_rsci_bawt),
      .chn_relu_in_rsci_wen_comp(chn_relu_in_rsci_wen_comp),
      .chn_relu_in_rsci_ld_core_psct(chn_relu_in_rsci_ld_core_psct),
      .chn_relu_in_rsci_d_mxwt(chn_relu_in_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  SDP_X_X_relu_core_chn_relu_out_rsci X_relu_core_chn_relu_out_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_relu_out_rsc_z(chn_relu_out_rsc_z),
      .chn_relu_out_rsc_vz(chn_relu_out_rsc_vz),
      .chn_relu_out_rsc_lz(chn_relu_out_rsc_lz),
      .chn_relu_out_rsci_oswt(chn_relu_out_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_relu_out_rsci_iswt0(reg_cfg_relu_bypass_rsc_triosy_obj_ld_core_psct_cse),
      .chn_relu_out_rsci_bawt(chn_relu_out_rsci_bawt),
      .chn_relu_out_rsci_wen_comp(chn_relu_out_rsci_wen_comp),
      .chn_relu_out_rsci_ld_core_psct(reg_chn_relu_out_rsci_ld_core_psct_cse),
      .chn_relu_out_rsci_d(nl_X_relu_core_chn_relu_out_rsci_inst_chn_relu_out_rsci_d[511:0])
    );
  SDP_X_X_relu_core_cfg_relu_bypass_rsc_triosy_obj X_relu_core_cfg_relu_bypass_rsc_triosy_obj_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_relu_bypass_rsc_triosy_lz(cfg_relu_bypass_rsc_triosy_lz),
      .cfg_relu_bypass_rsc_triosy_obj_oswt(cfg_relu_bypass_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_relu_bypass_rsc_triosy_obj_iswt0(reg_cfg_relu_bypass_rsc_triosy_obj_ld_core_psct_cse),
      .cfg_relu_bypass_rsc_triosy_obj_bawt(cfg_relu_bypass_rsc_triosy_obj_bawt)
    );
  SDP_X_X_relu_core_staller X_relu_core_staller_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .chn_relu_in_rsci_wen_comp(chn_relu_in_rsci_wen_comp),
      .core_wten(core_wten),
      .chn_relu_out_rsci_wen_comp(chn_relu_out_rsci_wen_comp)
    );
  SDP_X_X_relu_core_core_fsm X_relu_core_core_fsm_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign nor_cse = ~(relu_loop_asn_115 | or_dcpl_12);
  assign chn_relu_out_and_1_cse = core_wen & (~(or_dcpl_2 | (fsm_output[0])));
  assign nor_2_cse = ~(relu_loop_asn_115 | or_dcpl_13);
  assign chn_relu_out_and_5_cse = core_wen & (and_32_cse | and_34_cse);
  assign nor_4_cse = ~(relu_loop_asn_115 | or_dcpl_14);
  assign nor_6_cse = ~(relu_loop_asn_115 | or_dcpl_15);
  assign nor_8_cse = ~(relu_loop_asn_115 | or_dcpl_16);
  assign nor_10_cse = ~(relu_loop_asn_115 | or_dcpl_17);
  assign nor_12_cse = ~(relu_loop_asn_115 | or_dcpl_18);
  assign nor_14_cse = ~(relu_loop_asn_115 | or_dcpl_19);
  assign nor_16_cse = ~(relu_loop_asn_115 | or_dcpl_20);
  assign nor_18_cse = ~(relu_loop_asn_115 | or_dcpl_21);
  assign nor_20_cse = ~(relu_loop_asn_115 | or_dcpl_22);
  assign nor_22_cse = ~(relu_loop_asn_115 | or_dcpl_23);
  assign nor_24_cse = ~(relu_loop_asn_115 | or_dcpl_24);
  assign nor_26_cse = ~(relu_loop_asn_115 | or_dcpl_25);
  assign nor_28_cse = ~(relu_loop_asn_115 | or_dcpl_26);
  assign nor_30_cse = ~(relu_loop_asn_115 | or_dcpl_27);
  assign FpRelu_8U_23U_oelse_and_cse = core_wen & (~(or_dcpl_2 | cfg_relu_bypass_rsci_d
      | (cfg_precision!=2'b10) | (fsm_output[0])));
  assign FpRelu_8U_23U_lor_lpi_1_dfm_mx0w0 = ~((chn_relu_in_rsci_d_mxwt[511]) & ((~((chn_relu_in_rsci_d_mxwt[502:480]!=23'b00000000000000000000000)))
      | (chn_relu_in_rsci_d_mxwt[510:503]!=8'b11111111)));
  assign FpRelu_8U_23U_lor_15_lpi_1_dfm_mx0w0 = ~((chn_relu_in_rsci_d_mxwt[479])
      & ((~((chn_relu_in_rsci_d_mxwt[470:448]!=23'b00000000000000000000000))) | (chn_relu_in_rsci_d_mxwt[478:471]!=8'b11111111)));
  assign FpRelu_8U_23U_lor_14_lpi_1_dfm_mx0w0 = ~((chn_relu_in_rsci_d_mxwt[447])
      & ((~((chn_relu_in_rsci_d_mxwt[438:416]!=23'b00000000000000000000000))) | (chn_relu_in_rsci_d_mxwt[446:439]!=8'b11111111)));
  assign FpRelu_8U_23U_lor_13_lpi_1_dfm_mx0w0 = ~((chn_relu_in_rsci_d_mxwt[415])
      & ((~((chn_relu_in_rsci_d_mxwt[406:384]!=23'b00000000000000000000000))) | (chn_relu_in_rsci_d_mxwt[414:407]!=8'b11111111)));
  assign FpRelu_8U_23U_lor_12_lpi_1_dfm_mx0w0 = ~((chn_relu_in_rsci_d_mxwt[383])
      & ((~((chn_relu_in_rsci_d_mxwt[374:352]!=23'b00000000000000000000000))) | (chn_relu_in_rsci_d_mxwt[382:375]!=8'b11111111)));
  assign FpRelu_8U_23U_lor_11_lpi_1_dfm_mx0w0 = ~((chn_relu_in_rsci_d_mxwt[351])
      & ((~((chn_relu_in_rsci_d_mxwt[342:320]!=23'b00000000000000000000000))) | (chn_relu_in_rsci_d_mxwt[350:343]!=8'b11111111)));
  assign FpRelu_8U_23U_lor_10_lpi_1_dfm_mx0w0 = ~((chn_relu_in_rsci_d_mxwt[319])
      & ((~((chn_relu_in_rsci_d_mxwt[310:288]!=23'b00000000000000000000000))) | (chn_relu_in_rsci_d_mxwt[318:311]!=8'b11111111)));
  assign FpRelu_8U_23U_lor_9_lpi_1_dfm_mx0w0 = ~((chn_relu_in_rsci_d_mxwt[287]) &
      ((~((chn_relu_in_rsci_d_mxwt[278:256]!=23'b00000000000000000000000))) | (chn_relu_in_rsci_d_mxwt[286:279]!=8'b11111111)));
  assign FpRelu_8U_23U_lor_8_lpi_1_dfm_mx0w0 = ~((chn_relu_in_rsci_d_mxwt[255]) &
      ((~((chn_relu_in_rsci_d_mxwt[246:224]!=23'b00000000000000000000000))) | (chn_relu_in_rsci_d_mxwt[254:247]!=8'b11111111)));
  assign FpRelu_8U_23U_lor_7_lpi_1_dfm_mx0w0 = ~((chn_relu_in_rsci_d_mxwt[223]) &
      ((~((chn_relu_in_rsci_d_mxwt[214:192]!=23'b00000000000000000000000))) | (chn_relu_in_rsci_d_mxwt[222:215]!=8'b11111111)));
  assign FpRelu_8U_23U_lor_6_lpi_1_dfm_mx0w0 = ~((chn_relu_in_rsci_d_mxwt[191]) &
      ((~((chn_relu_in_rsci_d_mxwt[182:160]!=23'b00000000000000000000000))) | (chn_relu_in_rsci_d_mxwt[190:183]!=8'b11111111)));
  assign FpRelu_8U_23U_lor_5_lpi_1_dfm_mx0w0 = ~((chn_relu_in_rsci_d_mxwt[159]) &
      ((~((chn_relu_in_rsci_d_mxwt[150:128]!=23'b00000000000000000000000))) | (chn_relu_in_rsci_d_mxwt[158:151]!=8'b11111111)));
  assign FpRelu_8U_23U_lor_4_lpi_1_dfm_mx0w0 = ~((chn_relu_in_rsci_d_mxwt[127]) &
      ((~((chn_relu_in_rsci_d_mxwt[118:96]!=23'b00000000000000000000000))) | (chn_relu_in_rsci_d_mxwt[126:119]!=8'b11111111)));
  assign FpRelu_8U_23U_lor_3_lpi_1_dfm_mx0w0 = ~((chn_relu_in_rsci_d_mxwt[95]) &
      ((~((chn_relu_in_rsci_d_mxwt[86:64]!=23'b00000000000000000000000))) | (chn_relu_in_rsci_d_mxwt[94:87]!=8'b11111111)));
  assign FpRelu_8U_23U_lor_2_lpi_1_dfm_mx0w0 = ~((chn_relu_in_rsci_d_mxwt[63]) &
      ((~((chn_relu_in_rsci_d_mxwt[54:32]!=23'b00000000000000000000000))) | (chn_relu_in_rsci_d_mxwt[62:55]!=8'b11111111)));
  assign FpRelu_8U_23U_lor_1_lpi_1_dfm_mx0w0 = ~((chn_relu_in_rsci_d_mxwt[31]) &
      ((~((chn_relu_in_rsci_d_mxwt[22:0]!=23'b00000000000000000000000))) | (chn_relu_in_rsci_d_mxwt[30:23]!=8'b11111111)));
  assign nl_relu_loop_16_else_else_acc_nl = conv_s2u_32_33(~ (chn_relu_in_rsci_d_mxwt[511:480]))
      + 33'b1;
  assign relu_loop_16_else_else_acc_nl = nl_relu_loop_16_else_else_acc_nl[32:0];
  assign relu_loop_else_else_qr_30_0_lpi_1_dfm = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      (chn_relu_in_rsci_d_mxwt[510:480]), (readslicef_33_1_32((relu_loop_16_else_else_acc_nl))));
  assign nl_relu_loop_15_else_else_acc_nl = conv_s2u_32_33(~ (chn_relu_in_rsci_d_mxwt[479:448]))
      + 33'b1;
  assign relu_loop_15_else_else_acc_nl = nl_relu_loop_15_else_else_acc_nl[32:0];
  assign relu_loop_else_else_qr_30_0_15_lpi_1_dfm = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      (chn_relu_in_rsci_d_mxwt[478:448]), (readslicef_33_1_32((relu_loop_15_else_else_acc_nl))));
  assign nl_relu_loop_14_else_else_acc_nl = conv_s2u_32_33(~ (chn_relu_in_rsci_d_mxwt[447:416]))
      + 33'b1;
  assign relu_loop_14_else_else_acc_nl = nl_relu_loop_14_else_else_acc_nl[32:0];
  assign relu_loop_else_else_qr_30_0_14_lpi_1_dfm = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      (chn_relu_in_rsci_d_mxwt[446:416]), (readslicef_33_1_32((relu_loop_14_else_else_acc_nl))));
  assign nl_relu_loop_13_else_else_acc_nl = conv_s2u_32_33(~ (chn_relu_in_rsci_d_mxwt[415:384]))
      + 33'b1;
  assign relu_loop_13_else_else_acc_nl = nl_relu_loop_13_else_else_acc_nl[32:0];
  assign relu_loop_else_else_qr_30_0_13_lpi_1_dfm = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      (chn_relu_in_rsci_d_mxwt[414:384]), (readslicef_33_1_32((relu_loop_13_else_else_acc_nl))));
  assign nl_relu_loop_12_else_else_acc_nl = conv_s2u_32_33(~ (chn_relu_in_rsci_d_mxwt[383:352]))
      + 33'b1;
  assign relu_loop_12_else_else_acc_nl = nl_relu_loop_12_else_else_acc_nl[32:0];
  assign relu_loop_else_else_qr_30_0_12_lpi_1_dfm = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      (chn_relu_in_rsci_d_mxwt[382:352]), (readslicef_33_1_32((relu_loop_12_else_else_acc_nl))));
  assign nl_relu_loop_11_else_else_acc_nl = conv_s2u_32_33(~ (chn_relu_in_rsci_d_mxwt[351:320]))
      + 33'b1;
  assign relu_loop_11_else_else_acc_nl = nl_relu_loop_11_else_else_acc_nl[32:0];
  assign relu_loop_else_else_qr_30_0_11_lpi_1_dfm = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      (chn_relu_in_rsci_d_mxwt[350:320]), (readslicef_33_1_32((relu_loop_11_else_else_acc_nl))));
  assign nl_relu_loop_10_else_else_acc_nl = conv_s2u_32_33(~ (chn_relu_in_rsci_d_mxwt[319:288]))
      + 33'b1;
  assign relu_loop_10_else_else_acc_nl = nl_relu_loop_10_else_else_acc_nl[32:0];
  assign relu_loop_else_else_qr_30_0_10_lpi_1_dfm = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      (chn_relu_in_rsci_d_mxwt[318:288]), (readslicef_33_1_32((relu_loop_10_else_else_acc_nl))));
  assign nl_relu_loop_9_else_else_acc_nl = conv_s2u_32_33(~ (chn_relu_in_rsci_d_mxwt[287:256]))
      + 33'b1;
  assign relu_loop_9_else_else_acc_nl = nl_relu_loop_9_else_else_acc_nl[32:0];
  assign relu_loop_else_else_qr_30_0_9_lpi_1_dfm = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      (chn_relu_in_rsci_d_mxwt[286:256]), (readslicef_33_1_32((relu_loop_9_else_else_acc_nl))));
  assign nl_relu_loop_8_else_else_acc_nl = conv_s2u_32_33(~ (chn_relu_in_rsci_d_mxwt[255:224]))
      + 33'b1;
  assign relu_loop_8_else_else_acc_nl = nl_relu_loop_8_else_else_acc_nl[32:0];
  assign relu_loop_else_else_qr_30_0_8_lpi_1_dfm = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      (chn_relu_in_rsci_d_mxwt[254:224]), (readslicef_33_1_32((relu_loop_8_else_else_acc_nl))));
  assign nl_relu_loop_7_else_else_acc_nl = conv_s2u_32_33(~ (chn_relu_in_rsci_d_mxwt[223:192]))
      + 33'b1;
  assign relu_loop_7_else_else_acc_nl = nl_relu_loop_7_else_else_acc_nl[32:0];
  assign relu_loop_else_else_qr_30_0_7_lpi_1_dfm = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      (chn_relu_in_rsci_d_mxwt[222:192]), (readslicef_33_1_32((relu_loop_7_else_else_acc_nl))));
  assign nl_relu_loop_6_else_else_acc_nl = conv_s2u_32_33(~ (chn_relu_in_rsci_d_mxwt[191:160]))
      + 33'b1;
  assign relu_loop_6_else_else_acc_nl = nl_relu_loop_6_else_else_acc_nl[32:0];
  assign relu_loop_else_else_qr_30_0_6_lpi_1_dfm = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      (chn_relu_in_rsci_d_mxwt[190:160]), (readslicef_33_1_32((relu_loop_6_else_else_acc_nl))));
  assign nl_relu_loop_5_else_else_acc_nl = conv_s2u_32_33(~ (chn_relu_in_rsci_d_mxwt[159:128]))
      + 33'b1;
  assign relu_loop_5_else_else_acc_nl = nl_relu_loop_5_else_else_acc_nl[32:0];
  assign relu_loop_else_else_qr_30_0_5_lpi_1_dfm = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      (chn_relu_in_rsci_d_mxwt[158:128]), (readslicef_33_1_32((relu_loop_5_else_else_acc_nl))));
  assign nl_relu_loop_4_else_else_acc_nl = conv_s2u_32_33(~ (chn_relu_in_rsci_d_mxwt[127:96]))
      + 33'b1;
  assign relu_loop_4_else_else_acc_nl = nl_relu_loop_4_else_else_acc_nl[32:0];
  assign relu_loop_else_else_qr_30_0_4_lpi_1_dfm = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      (chn_relu_in_rsci_d_mxwt[126:96]), (readslicef_33_1_32((relu_loop_4_else_else_acc_nl))));
  assign nl_relu_loop_3_else_else_acc_nl = conv_s2u_32_33(~ (chn_relu_in_rsci_d_mxwt[95:64]))
      + 33'b1;
  assign relu_loop_3_else_else_acc_nl = nl_relu_loop_3_else_else_acc_nl[32:0];
  assign relu_loop_else_else_qr_30_0_3_lpi_1_dfm = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      (chn_relu_in_rsci_d_mxwt[94:64]), (readslicef_33_1_32((relu_loop_3_else_else_acc_nl))));
  assign nl_relu_loop_2_else_else_acc_nl = conv_s2u_32_33(~ (chn_relu_in_rsci_d_mxwt[63:32]))
      + 33'b1;
  assign relu_loop_2_else_else_acc_nl = nl_relu_loop_2_else_else_acc_nl[32:0];
  assign relu_loop_else_else_qr_30_0_2_lpi_1_dfm = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      (chn_relu_in_rsci_d_mxwt[62:32]), (readslicef_33_1_32((relu_loop_2_else_else_acc_nl))));
  assign nl_relu_loop_1_else_else_acc_nl = conv_s2u_32_33(~ (chn_relu_in_rsci_d_mxwt[31:0]))
      + 33'b1;
  assign relu_loop_1_else_else_acc_nl = nl_relu_loop_1_else_else_acc_nl[32:0];
  assign relu_loop_else_else_qr_30_0_1_lpi_1_dfm = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      (chn_relu_in_rsci_d_mxwt[30:0]), (readslicef_33_1_32((relu_loop_1_else_else_acc_nl))));
  assign relu_loop_else_unequal_tmp = ~((cfg_precision==2'b10));
  assign and_4_mdf = chn_relu_in_rsci_bawt & (chn_relu_out_rsci_bawt | (~ reg_chn_relu_out_rsci_ld_core_psct_cse))
      & (cfg_relu_bypass_rsc_triosy_obj_bawt | (~ reg_chn_relu_out_rsci_ld_core_psct_cse));
  assign relu_loop_asn_113 = ~(relu_loop_else_unequal_tmp | cfg_relu_bypass_rsci_d);
  assign relu_loop_asn_115 = relu_loop_else_unequal_tmp & (~ cfg_relu_bypass_rsci_d);
  assign and_dcpl_1 = chn_relu_out_rsci_bawt & cfg_relu_bypass_rsc_triosy_obj_bawt;
  assign or_dcpl = and_dcpl_1 | (~ reg_chn_relu_out_rsci_ld_core_psct_cse);
  assign and_dcpl_3 = and_dcpl_1 & reg_chn_relu_out_rsci_ld_core_psct_cse;
  assign or_dcpl_1 = ~(chn_relu_out_rsci_bawt & cfg_relu_bypass_rsc_triosy_obj_bawt);
  assign or_dcpl_2 = ~((~(or_dcpl_1 & reg_chn_relu_out_rsci_ld_core_psct_cse)) &
      chn_relu_in_rsci_bawt);
  assign and_dcpl_7 = chn_relu_in_rsci_bawt & cfg_relu_bypass_rsci_d;
  assign and_dcpl_10 = chn_relu_in_rsci_bawt & (~ cfg_relu_bypass_rsci_d);
  assign and_dcpl_15 = and_dcpl_1 & reg_chn_relu_out_rsci_ld_core_psct_cse & (~ chn_relu_in_rsci_bawt);
  assign or_dcpl_10 = (cfg_precision!=2'b10);
  assign and_32_cse = or_dcpl & and_dcpl_7 & (fsm_output[1]);
  assign and_34_cse = or_dcpl & and_dcpl_10 & (fsm_output[1]);
  assign or_tmp_85 = or_dcpl & chn_relu_in_rsci_bawt & (fsm_output[1]);
  assign chn_relu_in_rsci_ld_core_psct_mx0c0 = and_4_mdf | (fsm_output[0]);
  assign chn_relu_out_rsci_d_31_mx0c1 = and_34_cse | (and_dcpl_3 & and_dcpl_10);
  assign chn_relu_in_rsci_oswt_unreg = or_tmp_85;
  assign chn_relu_out_rsci_oswt_unreg_pff = and_dcpl_3;
  assign or_dcpl_12 = (relu_loop_asn_113 & FpRelu_8U_23U_lor_1_lpi_1_dfm_mx0w0) |
      cfg_relu_bypass_rsci_d;
  assign or_dcpl_13 = (relu_loop_asn_113 & FpRelu_8U_23U_lor_2_lpi_1_dfm_mx0w0) |
      cfg_relu_bypass_rsci_d;
  assign or_dcpl_14 = (relu_loop_asn_113 & FpRelu_8U_23U_lor_3_lpi_1_dfm_mx0w0) |
      cfg_relu_bypass_rsci_d;
  assign or_dcpl_15 = (relu_loop_asn_113 & FpRelu_8U_23U_lor_4_lpi_1_dfm_mx0w0) |
      cfg_relu_bypass_rsci_d;
  assign or_dcpl_16 = (relu_loop_asn_113 & FpRelu_8U_23U_lor_5_lpi_1_dfm_mx0w0) |
      cfg_relu_bypass_rsci_d;
  assign or_dcpl_17 = (relu_loop_asn_113 & FpRelu_8U_23U_lor_6_lpi_1_dfm_mx0w0) |
      cfg_relu_bypass_rsci_d;
  assign or_dcpl_18 = (relu_loop_asn_113 & FpRelu_8U_23U_lor_7_lpi_1_dfm_mx0w0) |
      cfg_relu_bypass_rsci_d;
  assign or_dcpl_19 = (relu_loop_asn_113 & FpRelu_8U_23U_lor_8_lpi_1_dfm_mx0w0) |
      cfg_relu_bypass_rsci_d;
  assign or_dcpl_20 = (relu_loop_asn_113 & FpRelu_8U_23U_lor_9_lpi_1_dfm_mx0w0) |
      cfg_relu_bypass_rsci_d;
  assign or_dcpl_21 = (relu_loop_asn_113 & FpRelu_8U_23U_lor_10_lpi_1_dfm_mx0w0)
      | cfg_relu_bypass_rsci_d;
  assign or_dcpl_22 = (relu_loop_asn_113 & FpRelu_8U_23U_lor_11_lpi_1_dfm_mx0w0)
      | cfg_relu_bypass_rsci_d;
  assign or_dcpl_23 = (relu_loop_asn_113 & FpRelu_8U_23U_lor_12_lpi_1_dfm_mx0w0)
      | cfg_relu_bypass_rsci_d;
  assign or_dcpl_24 = (relu_loop_asn_113 & FpRelu_8U_23U_lor_13_lpi_1_dfm_mx0w0)
      | cfg_relu_bypass_rsci_d;
  assign or_dcpl_25 = (relu_loop_asn_113 & FpRelu_8U_23U_lor_14_lpi_1_dfm_mx0w0)
      | cfg_relu_bypass_rsci_d;
  assign or_dcpl_26 = (relu_loop_asn_113 & FpRelu_8U_23U_lor_15_lpi_1_dfm_mx0w0)
      | cfg_relu_bypass_rsci_d;
  assign or_dcpl_27 = (relu_loop_asn_113 & FpRelu_8U_23U_lor_lpi_1_dfm_mx0w0) | cfg_relu_bypass_rsci_d;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_relu_in_rsci_iswt0 <= 1'b0;
      reg_cfg_relu_bypass_rsc_triosy_obj_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen ) begin
      chn_relu_in_rsci_iswt0 <= ~((~ and_4_mdf) & (fsm_output[1]));
      reg_cfg_relu_bypass_rsc_triosy_obj_ld_core_psct_cse <= or_tmp_85;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_relu_in_rsci_ld_core_psct <= 1'b0;
    end
    else if ( core_wen & chn_relu_in_rsci_ld_core_psct_mx0c0 ) begin
      chn_relu_in_rsci_ld_core_psct <= chn_relu_in_rsci_ld_core_psct_mx0c0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_relu_out_rsci_d_22_0 <= 23'b0;
    end
    else if ( core_wen & (~(or_dcpl_2 | ((or_dcpl_1 | (~ reg_chn_relu_out_rsci_ld_core_psct_cse)
        | (~ chn_relu_in_rsci_bawt)) & (fsm_output[0])))) ) begin
      chn_relu_out_rsci_d_22_0 <= MUX1HOT_v_23_3_2(({{22{FpRelu_8U_23U_lor_1_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_1_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_1_lpi_1_dfm[22:0]),
          (chn_relu_in_rsci_d_mxwt[22:0]), {nor_cse , relu_loop_asn_115 , or_dcpl_12});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_relu_out_rsci_d_30_23 <= 8'b0;
      chn_relu_out_rsci_d_54_32 <= 23'b0;
      chn_relu_out_rsci_d_62_55 <= 8'b0;
      chn_relu_out_rsci_d_86_64 <= 23'b0;
      chn_relu_out_rsci_d_94_87 <= 8'b0;
      chn_relu_out_rsci_d_118_96 <= 23'b0;
      chn_relu_out_rsci_d_126_119 <= 8'b0;
      chn_relu_out_rsci_d_150_128 <= 23'b0;
      chn_relu_out_rsci_d_158_151 <= 8'b0;
      chn_relu_out_rsci_d_182_160 <= 23'b0;
      chn_relu_out_rsci_d_190_183 <= 8'b0;
      chn_relu_out_rsci_d_214_192 <= 23'b0;
      chn_relu_out_rsci_d_222_215 <= 8'b0;
      chn_relu_out_rsci_d_246_224 <= 23'b0;
      chn_relu_out_rsci_d_254_247 <= 8'b0;
      chn_relu_out_rsci_d_278_256 <= 23'b0;
      chn_relu_out_rsci_d_286_279 <= 8'b0;
      chn_relu_out_rsci_d_310_288 <= 23'b0;
      chn_relu_out_rsci_d_318_311 <= 8'b0;
      chn_relu_out_rsci_d_342_320 <= 23'b0;
      chn_relu_out_rsci_d_350_343 <= 8'b0;
      chn_relu_out_rsci_d_374_352 <= 23'b0;
      chn_relu_out_rsci_d_382_375 <= 8'b0;
      chn_relu_out_rsci_d_406_384 <= 23'b0;
      chn_relu_out_rsci_d_414_407 <= 8'b0;
      chn_relu_out_rsci_d_438_416 <= 23'b0;
      chn_relu_out_rsci_d_446_439 <= 8'b0;
      chn_relu_out_rsci_d_470_448 <= 23'b0;
      chn_relu_out_rsci_d_478_471 <= 8'b0;
      chn_relu_out_rsci_d_502_480 <= 23'b0;
      chn_relu_out_rsci_d_510_503 <= 8'b0;
    end
    else if ( chn_relu_out_and_1_cse ) begin
      chn_relu_out_rsci_d_30_23 <= MUX1HOT_v_8_3_2(({{7{FpRelu_8U_23U_lor_1_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_1_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_1_lpi_1_dfm[30:23]),
          (chn_relu_in_rsci_d_mxwt[30:23]), {nor_cse , relu_loop_asn_115 , or_dcpl_12});
      chn_relu_out_rsci_d_54_32 <= MUX1HOT_v_23_3_2(({{22{FpRelu_8U_23U_lor_2_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_2_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_2_lpi_1_dfm[22:0]),
          (chn_relu_in_rsci_d_mxwt[54:32]), {nor_2_cse , relu_loop_asn_115 , or_dcpl_13});
      chn_relu_out_rsci_d_62_55 <= MUX1HOT_v_8_3_2(({{7{FpRelu_8U_23U_lor_2_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_2_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_2_lpi_1_dfm[30:23]),
          (chn_relu_in_rsci_d_mxwt[62:55]), {nor_2_cse , relu_loop_asn_115 , or_dcpl_13});
      chn_relu_out_rsci_d_86_64 <= MUX1HOT_v_23_3_2(({{22{FpRelu_8U_23U_lor_3_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_3_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_3_lpi_1_dfm[22:0]),
          (chn_relu_in_rsci_d_mxwt[86:64]), {nor_4_cse , relu_loop_asn_115 , or_dcpl_14});
      chn_relu_out_rsci_d_94_87 <= MUX1HOT_v_8_3_2(({{7{FpRelu_8U_23U_lor_3_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_3_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_3_lpi_1_dfm[30:23]),
          (chn_relu_in_rsci_d_mxwt[94:87]), {nor_4_cse , relu_loop_asn_115 , or_dcpl_14});
      chn_relu_out_rsci_d_118_96 <= MUX1HOT_v_23_3_2(({{22{FpRelu_8U_23U_lor_4_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_4_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_4_lpi_1_dfm[22:0]),
          (chn_relu_in_rsci_d_mxwt[118:96]), {nor_6_cse , relu_loop_asn_115 , or_dcpl_15});
      chn_relu_out_rsci_d_126_119 <= MUX1HOT_v_8_3_2(({{7{FpRelu_8U_23U_lor_4_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_4_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_4_lpi_1_dfm[30:23]),
          (chn_relu_in_rsci_d_mxwt[126:119]), {nor_6_cse , relu_loop_asn_115 , or_dcpl_15});
      chn_relu_out_rsci_d_150_128 <= MUX1HOT_v_23_3_2(({{22{FpRelu_8U_23U_lor_5_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_5_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_5_lpi_1_dfm[22:0]),
          (chn_relu_in_rsci_d_mxwt[150:128]), {nor_8_cse , relu_loop_asn_115 , or_dcpl_16});
      chn_relu_out_rsci_d_158_151 <= MUX1HOT_v_8_3_2(({{7{FpRelu_8U_23U_lor_5_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_5_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_5_lpi_1_dfm[30:23]),
          (chn_relu_in_rsci_d_mxwt[158:151]), {nor_8_cse , relu_loop_asn_115 , or_dcpl_16});
      chn_relu_out_rsci_d_182_160 <= MUX1HOT_v_23_3_2(({{22{FpRelu_8U_23U_lor_6_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_6_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_6_lpi_1_dfm[22:0]),
          (chn_relu_in_rsci_d_mxwt[182:160]), {nor_10_cse , relu_loop_asn_115 , or_dcpl_17});
      chn_relu_out_rsci_d_190_183 <= MUX1HOT_v_8_3_2(({{7{FpRelu_8U_23U_lor_6_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_6_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_6_lpi_1_dfm[30:23]),
          (chn_relu_in_rsci_d_mxwt[190:183]), {nor_10_cse , relu_loop_asn_115 , or_dcpl_17});
      chn_relu_out_rsci_d_214_192 <= MUX1HOT_v_23_3_2(({{22{FpRelu_8U_23U_lor_7_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_7_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_7_lpi_1_dfm[22:0]),
          (chn_relu_in_rsci_d_mxwt[214:192]), {nor_12_cse , relu_loop_asn_115 , or_dcpl_18});
      chn_relu_out_rsci_d_222_215 <= MUX1HOT_v_8_3_2(({{7{FpRelu_8U_23U_lor_7_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_7_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_7_lpi_1_dfm[30:23]),
          (chn_relu_in_rsci_d_mxwt[222:215]), {nor_12_cse , relu_loop_asn_115 , or_dcpl_18});
      chn_relu_out_rsci_d_246_224 <= MUX1HOT_v_23_3_2(({{22{FpRelu_8U_23U_lor_8_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_8_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_8_lpi_1_dfm[22:0]),
          (chn_relu_in_rsci_d_mxwt[246:224]), {nor_14_cse , relu_loop_asn_115 , or_dcpl_19});
      chn_relu_out_rsci_d_254_247 <= MUX1HOT_v_8_3_2(({{7{FpRelu_8U_23U_lor_8_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_8_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_8_lpi_1_dfm[30:23]),
          (chn_relu_in_rsci_d_mxwt[254:247]), {nor_14_cse , relu_loop_asn_115 , or_dcpl_19});
      chn_relu_out_rsci_d_278_256 <= MUX1HOT_v_23_3_2(({{22{FpRelu_8U_23U_lor_9_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_9_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_9_lpi_1_dfm[22:0]),
          (chn_relu_in_rsci_d_mxwt[278:256]), {nor_16_cse , relu_loop_asn_115 , or_dcpl_20});
      chn_relu_out_rsci_d_286_279 <= MUX1HOT_v_8_3_2(({{7{FpRelu_8U_23U_lor_9_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_9_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_9_lpi_1_dfm[30:23]),
          (chn_relu_in_rsci_d_mxwt[286:279]), {nor_16_cse , relu_loop_asn_115 , or_dcpl_20});
      chn_relu_out_rsci_d_310_288 <= MUX1HOT_v_23_3_2(({{22{FpRelu_8U_23U_lor_10_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_10_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_10_lpi_1_dfm[22:0]),
          (chn_relu_in_rsci_d_mxwt[310:288]), {nor_18_cse , relu_loop_asn_115 , or_dcpl_21});
      chn_relu_out_rsci_d_318_311 <= MUX1HOT_v_8_3_2(({{7{FpRelu_8U_23U_lor_10_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_10_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_10_lpi_1_dfm[30:23]),
          (chn_relu_in_rsci_d_mxwt[318:311]), {nor_18_cse , relu_loop_asn_115 , or_dcpl_21});
      chn_relu_out_rsci_d_342_320 <= MUX1HOT_v_23_3_2(({{22{FpRelu_8U_23U_lor_11_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_11_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_11_lpi_1_dfm[22:0]),
          (chn_relu_in_rsci_d_mxwt[342:320]), {nor_20_cse , relu_loop_asn_115 , or_dcpl_22});
      chn_relu_out_rsci_d_350_343 <= MUX1HOT_v_8_3_2(({{7{FpRelu_8U_23U_lor_11_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_11_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_11_lpi_1_dfm[30:23]),
          (chn_relu_in_rsci_d_mxwt[350:343]), {nor_20_cse , relu_loop_asn_115 , or_dcpl_22});
      chn_relu_out_rsci_d_374_352 <= MUX1HOT_v_23_3_2(({{22{FpRelu_8U_23U_lor_12_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_12_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_12_lpi_1_dfm[22:0]),
          (chn_relu_in_rsci_d_mxwt[374:352]), {nor_22_cse , relu_loop_asn_115 , or_dcpl_23});
      chn_relu_out_rsci_d_382_375 <= MUX1HOT_v_8_3_2(({{7{FpRelu_8U_23U_lor_12_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_12_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_12_lpi_1_dfm[30:23]),
          (chn_relu_in_rsci_d_mxwt[382:375]), {nor_22_cse , relu_loop_asn_115 , or_dcpl_23});
      chn_relu_out_rsci_d_406_384 <= MUX1HOT_v_23_3_2(({{22{FpRelu_8U_23U_lor_13_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_13_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_13_lpi_1_dfm[22:0]),
          (chn_relu_in_rsci_d_mxwt[406:384]), {nor_24_cse , relu_loop_asn_115 , or_dcpl_24});
      chn_relu_out_rsci_d_414_407 <= MUX1HOT_v_8_3_2(({{7{FpRelu_8U_23U_lor_13_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_13_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_13_lpi_1_dfm[30:23]),
          (chn_relu_in_rsci_d_mxwt[414:407]), {nor_24_cse , relu_loop_asn_115 , or_dcpl_24});
      chn_relu_out_rsci_d_438_416 <= MUX1HOT_v_23_3_2(({{22{FpRelu_8U_23U_lor_14_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_14_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_14_lpi_1_dfm[22:0]),
          (chn_relu_in_rsci_d_mxwt[438:416]), {nor_26_cse , relu_loop_asn_115 , or_dcpl_25});
      chn_relu_out_rsci_d_446_439 <= MUX1HOT_v_8_3_2(({{7{FpRelu_8U_23U_lor_14_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_14_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_14_lpi_1_dfm[30:23]),
          (chn_relu_in_rsci_d_mxwt[446:439]), {nor_26_cse , relu_loop_asn_115 , or_dcpl_25});
      chn_relu_out_rsci_d_470_448 <= MUX1HOT_v_23_3_2(({{22{FpRelu_8U_23U_lor_15_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_15_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_15_lpi_1_dfm[22:0]),
          (chn_relu_in_rsci_d_mxwt[470:448]), {nor_28_cse , relu_loop_asn_115 , or_dcpl_26});
      chn_relu_out_rsci_d_478_471 <= MUX1HOT_v_8_3_2(({{7{FpRelu_8U_23U_lor_15_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_15_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_15_lpi_1_dfm[30:23]),
          (chn_relu_in_rsci_d_mxwt[478:471]), {nor_28_cse , relu_loop_asn_115 , or_dcpl_26});
      chn_relu_out_rsci_d_502_480 <= MUX1HOT_v_23_3_2(({{22{FpRelu_8U_23U_lor_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_lpi_1_dfm[22:0]),
          (chn_relu_in_rsci_d_mxwt[502:480]), {nor_30_cse , relu_loop_asn_115 , or_dcpl_27});
      chn_relu_out_rsci_d_510_503 <= MUX1HOT_v_8_3_2(({{7{FpRelu_8U_23U_lor_lpi_1_dfm_mx0w0}},
          FpRelu_8U_23U_lor_lpi_1_dfm_mx0w0}), (relu_loop_else_else_qr_30_0_lpi_1_dfm[30:23]),
          (chn_relu_in_rsci_d_mxwt[510:503]), {nor_30_cse , relu_loop_asn_115 , or_dcpl_27});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_relu_out_rsci_d_31 <= 1'b0;
    end
    else if ( core_wen & (and_32_cse | (and_dcpl_3 & and_dcpl_7) | chn_relu_out_rsci_d_31_mx0c1)
        ) begin
      chn_relu_out_rsci_d_31 <= MUX_s_1_2_2((chn_relu_in_rsci_d_mxwt[31]), (relu_loop_else_relu_loop_else_and_16_nl),
          chn_relu_out_rsci_d_31_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_relu_out_rsci_d_63 <= 1'b0;
      chn_relu_out_rsci_d_95 <= 1'b0;
      chn_relu_out_rsci_d_127 <= 1'b0;
      chn_relu_out_rsci_d_159 <= 1'b0;
      chn_relu_out_rsci_d_191 <= 1'b0;
      chn_relu_out_rsci_d_223 <= 1'b0;
      chn_relu_out_rsci_d_255 <= 1'b0;
      chn_relu_out_rsci_d_287 <= 1'b0;
      chn_relu_out_rsci_d_319 <= 1'b0;
      chn_relu_out_rsci_d_351 <= 1'b0;
      chn_relu_out_rsci_d_383 <= 1'b0;
      chn_relu_out_rsci_d_415 <= 1'b0;
      chn_relu_out_rsci_d_447 <= 1'b0;
      chn_relu_out_rsci_d_479 <= 1'b0;
      chn_relu_out_rsci_d_511 <= 1'b0;
    end
    else if ( chn_relu_out_and_5_cse ) begin
      chn_relu_out_rsci_d_63 <= MUX_s_1_2_2((chn_relu_in_rsci_d_mxwt[63]), (relu_loop_else_relu_loop_else_and_17_nl),
          and_34_cse);
      chn_relu_out_rsci_d_95 <= MUX_s_1_2_2((chn_relu_in_rsci_d_mxwt[95]), (relu_loop_else_relu_loop_else_and_18_nl),
          and_34_cse);
      chn_relu_out_rsci_d_127 <= MUX_s_1_2_2((chn_relu_in_rsci_d_mxwt[127]), (relu_loop_else_relu_loop_else_and_19_nl),
          and_34_cse);
      chn_relu_out_rsci_d_159 <= MUX_s_1_2_2((chn_relu_in_rsci_d_mxwt[159]), (relu_loop_else_relu_loop_else_and_20_nl),
          and_34_cse);
      chn_relu_out_rsci_d_191 <= MUX_s_1_2_2((chn_relu_in_rsci_d_mxwt[191]), (relu_loop_else_relu_loop_else_and_21_nl),
          and_34_cse);
      chn_relu_out_rsci_d_223 <= MUX_s_1_2_2((chn_relu_in_rsci_d_mxwt[223]), (relu_loop_else_relu_loop_else_and_22_nl),
          and_34_cse);
      chn_relu_out_rsci_d_255 <= MUX_s_1_2_2((chn_relu_in_rsci_d_mxwt[255]), (relu_loop_else_relu_loop_else_and_23_nl),
          and_34_cse);
      chn_relu_out_rsci_d_287 <= MUX_s_1_2_2((chn_relu_in_rsci_d_mxwt[287]), (relu_loop_else_relu_loop_else_and_24_nl),
          and_34_cse);
      chn_relu_out_rsci_d_319 <= MUX_s_1_2_2((chn_relu_in_rsci_d_mxwt[319]), (relu_loop_else_relu_loop_else_and_25_nl),
          and_34_cse);
      chn_relu_out_rsci_d_351 <= MUX_s_1_2_2((chn_relu_in_rsci_d_mxwt[351]), (relu_loop_else_relu_loop_else_and_26_nl),
          and_34_cse);
      chn_relu_out_rsci_d_383 <= MUX_s_1_2_2((chn_relu_in_rsci_d_mxwt[383]), (relu_loop_else_relu_loop_else_and_27_nl),
          and_34_cse);
      chn_relu_out_rsci_d_415 <= MUX_s_1_2_2((chn_relu_in_rsci_d_mxwt[415]), (relu_loop_else_relu_loop_else_and_28_nl),
          and_34_cse);
      chn_relu_out_rsci_d_447 <= MUX_s_1_2_2((chn_relu_in_rsci_d_mxwt[447]), (relu_loop_else_relu_loop_else_and_29_nl),
          and_34_cse);
      chn_relu_out_rsci_d_479 <= MUX_s_1_2_2((chn_relu_in_rsci_d_mxwt[479]), (relu_loop_else_relu_loop_else_and_30_nl),
          and_34_cse);
      chn_relu_out_rsci_d_511 <= MUX_s_1_2_2((chn_relu_in_rsci_d_mxwt[511]), (relu_loop_else_relu_loop_else_and_31_nl),
          and_34_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_relu_out_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (or_tmp_85 | and_dcpl_15) ) begin
      reg_chn_relu_out_rsci_ld_core_psct_cse <= ~ and_dcpl_15;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpRelu_8U_23U_lor_lpi_1_dfm <= 1'b0;
      FpRelu_8U_23U_lor_15_lpi_1_dfm <= 1'b0;
      FpRelu_8U_23U_lor_14_lpi_1_dfm <= 1'b0;
      FpRelu_8U_23U_lor_13_lpi_1_dfm <= 1'b0;
      FpRelu_8U_23U_lor_12_lpi_1_dfm <= 1'b0;
      FpRelu_8U_23U_lor_11_lpi_1_dfm <= 1'b0;
      FpRelu_8U_23U_lor_10_lpi_1_dfm <= 1'b0;
      FpRelu_8U_23U_lor_9_lpi_1_dfm <= 1'b0;
      FpRelu_8U_23U_lor_8_lpi_1_dfm <= 1'b0;
      FpRelu_8U_23U_lor_7_lpi_1_dfm <= 1'b0;
      FpRelu_8U_23U_lor_6_lpi_1_dfm <= 1'b0;
      FpRelu_8U_23U_lor_5_lpi_1_dfm <= 1'b0;
      FpRelu_8U_23U_lor_4_lpi_1_dfm <= 1'b0;
      FpRelu_8U_23U_lor_3_lpi_1_dfm <= 1'b0;
      FpRelu_8U_23U_lor_2_lpi_1_dfm <= 1'b0;
      FpRelu_8U_23U_lor_1_lpi_1_dfm <= 1'b0;
    end
    else if ( FpRelu_8U_23U_oelse_and_cse ) begin
      FpRelu_8U_23U_lor_lpi_1_dfm <= FpRelu_8U_23U_lor_lpi_1_dfm_mx0w0;
      FpRelu_8U_23U_lor_15_lpi_1_dfm <= FpRelu_8U_23U_lor_15_lpi_1_dfm_mx0w0;
      FpRelu_8U_23U_lor_14_lpi_1_dfm <= FpRelu_8U_23U_lor_14_lpi_1_dfm_mx0w0;
      FpRelu_8U_23U_lor_13_lpi_1_dfm <= FpRelu_8U_23U_lor_13_lpi_1_dfm_mx0w0;
      FpRelu_8U_23U_lor_12_lpi_1_dfm <= FpRelu_8U_23U_lor_12_lpi_1_dfm_mx0w0;
      FpRelu_8U_23U_lor_11_lpi_1_dfm <= FpRelu_8U_23U_lor_11_lpi_1_dfm_mx0w0;
      FpRelu_8U_23U_lor_10_lpi_1_dfm <= FpRelu_8U_23U_lor_10_lpi_1_dfm_mx0w0;
      FpRelu_8U_23U_lor_9_lpi_1_dfm <= FpRelu_8U_23U_lor_9_lpi_1_dfm_mx0w0;
      FpRelu_8U_23U_lor_8_lpi_1_dfm <= FpRelu_8U_23U_lor_8_lpi_1_dfm_mx0w0;
      FpRelu_8U_23U_lor_7_lpi_1_dfm <= FpRelu_8U_23U_lor_7_lpi_1_dfm_mx0w0;
      FpRelu_8U_23U_lor_6_lpi_1_dfm <= FpRelu_8U_23U_lor_6_lpi_1_dfm_mx0w0;
      FpRelu_8U_23U_lor_5_lpi_1_dfm <= FpRelu_8U_23U_lor_5_lpi_1_dfm_mx0w0;
      FpRelu_8U_23U_lor_4_lpi_1_dfm <= FpRelu_8U_23U_lor_4_lpi_1_dfm_mx0w0;
      FpRelu_8U_23U_lor_3_lpi_1_dfm <= FpRelu_8U_23U_lor_3_lpi_1_dfm_mx0w0;
      FpRelu_8U_23U_lor_2_lpi_1_dfm <= FpRelu_8U_23U_lor_2_lpi_1_dfm_mx0w0;
      FpRelu_8U_23U_lor_1_lpi_1_dfm <= FpRelu_8U_23U_lor_1_lpi_1_dfm_mx0w0;
    end
  end
  assign FpRelu_8U_23U_oelse_mux_32_nl = MUX_s_1_2_2(FpRelu_8U_23U_lor_1_lpi_1_dfm_mx0w0,
      FpRelu_8U_23U_lor_1_lpi_1_dfm, or_dcpl_10);
  assign relu_loop_else_relu_loop_else_and_16_nl = (chn_relu_in_rsci_d_mxwt[31])
      & (FpRelu_8U_23U_oelse_mux_32_nl) & (~ relu_loop_else_unequal_tmp);
  assign FpRelu_8U_23U_oelse_mux_30_nl = MUX_s_1_2_2(FpRelu_8U_23U_lor_2_lpi_1_dfm_mx0w0,
      FpRelu_8U_23U_lor_2_lpi_1_dfm, or_dcpl_10);
  assign relu_loop_else_relu_loop_else_and_17_nl = (chn_relu_in_rsci_d_mxwt[63])
      & (FpRelu_8U_23U_oelse_mux_30_nl) & (~ relu_loop_else_unequal_tmp);
  assign FpRelu_8U_23U_oelse_mux_28_nl = MUX_s_1_2_2(FpRelu_8U_23U_lor_3_lpi_1_dfm_mx0w0,
      FpRelu_8U_23U_lor_3_lpi_1_dfm, or_dcpl_10);
  assign relu_loop_else_relu_loop_else_and_18_nl = (chn_relu_in_rsci_d_mxwt[95])
      & (FpRelu_8U_23U_oelse_mux_28_nl) & (~ relu_loop_else_unequal_tmp);
  assign FpRelu_8U_23U_oelse_mux_26_nl = MUX_s_1_2_2(FpRelu_8U_23U_lor_4_lpi_1_dfm_mx0w0,
      FpRelu_8U_23U_lor_4_lpi_1_dfm, or_dcpl_10);
  assign relu_loop_else_relu_loop_else_and_19_nl = (chn_relu_in_rsci_d_mxwt[127])
      & (FpRelu_8U_23U_oelse_mux_26_nl) & (~ relu_loop_else_unequal_tmp);
  assign FpRelu_8U_23U_oelse_mux_24_nl = MUX_s_1_2_2(FpRelu_8U_23U_lor_5_lpi_1_dfm_mx0w0,
      FpRelu_8U_23U_lor_5_lpi_1_dfm, or_dcpl_10);
  assign relu_loop_else_relu_loop_else_and_20_nl = (chn_relu_in_rsci_d_mxwt[159])
      & (FpRelu_8U_23U_oelse_mux_24_nl) & (~ relu_loop_else_unequal_tmp);
  assign FpRelu_8U_23U_oelse_mux_22_nl = MUX_s_1_2_2(FpRelu_8U_23U_lor_6_lpi_1_dfm_mx0w0,
      FpRelu_8U_23U_lor_6_lpi_1_dfm, or_dcpl_10);
  assign relu_loop_else_relu_loop_else_and_21_nl = (chn_relu_in_rsci_d_mxwt[191])
      & (FpRelu_8U_23U_oelse_mux_22_nl) & (~ relu_loop_else_unequal_tmp);
  assign FpRelu_8U_23U_oelse_mux_20_nl = MUX_s_1_2_2(FpRelu_8U_23U_lor_7_lpi_1_dfm_mx0w0,
      FpRelu_8U_23U_lor_7_lpi_1_dfm, or_dcpl_10);
  assign relu_loop_else_relu_loop_else_and_22_nl = (chn_relu_in_rsci_d_mxwt[223])
      & (FpRelu_8U_23U_oelse_mux_20_nl) & (~ relu_loop_else_unequal_tmp);
  assign FpRelu_8U_23U_oelse_mux_18_nl = MUX_s_1_2_2(FpRelu_8U_23U_lor_8_lpi_1_dfm_mx0w0,
      FpRelu_8U_23U_lor_8_lpi_1_dfm, or_dcpl_10);
  assign relu_loop_else_relu_loop_else_and_23_nl = (chn_relu_in_rsci_d_mxwt[255])
      & (FpRelu_8U_23U_oelse_mux_18_nl) & (~ relu_loop_else_unequal_tmp);
  assign FpRelu_8U_23U_oelse_mux_16_nl = MUX_s_1_2_2(FpRelu_8U_23U_lor_9_lpi_1_dfm_mx0w0,
      FpRelu_8U_23U_lor_9_lpi_1_dfm, or_dcpl_10);
  assign relu_loop_else_relu_loop_else_and_24_nl = (chn_relu_in_rsci_d_mxwt[287])
      & (FpRelu_8U_23U_oelse_mux_16_nl) & (~ relu_loop_else_unequal_tmp);
  assign FpRelu_8U_23U_oelse_mux_14_nl = MUX_s_1_2_2(FpRelu_8U_23U_lor_10_lpi_1_dfm_mx0w0,
      FpRelu_8U_23U_lor_10_lpi_1_dfm, or_dcpl_10);
  assign relu_loop_else_relu_loop_else_and_25_nl = (chn_relu_in_rsci_d_mxwt[319])
      & (FpRelu_8U_23U_oelse_mux_14_nl) & (~ relu_loop_else_unequal_tmp);
  assign FpRelu_8U_23U_oelse_mux_12_nl = MUX_s_1_2_2(FpRelu_8U_23U_lor_11_lpi_1_dfm_mx0w0,
      FpRelu_8U_23U_lor_11_lpi_1_dfm, or_dcpl_10);
  assign relu_loop_else_relu_loop_else_and_26_nl = (chn_relu_in_rsci_d_mxwt[351])
      & (FpRelu_8U_23U_oelse_mux_12_nl) & (~ relu_loop_else_unequal_tmp);
  assign FpRelu_8U_23U_oelse_mux_10_nl = MUX_s_1_2_2(FpRelu_8U_23U_lor_12_lpi_1_dfm_mx0w0,
      FpRelu_8U_23U_lor_12_lpi_1_dfm, or_dcpl_10);
  assign relu_loop_else_relu_loop_else_and_27_nl = (chn_relu_in_rsci_d_mxwt[383])
      & (FpRelu_8U_23U_oelse_mux_10_nl) & (~ relu_loop_else_unequal_tmp);
  assign FpRelu_8U_23U_oelse_mux_8_nl = MUX_s_1_2_2(FpRelu_8U_23U_lor_13_lpi_1_dfm_mx0w0,
      FpRelu_8U_23U_lor_13_lpi_1_dfm, or_dcpl_10);
  assign relu_loop_else_relu_loop_else_and_28_nl = (chn_relu_in_rsci_d_mxwt[415])
      & (FpRelu_8U_23U_oelse_mux_8_nl) & (~ relu_loop_else_unequal_tmp);
  assign FpRelu_8U_23U_oelse_mux_6_nl = MUX_s_1_2_2(FpRelu_8U_23U_lor_14_lpi_1_dfm_mx0w0,
      FpRelu_8U_23U_lor_14_lpi_1_dfm, or_dcpl_10);
  assign relu_loop_else_relu_loop_else_and_29_nl = (chn_relu_in_rsci_d_mxwt[447])
      & (FpRelu_8U_23U_oelse_mux_6_nl) & (~ relu_loop_else_unequal_tmp);
  assign FpRelu_8U_23U_oelse_mux_4_nl = MUX_s_1_2_2(FpRelu_8U_23U_lor_15_lpi_1_dfm_mx0w0,
      FpRelu_8U_23U_lor_15_lpi_1_dfm, or_dcpl_10);
  assign relu_loop_else_relu_loop_else_and_30_nl = (chn_relu_in_rsci_d_mxwt[479])
      & (FpRelu_8U_23U_oelse_mux_4_nl) & (~ relu_loop_else_unequal_tmp);
  assign FpRelu_8U_23U_oelse_mux_2_nl = MUX_s_1_2_2(FpRelu_8U_23U_lor_lpi_1_dfm_mx0w0,
      FpRelu_8U_23U_lor_lpi_1_dfm, or_dcpl_10);
  assign relu_loop_else_relu_loop_else_and_31_nl = (chn_relu_in_rsci_d_mxwt[511])
      & (FpRelu_8U_23U_oelse_mux_2_nl) & (~ relu_loop_else_unequal_tmp);
  function [22:0] MUX1HOT_v_23_3_2;
    input [22:0] input_2;
    input [22:0] input_1;
    input [22:0] input_0;
    input [2:0] sel;
    reg [22:0] result;
  begin
    result = input_0 & {23{sel[0]}};
    result = result | ( input_1 & {23{sel[1]}});
    result = result | ( input_2 & {23{sel[2]}});
    MUX1HOT_v_23_3_2 = result;
  end
  endfunction
  function [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction
  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction
  function [30:0] MUX_v_31_2_2;
    input [30:0] input_0;
    input [30:0] input_1;
    input [0:0] sel;
    reg [30:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_31_2_2 = result;
  end
  endfunction
  function [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction
  function [32:0] conv_s2u_32_33 ;
    input [31:0] vector ;
  begin
    conv_s2u_32_33 = {vector[31], vector};
  end
  endfunction
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_alu
// ------------------------------------------------------------------
module SDP_X_X_alu (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_in_rsc_z, chn_alu_in_rsc_vz, chn_alu_in_rsc_lz,
      chn_alu_op_rsc_z, chn_alu_op_rsc_vz, chn_alu_op_rsc_lz, cfg_alu_op_rsc_z, cfg_alu_op_rsc_triosy_lz,
      cfg_alu_bypass_rsc_z, cfg_alu_bypass_rsc_triosy_lz, cfg_alu_algo_rsc_z, cfg_alu_algo_rsc_triosy_lz,
      cfg_alu_src_rsc_z, cfg_alu_src_rsc_triosy_lz, cfg_alu_shift_value_rsc_z, cfg_alu_shift_value_rsc_triosy_lz,
      cfg_nan_to_zero, cfg_precision, chn_alu_out_rsc_z, chn_alu_out_rsc_vz, chn_alu_out_rsc_lz
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [511:0] chn_alu_in_rsc_z;
  input chn_alu_in_rsc_vz;
  output chn_alu_in_rsc_lz;
  input [255:0] chn_alu_op_rsc_z;
  input chn_alu_op_rsc_vz;
  output chn_alu_op_rsc_lz;
  input [15:0] cfg_alu_op_rsc_z;
  output cfg_alu_op_rsc_triosy_lz;
  input cfg_alu_bypass_rsc_z;
  output cfg_alu_bypass_rsc_triosy_lz;
  input [1:0] cfg_alu_algo_rsc_z;
  output cfg_alu_algo_rsc_triosy_lz;
  input cfg_alu_src_rsc_z;
  output cfg_alu_src_rsc_triosy_lz;
  input [5:0] cfg_alu_shift_value_rsc_z;
  output cfg_alu_shift_value_rsc_triosy_lz;
  input cfg_nan_to_zero;
  input [1:0] cfg_precision;
  output [527:0] chn_alu_out_rsc_z;
  input chn_alu_out_rsc_vz;
  output chn_alu_out_rsc_lz;
// Interconnect Declarations
  wire chn_alu_in_rsci_oswt;
  wire chn_alu_in_rsci_oswt_unreg;
  wire chn_alu_op_rsci_oswt;
  wire chn_alu_op_rsci_oswt_unreg;
  wire [15:0] cfg_alu_op_rsci_d;
  wire cfg_alu_bypass_rsci_d;
  wire [1:0] cfg_alu_algo_rsci_d;
  wire cfg_alu_src_rsci_d;
  wire [5:0] cfg_alu_shift_value_rsci_d;
  wire chn_alu_out_rsci_oswt;
  wire chn_alu_out_rsci_oswt_unreg;
  wire cfg_alu_op_rsc_triosy_obj_oswt;
  wire cfg_alu_bypass_rsc_triosy_obj_oswt;
  wire cfg_alu_algo_rsc_triosy_obj_oswt;
  wire cfg_alu_src_rsc_triosy_obj_oswt;
  wire cfg_alu_shift_value_rsc_triosy_obj_oswt;
  wire cfg_alu_op_rsc_triosy_obj_oswt_unreg_iff;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_in_wire_v1 #(.rscid(32'sd3),
  .width(32'sd16)) cfg_alu_op_rsci (
      .d(cfg_alu_op_rsci_d),
      .z(cfg_alu_op_rsc_z)
    );
  SDP_X_mgc_in_wire_v1 #(.rscid(32'sd4),
  .width(32'sd1)) cfg_alu_bypass_rsci (
      .d(cfg_alu_bypass_rsci_d),
      .z(cfg_alu_bypass_rsc_z)
    );
  SDP_X_mgc_in_wire_v1 #(.rscid(32'sd5),
  .width(32'sd2)) cfg_alu_algo_rsci (
      .d(cfg_alu_algo_rsci_d),
      .z(cfg_alu_algo_rsc_z)
    );
  SDP_X_mgc_in_wire_v1 #(.rscid(32'sd6),
  .width(32'sd1)) cfg_alu_src_rsci (
      .d(cfg_alu_src_rsci_d),
      .z(cfg_alu_src_rsc_z)
    );
  SDP_X_mgc_in_wire_v1 #(.rscid(32'sd7),
  .width(32'sd6)) cfg_alu_shift_value_rsci (
      .d(cfg_alu_shift_value_rsci_d),
      .z(cfg_alu_shift_value_rsc_z)
    );
  SDP_X_chn_alu_in_rsci_unreg chn_alu_in_rsci_unreg_inst (
      .in_0(chn_alu_in_rsci_oswt_unreg),
      .outsig(chn_alu_in_rsci_oswt)
    );
  SDP_X_chn_alu_op_rsci_unreg chn_alu_op_rsci_unreg_inst (
      .in_0(chn_alu_op_rsci_oswt_unreg),
      .outsig(chn_alu_op_rsci_oswt)
    );
  SDP_X_chn_alu_out_rsci_unreg chn_alu_out_rsci_unreg_inst (
      .in_0(chn_alu_out_rsci_oswt_unreg),
      .outsig(chn_alu_out_rsci_oswt)
    );
  SDP_X_cfg_alu_op_rsc_triosy_obj_unreg cfg_alu_op_rsc_triosy_obj_unreg_inst (
      .in_0(cfg_alu_op_rsc_triosy_obj_oswt_unreg_iff),
      .outsig(cfg_alu_op_rsc_triosy_obj_oswt)
    );
  SDP_X_cfg_alu_bypass_rsc_triosy_obj_unreg cfg_alu_bypass_rsc_triosy_obj_unreg_inst (
      .in_0(cfg_alu_op_rsc_triosy_obj_oswt_unreg_iff),
      .outsig(cfg_alu_bypass_rsc_triosy_obj_oswt)
    );
  SDP_X_cfg_alu_algo_rsc_triosy_obj_unreg cfg_alu_algo_rsc_triosy_obj_unreg_inst (
      .in_0(cfg_alu_op_rsc_triosy_obj_oswt_unreg_iff),
      .outsig(cfg_alu_algo_rsc_triosy_obj_oswt)
    );
  SDP_X_cfg_alu_src_rsc_triosy_obj_unreg cfg_alu_src_rsc_triosy_obj_unreg_inst (
      .in_0(cfg_alu_op_rsc_triosy_obj_oswt_unreg_iff),
      .outsig(cfg_alu_src_rsc_triosy_obj_oswt)
    );
  SDP_X_cfg_alu_shift_value_rsc_triosy_obj_unreg cfg_alu_shift_value_rsc_triosy_obj_unreg_inst
      (
      .in_0(cfg_alu_op_rsc_triosy_obj_oswt_unreg_iff),
      .outsig(cfg_alu_shift_value_rsc_triosy_obj_oswt)
    );
  SDP_X_X_alu_core X_alu_core_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_in_rsc_z(chn_alu_in_rsc_z),
      .chn_alu_in_rsc_vz(chn_alu_in_rsc_vz),
      .chn_alu_in_rsc_lz(chn_alu_in_rsc_lz),
      .chn_alu_op_rsc_z(chn_alu_op_rsc_z),
      .chn_alu_op_rsc_vz(chn_alu_op_rsc_vz),
      .chn_alu_op_rsc_lz(chn_alu_op_rsc_lz),
      .cfg_alu_op_rsc_triosy_lz(cfg_alu_op_rsc_triosy_lz),
      .cfg_alu_bypass_rsc_triosy_lz(cfg_alu_bypass_rsc_triosy_lz),
      .cfg_alu_algo_rsc_triosy_lz(cfg_alu_algo_rsc_triosy_lz),
      .cfg_alu_src_rsc_triosy_lz(cfg_alu_src_rsc_triosy_lz),
      .cfg_alu_shift_value_rsc_triosy_lz(cfg_alu_shift_value_rsc_triosy_lz),
      .cfg_nan_to_zero(cfg_nan_to_zero),
      .cfg_precision(cfg_precision),
      .chn_alu_out_rsc_z(chn_alu_out_rsc_z),
      .chn_alu_out_rsc_vz(chn_alu_out_rsc_vz),
      .chn_alu_out_rsc_lz(chn_alu_out_rsc_lz),
      .chn_alu_in_rsci_oswt(chn_alu_in_rsci_oswt),
      .chn_alu_in_rsci_oswt_unreg(chn_alu_in_rsci_oswt_unreg),
      .chn_alu_op_rsci_oswt(chn_alu_op_rsci_oswt),
      .chn_alu_op_rsci_oswt_unreg(chn_alu_op_rsci_oswt_unreg),
      .cfg_alu_op_rsci_d(cfg_alu_op_rsci_d),
      .cfg_alu_bypass_rsci_d(cfg_alu_bypass_rsci_d),
      .cfg_alu_algo_rsci_d(cfg_alu_algo_rsci_d),
      .cfg_alu_src_rsci_d(cfg_alu_src_rsci_d),
      .cfg_alu_shift_value_rsci_d(cfg_alu_shift_value_rsci_d),
      .chn_alu_out_rsci_oswt(chn_alu_out_rsci_oswt),
      .chn_alu_out_rsci_oswt_unreg(chn_alu_out_rsci_oswt_unreg),
      .cfg_alu_op_rsc_triosy_obj_oswt(cfg_alu_op_rsc_triosy_obj_oswt),
      .cfg_alu_bypass_rsc_triosy_obj_oswt(cfg_alu_bypass_rsc_triosy_obj_oswt),
      .cfg_alu_algo_rsc_triosy_obj_oswt(cfg_alu_algo_rsc_triosy_obj_oswt),
      .cfg_alu_src_rsc_triosy_obj_oswt(cfg_alu_src_rsc_triosy_obj_oswt),
      .cfg_alu_shift_value_rsc_triosy_obj_oswt(cfg_alu_shift_value_rsc_triosy_obj_oswt),
      .cfg_alu_op_rsc_triosy_obj_oswt_unreg_pff(cfg_alu_op_rsc_triosy_obj_oswt_unreg_iff)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_mul
// ------------------------------------------------------------------
module SDP_X_X_mul (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_in_rsc_slz, chn_mul_in_rsc_sz, chn_mul_in_rsc_z,
      chn_mul_in_rsc_vz, chn_mul_in_rsc_lz, chn_mul_op_rsc_z, chn_mul_op_rsc_vz,
      chn_mul_op_rsc_lz, cfg_mul_op_rsc_z, cfg_mul_op_rsc_triosy_lz, cfg_mul_bypass_rsc_z,
      cfg_mul_bypass_rsc_triosy_lz, cfg_mul_prelu_rsc_z, cfg_mul_prelu_rsc_triosy_lz,
      cfg_mul_src_rsc_z, cfg_mul_src_rsc_triosy_lz, cfg_nan_to_zero, cfg_precision,
      chn_mul_out_rsc_z, chn_mul_out_rsc_vz, chn_mul_out_rsc_lz
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output chn_mul_in_rsc_slz;
  input chn_mul_in_rsc_sz;
  input [527:0] chn_mul_in_rsc_z;
  input chn_mul_in_rsc_vz;
  output chn_mul_in_rsc_lz;
  input [255:0] chn_mul_op_rsc_z;
  input chn_mul_op_rsc_vz;
  output chn_mul_op_rsc_lz;
  input [15:0] cfg_mul_op_rsc_z;
  output cfg_mul_op_rsc_triosy_lz;
  input cfg_mul_bypass_rsc_z;
  output cfg_mul_bypass_rsc_triosy_lz;
  input cfg_mul_prelu_rsc_z;
  output cfg_mul_prelu_rsc_triosy_lz;
  input cfg_mul_src_rsc_z;
  output cfg_mul_src_rsc_triosy_lz;
  input cfg_nan_to_zero;
  input [1:0] cfg_precision;
  output [799:0] chn_mul_out_rsc_z;
  input chn_mul_out_rsc_vz;
  output chn_mul_out_rsc_lz;
// Interconnect Declarations
  wire chn_mul_in_rsci_oswt;
  wire chn_mul_in_rsci_oswt_unreg;
  wire chn_mul_op_rsci_oswt;
  wire chn_mul_op_rsci_oswt_unreg;
  wire [15:0] cfg_mul_op_rsci_d;
  wire cfg_mul_bypass_rsci_d;
  wire cfg_mul_prelu_rsci_d;
  wire cfg_mul_src_rsci_d;
  wire chn_mul_out_rsci_oswt;
  wire chn_mul_out_rsci_oswt_unreg;
  wire cfg_mul_op_rsc_triosy_obj_oswt;
  wire cfg_mul_bypass_rsc_triosy_obj_oswt;
  wire cfg_mul_prelu_rsc_triosy_obj_oswt;
  wire cfg_mul_src_rsc_triosy_obj_oswt;
  wire cfg_mul_op_rsc_triosy_obj_oswt_unreg_iff;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_in_wire_v1 #(.rscid(32'sd16),
  .width(32'sd16)) cfg_mul_op_rsci (
      .d(cfg_mul_op_rsci_d),
      .z(cfg_mul_op_rsc_z)
    );
  SDP_X_mgc_in_wire_v1 #(.rscid(32'sd17),
  .width(32'sd1)) cfg_mul_bypass_rsci (
      .d(cfg_mul_bypass_rsci_d),
      .z(cfg_mul_bypass_rsc_z)
    );
  SDP_X_mgc_in_wire_v1 #(.rscid(32'sd18),
  .width(32'sd1)) cfg_mul_prelu_rsci (
      .d(cfg_mul_prelu_rsci_d),
      .z(cfg_mul_prelu_rsc_z)
    );
  SDP_X_mgc_in_wire_v1 #(.rscid(32'sd19),
  .width(32'sd1)) cfg_mul_src_rsci (
      .d(cfg_mul_src_rsci_d),
      .z(cfg_mul_src_rsc_z)
    );
  SDP_X_chn_mul_in_rsci_unreg chn_mul_in_rsci_unreg_inst (
      .in_0(chn_mul_in_rsci_oswt_unreg),
      .outsig(chn_mul_in_rsci_oswt)
    );
  SDP_X_chn_mul_op_rsci_unreg chn_mul_op_rsci_unreg_inst (
      .in_0(chn_mul_op_rsci_oswt_unreg),
      .outsig(chn_mul_op_rsci_oswt)
    );
  SDP_X_chn_mul_out_rsci_unreg chn_mul_out_rsci_unreg_inst (
      .in_0(chn_mul_out_rsci_oswt_unreg),
      .outsig(chn_mul_out_rsci_oswt)
    );
  SDP_X_cfg_mul_op_rsc_triosy_obj_unreg cfg_mul_op_rsc_triosy_obj_unreg_inst (
      .in_0(cfg_mul_op_rsc_triosy_obj_oswt_unreg_iff),
      .outsig(cfg_mul_op_rsc_triosy_obj_oswt)
    );
  SDP_X_cfg_mul_bypass_rsc_triosy_obj_unreg cfg_mul_bypass_rsc_triosy_obj_unreg_inst (
      .in_0(cfg_mul_op_rsc_triosy_obj_oswt_unreg_iff),
      .outsig(cfg_mul_bypass_rsc_triosy_obj_oswt)
    );
  SDP_X_cfg_mul_prelu_rsc_triosy_obj_unreg cfg_mul_prelu_rsc_triosy_obj_unreg_inst (
      .in_0(cfg_mul_op_rsc_triosy_obj_oswt_unreg_iff),
      .outsig(cfg_mul_prelu_rsc_triosy_obj_oswt)
    );
  SDP_X_cfg_mul_src_rsc_triosy_obj_unreg cfg_mul_src_rsc_triosy_obj_unreg_inst (
      .in_0(cfg_mul_op_rsc_triosy_obj_oswt_unreg_iff),
      .outsig(cfg_mul_src_rsc_triosy_obj_oswt)
    );
  SDP_X_X_mul_core X_mul_core_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_in_rsc_slz(chn_mul_in_rsc_slz),
      .chn_mul_in_rsc_sz(chn_mul_in_rsc_sz),
      .chn_mul_in_rsc_z(chn_mul_in_rsc_z),
      .chn_mul_in_rsc_vz(chn_mul_in_rsc_vz),
      .chn_mul_in_rsc_lz(chn_mul_in_rsc_lz),
      .chn_mul_op_rsc_z(chn_mul_op_rsc_z),
      .chn_mul_op_rsc_vz(chn_mul_op_rsc_vz),
      .chn_mul_op_rsc_lz(chn_mul_op_rsc_lz),
      .cfg_mul_op_rsc_triosy_lz(cfg_mul_op_rsc_triosy_lz),
      .cfg_mul_bypass_rsc_triosy_lz(cfg_mul_bypass_rsc_triosy_lz),
      .cfg_mul_prelu_rsc_triosy_lz(cfg_mul_prelu_rsc_triosy_lz),
      .cfg_mul_src_rsc_triosy_lz(cfg_mul_src_rsc_triosy_lz),
      .cfg_nan_to_zero(cfg_nan_to_zero),
      .cfg_precision(cfg_precision),
      .chn_mul_out_rsc_z(chn_mul_out_rsc_z),
      .chn_mul_out_rsc_vz(chn_mul_out_rsc_vz),
      .chn_mul_out_rsc_lz(chn_mul_out_rsc_lz),
      .chn_mul_in_rsci_oswt(chn_mul_in_rsci_oswt),
      .chn_mul_in_rsci_oswt_unreg(chn_mul_in_rsci_oswt_unreg),
      .chn_mul_op_rsci_oswt(chn_mul_op_rsci_oswt),
      .chn_mul_op_rsci_oswt_unreg(chn_mul_op_rsci_oswt_unreg),
      .cfg_mul_op_rsci_d(cfg_mul_op_rsci_d),
      .cfg_mul_bypass_rsci_d(cfg_mul_bypass_rsci_d),
      .cfg_mul_prelu_rsci_d(cfg_mul_prelu_rsci_d),
      .cfg_mul_src_rsci_d(cfg_mul_src_rsci_d),
      .chn_mul_out_rsci_oswt(chn_mul_out_rsci_oswt),
      .chn_mul_out_rsci_oswt_unreg(chn_mul_out_rsci_oswt_unreg),
      .cfg_mul_op_rsc_triosy_obj_oswt(cfg_mul_op_rsc_triosy_obj_oswt),
      .cfg_mul_bypass_rsc_triosy_obj_oswt(cfg_mul_bypass_rsc_triosy_obj_oswt),
      .cfg_mul_prelu_rsc_triosy_obj_oswt(cfg_mul_prelu_rsc_triosy_obj_oswt),
      .cfg_mul_src_rsc_triosy_obj_oswt(cfg_mul_src_rsc_triosy_obj_oswt),
      .cfg_mul_op_rsc_triosy_obj_oswt_unreg_pff(cfg_mul_op_rsc_triosy_obj_oswt_unreg_iff)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_trt
// ------------------------------------------------------------------
module SDP_X_X_trt (
  nvdla_core_clk, nvdla_core_rstn, chn_trt_in_rsc_slz, chn_trt_in_rsc_sz, chn_trt_in_rsc_z,
      chn_trt_in_rsc_vz, chn_trt_in_rsc_lz, cfg_mul_shift_value_rsc_z, cfg_mul_shift_value_rsc_triosy_lz,
      cfg_precision, chn_trt_out_rsc_z, chn_trt_out_rsc_vz, chn_trt_out_rsc_lz
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output chn_trt_in_rsc_slz;
  input chn_trt_in_rsc_sz;
  input [799:0] chn_trt_in_rsc_z;
  input chn_trt_in_rsc_vz;
  output chn_trt_in_rsc_lz;
  input [5:0] cfg_mul_shift_value_rsc_z;
  output cfg_mul_shift_value_rsc_triosy_lz;
  input [1:0] cfg_precision;
  output [511:0] chn_trt_out_rsc_z;
  input chn_trt_out_rsc_vz;
  output chn_trt_out_rsc_lz;
// Interconnect Declarations
  wire chn_trt_in_rsci_oswt;
  wire chn_trt_in_rsci_oswt_unreg;
  wire [5:0] cfg_mul_shift_value_rsci_d;
  wire chn_trt_out_rsci_oswt;
  wire cfg_mul_shift_value_rsc_triosy_obj_oswt;
  wire chn_trt_out_rsci_oswt_unreg_iff;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_in_wire_v1 #(.rscid(32'sd28),
  .width(32'sd6)) cfg_mul_shift_value_rsci (
      .d(cfg_mul_shift_value_rsci_d),
      .z(cfg_mul_shift_value_rsc_z)
    );
  SDP_X_chn_trt_in_rsci_unreg chn_trt_in_rsci_unreg_inst (
      .in_0(chn_trt_in_rsci_oswt_unreg),
      .outsig(chn_trt_in_rsci_oswt)
    );
  SDP_X_chn_trt_out_rsci_unreg chn_trt_out_rsci_unreg_inst (
      .in_0(chn_trt_out_rsci_oswt_unreg_iff),
      .outsig(chn_trt_out_rsci_oswt)
    );
  SDP_X_cfg_mul_shift_value_rsc_triosy_obj_unreg cfg_mul_shift_value_rsc_triosy_obj_unreg_inst
      (
      .in_0(chn_trt_out_rsci_oswt_unreg_iff),
      .outsig(cfg_mul_shift_value_rsc_triosy_obj_oswt)
    );
  SDP_X_X_trt_core X_trt_core_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_trt_in_rsc_slz(chn_trt_in_rsc_slz),
      .chn_trt_in_rsc_sz(chn_trt_in_rsc_sz),
      .chn_trt_in_rsc_z(chn_trt_in_rsc_z),
      .chn_trt_in_rsc_vz(chn_trt_in_rsc_vz),
      .chn_trt_in_rsc_lz(chn_trt_in_rsc_lz),
      .cfg_mul_shift_value_rsc_triosy_lz(cfg_mul_shift_value_rsc_triosy_lz),
      .cfg_precision(cfg_precision),
      .chn_trt_out_rsc_z(chn_trt_out_rsc_z),
      .chn_trt_out_rsc_vz(chn_trt_out_rsc_vz),
      .chn_trt_out_rsc_lz(chn_trt_out_rsc_lz),
      .chn_trt_in_rsci_oswt(chn_trt_in_rsci_oswt),
      .chn_trt_in_rsci_oswt_unreg(chn_trt_in_rsci_oswt_unreg),
      .cfg_mul_shift_value_rsci_d(cfg_mul_shift_value_rsci_d),
      .chn_trt_out_rsci_oswt(chn_trt_out_rsci_oswt),
      .cfg_mul_shift_value_rsc_triosy_obj_oswt(cfg_mul_shift_value_rsc_triosy_obj_oswt),
      .chn_trt_out_rsci_oswt_unreg_pff(chn_trt_out_rsci_oswt_unreg_iff)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_X_X_relu
// ------------------------------------------------------------------
module SDP_X_X_relu (
  nvdla_core_clk, nvdla_core_rstn, chn_relu_in_rsc_z, chn_relu_in_rsc_vz, chn_relu_in_rsc_lz,
      cfg_relu_bypass_rsc_z, cfg_relu_bypass_rsc_triosy_lz, cfg_precision, chn_relu_out_rsc_z,
      chn_relu_out_rsc_vz, chn_relu_out_rsc_lz
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [511:0] chn_relu_in_rsc_z;
  input chn_relu_in_rsc_vz;
  output chn_relu_in_rsc_lz;
  input cfg_relu_bypass_rsc_z;
  output cfg_relu_bypass_rsc_triosy_lz;
  input [1:0] cfg_precision;
  output [511:0] chn_relu_out_rsc_z;
  input chn_relu_out_rsc_vz;
  output chn_relu_out_rsc_lz;
// Interconnect Declarations
  wire chn_relu_in_rsci_oswt;
  wire chn_relu_in_rsci_oswt_unreg;
  wire cfg_relu_bypass_rsci_d;
  wire chn_relu_out_rsci_oswt;
  wire cfg_relu_bypass_rsc_triosy_obj_oswt;
  wire chn_relu_out_rsci_oswt_unreg_iff;
// Interconnect Declarations for Component Instantiations
  SDP_X_mgc_in_wire_v1 #(.rscid(32'sd34),
  .width(32'sd1)) cfg_relu_bypass_rsci (
      .d(cfg_relu_bypass_rsci_d),
      .z(cfg_relu_bypass_rsc_z)
    );
  SDP_X_chn_relu_in_rsci_unreg chn_relu_in_rsci_unreg_inst (
      .in_0(chn_relu_in_rsci_oswt_unreg),
      .outsig(chn_relu_in_rsci_oswt)
    );
  SDP_X_chn_relu_out_rsci_unreg chn_relu_out_rsci_unreg_inst (
      .in_0(chn_relu_out_rsci_oswt_unreg_iff),
      .outsig(chn_relu_out_rsci_oswt)
    );
  SDP_X_cfg_relu_bypass_rsc_triosy_obj_unreg cfg_relu_bypass_rsc_triosy_obj_unreg_inst
      (
      .in_0(chn_relu_out_rsci_oswt_unreg_iff),
      .outsig(cfg_relu_bypass_rsc_triosy_obj_oswt)
    );
  SDP_X_X_relu_core X_relu_core_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_relu_in_rsc_z(chn_relu_in_rsc_z),
      .chn_relu_in_rsc_vz(chn_relu_in_rsc_vz),
      .chn_relu_in_rsc_lz(chn_relu_in_rsc_lz),
      .cfg_relu_bypass_rsc_triosy_lz(cfg_relu_bypass_rsc_triosy_lz),
      .cfg_precision(cfg_precision),
      .chn_relu_out_rsc_z(chn_relu_out_rsc_z),
      .chn_relu_out_rsc_vz(chn_relu_out_rsc_vz),
      .chn_relu_out_rsc_lz(chn_relu_out_rsc_lz),
      .chn_relu_in_rsci_oswt(chn_relu_in_rsci_oswt),
      .chn_relu_in_rsci_oswt_unreg(chn_relu_in_rsci_oswt_unreg),
      .cfg_relu_bypass_rsci_d(cfg_relu_bypass_rsci_d),
      .chn_relu_out_rsci_oswt(chn_relu_out_rsci_oswt),
      .cfg_relu_bypass_rsc_triosy_obj_oswt(cfg_relu_bypass_rsc_triosy_obj_oswt),
      .chn_relu_out_rsci_oswt_unreg_pff(chn_relu_out_rsci_oswt_unreg_iff)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_x
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_x (
  nvdla_core_clk, nvdla_core_rstn, chn_data_in_rsc_z, chn_data_in_rsc_vz, chn_data_in_rsc_lz,
      chn_alu_op_rsc_z, chn_alu_op_rsc_vz, chn_alu_op_rsc_lz, chn_mul_op_rsc_z, chn_mul_op_rsc_vz,
      chn_mul_op_rsc_lz, cfg_mul_op_rsc_z, cfg_mul_op_rsc_triosy_lz, cfg_alu_op_rsc_z,
      cfg_alu_op_rsc_triosy_lz, cfg_alu_bypass_rsc_z, cfg_alu_bypass_rsc_triosy_lz,
      cfg_alu_algo_rsc_z, cfg_alu_algo_rsc_triosy_lz, cfg_alu_src_rsc_z, cfg_alu_src_rsc_triosy_lz,
      cfg_alu_shift_value_rsc_z, cfg_alu_shift_value_rsc_triosy_lz, cfg_mul_bypass_rsc_z,
      cfg_mul_bypass_rsc_triosy_lz, cfg_mul_prelu_rsc_z, cfg_mul_prelu_rsc_triosy_lz,
      cfg_mul_src_rsc_z, cfg_mul_src_rsc_triosy_lz, cfg_mul_shift_value_rsc_z, cfg_mul_shift_value_rsc_triosy_lz,
      cfg_relu_bypass_rsc_z, cfg_relu_bypass_rsc_triosy_lz, cfg_nan_to_zero, cfg_precision,
      chn_data_out_rsc_z, chn_data_out_rsc_vz, chn_data_out_rsc_lz
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [511:0] chn_data_in_rsc_z;
  input chn_data_in_rsc_vz;
  output chn_data_in_rsc_lz;
  input [255:0] chn_alu_op_rsc_z;
  input chn_alu_op_rsc_vz;
  output chn_alu_op_rsc_lz;
  input [255:0] chn_mul_op_rsc_z;
  input chn_mul_op_rsc_vz;
  output chn_mul_op_rsc_lz;
  input [15:0] cfg_mul_op_rsc_z;
  output cfg_mul_op_rsc_triosy_lz;
  input [15:0] cfg_alu_op_rsc_z;
  output cfg_alu_op_rsc_triosy_lz;
  input cfg_alu_bypass_rsc_z;
  output cfg_alu_bypass_rsc_triosy_lz;
  input [1:0] cfg_alu_algo_rsc_z;
  output cfg_alu_algo_rsc_triosy_lz;
  input cfg_alu_src_rsc_z;
  output cfg_alu_src_rsc_triosy_lz;
  input [5:0] cfg_alu_shift_value_rsc_z;
  output cfg_alu_shift_value_rsc_triosy_lz;
  input cfg_mul_bypass_rsc_z;
  output cfg_mul_bypass_rsc_triosy_lz;
  input cfg_mul_prelu_rsc_z;
  output cfg_mul_prelu_rsc_triosy_lz;
  input cfg_mul_src_rsc_z;
  output cfg_mul_src_rsc_triosy_lz;
  input [5:0] cfg_mul_shift_value_rsc_z;
  output cfg_mul_shift_value_rsc_triosy_lz;
  input cfg_relu_bypass_rsc_z;
  output cfg_relu_bypass_rsc_triosy_lz;
  input cfg_nan_to_zero;
  input [1:0] cfg_precision;
  output [511:0] chn_data_out_rsc_z;
  input chn_data_out_rsc_vz;
  output chn_data_out_rsc_lz;
// Interconnect Declarations
  wire [527:0] chn_alu_out_rsc_z_nX_alu_inst;
  wire chn_alu_out_rsc_vz_nX_alu_inst;
  wire [1:0] chn_mul_in_rsc_sz_nX_mul_inst;
  wire [527:0] chn_mul_in_rsc_z_nX_mul_inst;
  wire chn_mul_in_rsc_vz_nX_mul_inst;
  wire [799:0] chn_mul_out_rsc_z_nX_mul_inst;
  wire chn_mul_out_rsc_vz_nX_mul_inst;
  wire [1:0] chn_trt_in_rsc_sz_nX_trt_inst;
  wire [799:0] chn_trt_in_rsc_z_nX_trt_inst;
  wire chn_trt_in_rsc_vz_nX_trt_inst;
  wire [511:0] chn_trt_out_rsc_z_nX_trt_inst;
  wire chn_trt_out_rsc_vz_nX_trt_inst;
  wire [511:0] chn_relu_in_rsc_z_nX_relu_inst;
  wire chn_relu_in_rsc_vz_nX_relu_inst;
  wire [511:0] chn_relu_out_rsc_z_nX_relu_inst;
  wire chn_alu_in_rsc_lz_nX_alu_inst_bud;
  wire chn_alu_op_rsc_lz_nX_alu_inst_bud;
  wire cfg_alu_op_rsc_triosy_lz_nX_alu_inst_bud;
  wire cfg_alu_bypass_rsc_triosy_lz_nX_alu_inst_bud;
  wire cfg_alu_algo_rsc_triosy_lz_nX_alu_inst_bud;
  wire cfg_alu_src_rsc_triosy_lz_nX_alu_inst_bud;
  wire cfg_alu_shift_value_rsc_triosy_lz_nX_alu_inst_bud;
  wire chn_alu_out_rsc_lz_nX_alu_inst_bud;
  wire chn_mul_in_rsc_lz_nX_mul_inst_bud;
  wire chn_mul_in_rsc_slz_nX_mul_inst_bud;
  wire chn_mul_op_rsc_lz_nX_mul_inst_bud;
  wire cfg_mul_op_rsc_triosy_lz_nX_mul_inst_bud;
  wire cfg_mul_bypass_rsc_triosy_lz_nX_mul_inst_bud;
  wire cfg_mul_prelu_rsc_triosy_lz_nX_mul_inst_bud;
  wire cfg_mul_src_rsc_triosy_lz_nX_mul_inst_bud;
  wire chn_mul_out_rsc_lz_nX_mul_inst_bud;
  wire chn_trt_in_rsc_lz_nX_trt_inst_bud;
  wire chn_trt_in_rsc_slz_nX_trt_inst_bud;
  wire cfg_mul_shift_value_rsc_triosy_lz_nX_trt_inst_bud;
  wire chn_trt_out_rsc_lz_nX_trt_inst_bud;
  wire chn_relu_in_rsc_lz_nX_relu_inst_bud;
  wire cfg_relu_bypass_rsc_triosy_lz_nX_relu_inst_bud;
  wire chn_relu_out_rsc_lz_nX_relu_inst_bud;
  wire chn_trt_out_unc_2;
// Interconnect Declarations for Component Instantiations
  wire [0:0] nl_X_mul_inst_chn_mul_in_rsc_sz;
  assign nl_X_mul_inst_chn_mul_in_rsc_sz = chn_mul_in_rsc_sz_nX_mul_inst[0];
  wire [0:0] nl_X_trt_inst_chn_trt_in_rsc_sz;
  assign nl_X_trt_inst_chn_trt_in_rsc_sz = chn_trt_in_rsc_sz_nX_trt_inst[0];
  SDP_X_mgc_pipe_v10 #(.rscid(32'sd56),
  .width(32'sd528),
  .sz_width(32'sd2),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) chn_alu_out_cns_pipe (
      .clk(nvdla_core_clk),
      .en(1'b0),
      .arst(nvdla_core_rstn),
      .srst(1'b1),
      .ldin(chn_mul_in_rsc_lz_nX_mul_inst_bud),
      .vdin(chn_mul_in_rsc_vz_nX_mul_inst),
      .din(chn_mul_in_rsc_z_nX_mul_inst),
      .ldout(chn_alu_out_rsc_lz_nX_alu_inst_bud),
      .vdout(chn_alu_out_rsc_vz_nX_alu_inst),
      .dout(chn_alu_out_rsc_z_nX_alu_inst),
      .sd(chn_mul_in_rsc_sz_nX_mul_inst)
    );
  SDP_X_mgc_pipe_v10 #(.rscid(32'sd57),
  .width(32'sd800),
  .sz_width(32'sd2),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) chn_mul_out_cns_pipe (
      .clk(nvdla_core_clk),
      .en(1'b0),
      .arst(nvdla_core_rstn),
      .srst(1'b1),
      .ldin(chn_trt_in_rsc_lz_nX_trt_inst_bud),
      .vdin(chn_trt_in_rsc_vz_nX_trt_inst),
      .din(chn_trt_in_rsc_z_nX_trt_inst),
      .ldout(chn_mul_out_rsc_lz_nX_mul_inst_bud),
      .vdout(chn_mul_out_rsc_vz_nX_mul_inst),
      .dout(chn_mul_out_rsc_z_nX_mul_inst),
      .sd(chn_trt_in_rsc_sz_nX_trt_inst)
    );
  SDP_X_mgc_pipe_v10 #(.rscid(32'sd58),
  .width(32'sd512),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) chn_trt_out_cns_pipe (
      .clk(nvdla_core_clk),
      .en(1'b0),
      .arst(nvdla_core_rstn),
      .srst(1'b1),
      .ldin(chn_relu_in_rsc_lz_nX_relu_inst_bud),
      .vdin(chn_relu_in_rsc_vz_nX_relu_inst),
      .din(chn_relu_in_rsc_z_nX_relu_inst),
      .ldout(chn_trt_out_rsc_lz_nX_trt_inst_bud),
      .vdout(chn_trt_out_rsc_vz_nX_trt_inst),
      .dout(chn_trt_out_rsc_z_nX_trt_inst),
      .sd(chn_trt_out_unc_2)
    );
  SDP_X_X_alu X_alu_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_in_rsc_z(chn_data_in_rsc_z),
      .chn_alu_in_rsc_vz(chn_data_in_rsc_vz),
      .chn_alu_in_rsc_lz(chn_alu_in_rsc_lz_nX_alu_inst_bud),
      .chn_alu_op_rsc_z(chn_alu_op_rsc_z),
      .chn_alu_op_rsc_vz(chn_alu_op_rsc_vz),
      .chn_alu_op_rsc_lz(chn_alu_op_rsc_lz_nX_alu_inst_bud),
      .cfg_alu_op_rsc_z(cfg_alu_op_rsc_z),
      .cfg_alu_op_rsc_triosy_lz(cfg_alu_op_rsc_triosy_lz_nX_alu_inst_bud),
      .cfg_alu_bypass_rsc_z(cfg_alu_bypass_rsc_z),
      .cfg_alu_bypass_rsc_triosy_lz(cfg_alu_bypass_rsc_triosy_lz_nX_alu_inst_bud),
      .cfg_alu_algo_rsc_z(cfg_alu_algo_rsc_z),
      .cfg_alu_algo_rsc_triosy_lz(cfg_alu_algo_rsc_triosy_lz_nX_alu_inst_bud),
      .cfg_alu_src_rsc_z(cfg_alu_src_rsc_z),
      .cfg_alu_src_rsc_triosy_lz(cfg_alu_src_rsc_triosy_lz_nX_alu_inst_bud),
      .cfg_alu_shift_value_rsc_z(cfg_alu_shift_value_rsc_z),
      .cfg_alu_shift_value_rsc_triosy_lz(cfg_alu_shift_value_rsc_triosy_lz_nX_alu_inst_bud),
      .cfg_nan_to_zero(cfg_nan_to_zero),
      .cfg_precision(cfg_precision),
      .chn_alu_out_rsc_z(chn_alu_out_rsc_z_nX_alu_inst),
      .chn_alu_out_rsc_vz(chn_alu_out_rsc_vz_nX_alu_inst),
      .chn_alu_out_rsc_lz(chn_alu_out_rsc_lz_nX_alu_inst_bud)
    );
  SDP_X_X_mul X_mul_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_in_rsc_slz(chn_mul_in_rsc_slz_nX_mul_inst_bud),
      .chn_mul_in_rsc_sz(nl_X_mul_inst_chn_mul_in_rsc_sz[0:0]),
      .chn_mul_in_rsc_z(chn_mul_in_rsc_z_nX_mul_inst),
      .chn_mul_in_rsc_vz(chn_mul_in_rsc_vz_nX_mul_inst),
      .chn_mul_in_rsc_lz(chn_mul_in_rsc_lz_nX_mul_inst_bud),
      .chn_mul_op_rsc_z(chn_mul_op_rsc_z),
      .chn_mul_op_rsc_vz(chn_mul_op_rsc_vz),
      .chn_mul_op_rsc_lz(chn_mul_op_rsc_lz_nX_mul_inst_bud),
      .cfg_mul_op_rsc_z(cfg_mul_op_rsc_z),
      .cfg_mul_op_rsc_triosy_lz(cfg_mul_op_rsc_triosy_lz_nX_mul_inst_bud),
      .cfg_mul_bypass_rsc_z(cfg_mul_bypass_rsc_z),
      .cfg_mul_bypass_rsc_triosy_lz(cfg_mul_bypass_rsc_triosy_lz_nX_mul_inst_bud),
      .cfg_mul_prelu_rsc_z(cfg_mul_prelu_rsc_z),
      .cfg_mul_prelu_rsc_triosy_lz(cfg_mul_prelu_rsc_triosy_lz_nX_mul_inst_bud),
      .cfg_mul_src_rsc_z(cfg_mul_src_rsc_z),
      .cfg_mul_src_rsc_triosy_lz(cfg_mul_src_rsc_triosy_lz_nX_mul_inst_bud),
      .cfg_nan_to_zero(cfg_nan_to_zero),
      .cfg_precision(cfg_precision),
      .chn_mul_out_rsc_z(chn_mul_out_rsc_z_nX_mul_inst),
      .chn_mul_out_rsc_vz(chn_mul_out_rsc_vz_nX_mul_inst),
      .chn_mul_out_rsc_lz(chn_mul_out_rsc_lz_nX_mul_inst_bud)
    );
  SDP_X_X_trt X_trt_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_trt_in_rsc_slz(chn_trt_in_rsc_slz_nX_trt_inst_bud),
      .chn_trt_in_rsc_sz(nl_X_trt_inst_chn_trt_in_rsc_sz[0:0]),
      .chn_trt_in_rsc_z(chn_trt_in_rsc_z_nX_trt_inst),
      .chn_trt_in_rsc_vz(chn_trt_in_rsc_vz_nX_trt_inst),
      .chn_trt_in_rsc_lz(chn_trt_in_rsc_lz_nX_trt_inst_bud),
      .cfg_mul_shift_value_rsc_z(cfg_mul_shift_value_rsc_z),
      .cfg_mul_shift_value_rsc_triosy_lz(cfg_mul_shift_value_rsc_triosy_lz_nX_trt_inst_bud),
      .cfg_precision(cfg_precision),
      .chn_trt_out_rsc_z(chn_trt_out_rsc_z_nX_trt_inst),
      .chn_trt_out_rsc_vz(chn_trt_out_rsc_vz_nX_trt_inst),
      .chn_trt_out_rsc_lz(chn_trt_out_rsc_lz_nX_trt_inst_bud)
    );
  SDP_X_X_relu X_relu_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_relu_in_rsc_z(chn_relu_in_rsc_z_nX_relu_inst),
      .chn_relu_in_rsc_vz(chn_relu_in_rsc_vz_nX_relu_inst),
      .chn_relu_in_rsc_lz(chn_relu_in_rsc_lz_nX_relu_inst_bud),
      .cfg_relu_bypass_rsc_z(cfg_relu_bypass_rsc_z),
      .cfg_relu_bypass_rsc_triosy_lz(cfg_relu_bypass_rsc_triosy_lz_nX_relu_inst_bud),
      .cfg_precision(cfg_precision),
      .chn_relu_out_rsc_z(chn_relu_out_rsc_z_nX_relu_inst),
      .chn_relu_out_rsc_vz(chn_data_out_rsc_vz),
      .chn_relu_out_rsc_lz(chn_relu_out_rsc_lz_nX_relu_inst_bud)
    );
  assign chn_data_in_rsc_lz = chn_alu_in_rsc_lz_nX_alu_inst_bud;
  assign chn_alu_op_rsc_lz = chn_alu_op_rsc_lz_nX_alu_inst_bud;
  assign cfg_alu_op_rsc_triosy_lz = cfg_alu_op_rsc_triosy_lz_nX_alu_inst_bud;
  assign cfg_alu_bypass_rsc_triosy_lz = cfg_alu_bypass_rsc_triosy_lz_nX_alu_inst_bud;
  assign cfg_alu_algo_rsc_triosy_lz = cfg_alu_algo_rsc_triosy_lz_nX_alu_inst_bud;
  assign cfg_alu_src_rsc_triosy_lz = cfg_alu_src_rsc_triosy_lz_nX_alu_inst_bud;
  assign cfg_alu_shift_value_rsc_triosy_lz = cfg_alu_shift_value_rsc_triosy_lz_nX_alu_inst_bud;
  assign chn_mul_op_rsc_lz = chn_mul_op_rsc_lz_nX_mul_inst_bud;
  assign cfg_mul_op_rsc_triosy_lz = cfg_mul_op_rsc_triosy_lz_nX_mul_inst_bud;
  assign cfg_mul_bypass_rsc_triosy_lz = cfg_mul_bypass_rsc_triosy_lz_nX_mul_inst_bud;
  assign cfg_mul_prelu_rsc_triosy_lz = cfg_mul_prelu_rsc_triosy_lz_nX_mul_inst_bud;
  assign cfg_mul_src_rsc_triosy_lz = cfg_mul_src_rsc_triosy_lz_nX_mul_inst_bud;
  assign cfg_mul_shift_value_rsc_triosy_lz = cfg_mul_shift_value_rsc_triosy_lz_nX_trt_inst_bud;
  assign cfg_relu_bypass_rsc_triosy_lz = cfg_relu_bypass_rsc_triosy_lz_nX_relu_inst_bud;
  assign chn_data_out_rsc_lz = chn_relu_out_rsc_lz_nX_relu_inst_bud;
  assign chn_data_out_rsc_z = chn_relu_out_rsc_z_nX_relu_inst;
endmodule
